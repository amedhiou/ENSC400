
module up_island_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  OAI21_X4 U1 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  AOI21_X4 U3 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  AOI21_X4 U7 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  OAI21_X4 U9 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  NOR2_X4 U10 ( .A1(n151), .A2(B[31]), .ZN(n14) );
  NAND2_X4 U11 ( .A1(n151), .A2(B[31]), .ZN(n15) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U14 ( .A1(n22), .A2(n20), .ZN(n18) );
  OAI21_X4 U15 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  AOI21_X4 U21 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  NOR2_X4 U22 ( .A1(n28), .A2(n26), .ZN(n24) );
  OAI21_X4 U23 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U28 ( .A1(n34), .A2(n32), .ZN(n30) );
  OAI21_X4 U29 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NAND2_X4 U33 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  OAI21_X4 U35 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NOR2_X4 U48 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  NAND2_X4 U49 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  NAND2_X4 U50 ( .A1(n58), .A2(n52), .ZN(n50) );
  AOI21_X4 U51 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NOR2_X4 U52 ( .A1(n56), .A2(n54), .ZN(n52) );
  OAI21_X4 U53 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X4 U54 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NAND2_X4 U55 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X4 U56 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X4 U57 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  NOR2_X4 U60 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NAND2_X4 U61 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X4 U62 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X4 U63 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U71 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  NAND2_X4 U72 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X4 U73 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NAND2_X4 U74 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NOR2_X4 U77 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  NAND2_X4 U78 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X4 U79 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X4 U80 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U85 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  NAND2_X4 U86 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X4 U87 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NAND2_X4 U88 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  NOR2_X4 U91 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X4 U92 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X4 U93 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X4 U94 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U100 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NAND2_X4 U101 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X4 U102 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  NAND2_X4 U103 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  NOR2_X4 U106 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  NAND2_X4 U107 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X4 U108 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  NAND2_X4 U109 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  INV_X32 U121 ( .A(A[31]), .ZN(n151) );
  INV_X1 U157 ( .A(A[18]), .ZN(n138) );
  INV_X1 U158 ( .A(A[15]), .ZN(n135) );
  INV_X1 U159 ( .A(A[19]), .ZN(n139) );
  INV_X1 U160 ( .A(A[20]), .ZN(n140) );
  INV_X1 U161 ( .A(A[21]), .ZN(n141) );
  INV_X1 U162 ( .A(A[9]), .ZN(n129) );
  INV_X1 U163 ( .A(A[10]), .ZN(n130) );
  INV_X1 U164 ( .A(A[22]), .ZN(n142) );
  INV_X1 U165 ( .A(A[23]), .ZN(n143) );
  INV_X1 U166 ( .A(A[8]), .ZN(n128) );
  INV_X1 U167 ( .A(A[16]), .ZN(n136) );
  INV_X1 U168 ( .A(A[17]), .ZN(n137) );
  INV_X1 U169 ( .A(A[28]), .ZN(n148) );
  INV_X1 U170 ( .A(A[27]), .ZN(n147) );
  INV_X1 U171 ( .A(A[25]), .ZN(n145) );
  INV_X1 U172 ( .A(A[30]), .ZN(n150) );
  INV_X1 U173 ( .A(A[7]), .ZN(n127) );
  INV_X1 U174 ( .A(A[14]), .ZN(n134) );
  INV_X1 U175 ( .A(A[13]), .ZN(n133) );
  INV_X1 U176 ( .A(A[11]), .ZN(n131) );
  INV_X1 U177 ( .A(A[12]), .ZN(n132) );
  INV_X1 U178 ( .A(A[29]), .ZN(n149) );
  INV_X1 U179 ( .A(A[5]), .ZN(n125) );
  INV_X1 U180 ( .A(A[26]), .ZN(n146) );
  INV_X1 U181 ( .A(A[24]), .ZN(n144) );
  INV_X1 U182 ( .A(A[6]), .ZN(n126) );
  INV_X4 U183 ( .A(A[4]), .ZN(n124) );
  INV_X1 U184 ( .A(A[1]), .ZN(n121) );
  INV_X1 U185 ( .A(A[3]), .ZN(n123) );
  INV_X4 U186 ( .A(A[2]), .ZN(n122) );
  NAND2_X1 U187 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NOR2_X1 U188 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X1 U189 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  INV_X1 U190 ( .A(A[0]), .ZN(n120) );
endmodule


module up_island_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  OAI21_X4 U1 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  AOI21_X4 U3 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  AOI21_X4 U7 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  OAI21_X4 U9 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  NOR2_X4 U10 ( .A1(n151), .A2(A[31]), .ZN(n14) );
  NAND2_X4 U11 ( .A1(n151), .A2(A[31]), .ZN(n15) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U14 ( .A1(n22), .A2(n20), .ZN(n18) );
  OAI21_X4 U15 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  AOI21_X4 U21 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  NOR2_X4 U22 ( .A1(n28), .A2(n26), .ZN(n24) );
  OAI21_X4 U23 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U28 ( .A1(n34), .A2(n32), .ZN(n30) );
  OAI21_X4 U29 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NAND2_X4 U33 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  OAI21_X4 U35 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NOR2_X4 U48 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  NAND2_X4 U49 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  NAND2_X4 U50 ( .A1(n58), .A2(n52), .ZN(n50) );
  AOI21_X4 U51 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NOR2_X4 U52 ( .A1(n56), .A2(n54), .ZN(n52) );
  OAI21_X4 U53 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X4 U54 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NAND2_X4 U55 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X4 U56 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X4 U57 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  NOR2_X4 U60 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NAND2_X4 U61 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X4 U62 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X4 U63 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U71 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  NAND2_X4 U72 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X4 U73 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NAND2_X4 U74 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NOR2_X4 U77 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  NAND2_X4 U78 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X4 U79 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X4 U80 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U85 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  NAND2_X4 U86 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X4 U87 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NAND2_X4 U88 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  NOR2_X4 U91 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X4 U92 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X4 U93 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X4 U94 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U100 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NAND2_X4 U101 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X4 U102 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  NAND2_X4 U103 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  NOR2_X4 U106 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  NAND2_X4 U107 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X4 U108 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  NAND2_X4 U109 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  INV_X32 U152 ( .A(B[31]), .ZN(n151) );
  INV_X1 U157 ( .A(A[18]), .ZN(n138) );
  INV_X1 U158 ( .A(A[15]), .ZN(n135) );
  INV_X1 U159 ( .A(A[19]), .ZN(n139) );
  INV_X1 U160 ( .A(A[20]), .ZN(n140) );
  INV_X1 U161 ( .A(A[21]), .ZN(n141) );
  INV_X1 U162 ( .A(A[9]), .ZN(n129) );
  INV_X1 U163 ( .A(A[10]), .ZN(n130) );
  INV_X1 U164 ( .A(A[22]), .ZN(n142) );
  INV_X1 U165 ( .A(A[23]), .ZN(n143) );
  INV_X1 U166 ( .A(A[8]), .ZN(n128) );
  INV_X1 U167 ( .A(A[16]), .ZN(n136) );
  INV_X1 U168 ( .A(A[17]), .ZN(n137) );
  INV_X1 U169 ( .A(A[28]), .ZN(n148) );
  INV_X1 U170 ( .A(A[27]), .ZN(n147) );
  INV_X1 U171 ( .A(A[25]), .ZN(n145) );
  INV_X1 U172 ( .A(A[30]), .ZN(n150) );
  INV_X1 U173 ( .A(A[7]), .ZN(n127) );
  INV_X1 U174 ( .A(A[14]), .ZN(n134) );
  INV_X1 U175 ( .A(A[13]), .ZN(n133) );
  INV_X1 U176 ( .A(A[11]), .ZN(n131) );
  INV_X1 U177 ( .A(A[12]), .ZN(n132) );
  INV_X1 U178 ( .A(A[29]), .ZN(n149) );
  INV_X1 U179 ( .A(A[5]), .ZN(n125) );
  INV_X1 U180 ( .A(A[26]), .ZN(n146) );
  INV_X1 U181 ( .A(A[24]), .ZN(n144) );
  INV_X1 U182 ( .A(A[6]), .ZN(n126) );
  INV_X4 U183 ( .A(A[4]), .ZN(n124) );
  INV_X1 U184 ( .A(A[1]), .ZN(n121) );
  INV_X1 U185 ( .A(A[3]), .ZN(n123) );
  INV_X4 U186 ( .A(A[2]), .ZN(n122) );
  NAND2_X1 U187 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NOR2_X1 U188 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X1 U189 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  INV_X1 U190 ( .A(A[0]), .ZN(n120) );
endmodule


module up_island_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604;

  INV_X1 U173 ( .A(A[18]), .ZN(n549) );
  NAND2_X1 U174 ( .A1(A[15]), .A2(n378), .ZN(n555) );
  INV_X1 U175 ( .A(A[19]), .ZN(n542) );
  INV_X1 U176 ( .A(A[20]), .ZN(n529) );
  INV_X1 U177 ( .A(A[21]), .ZN(n522) );
  INV_X1 U178 ( .A(A[9]), .ZN(n494) );
  NAND2_X1 U179 ( .A1(A[9]), .A2(n377), .ZN(n595) );
  INV_X1 U180 ( .A(A[10]), .ZN(n486) );
  NAND2_X1 U181 ( .A1(A[10]), .A2(n377), .ZN(n587) );
  INV_X1 U182 ( .A(A[22]), .ZN(n515) );
  INV_X1 U183 ( .A(A[23]), .ZN(n508) );
  INV_X1 U184 ( .A(A[8]), .ZN(n502) );
  NAND2_X1 U185 ( .A1(A[8]), .A2(n377), .ZN(n583) );
  INV_X1 U186 ( .A(A[16]), .ZN(n563) );
  INV_X1 U187 ( .A(A[17]), .ZN(n556) );
  INV_X1 U188 ( .A(A[28]), .ZN(n469) );
  INV_X1 U189 ( .A(A[27]), .ZN(n477) );
  INV_X1 U190 ( .A(A[25]), .ZN(n493) );
  INV_X1 U191 ( .A(A[30]), .ZN(n446) );
  INV_X1 U192 ( .A(A[7]), .ZN(n509) );
  NAND2_X1 U193 ( .A1(A[7]), .A2(n377), .ZN(n591) );
  INV_X1 U194 ( .A(A[14]), .ZN(n447) );
  NAND2_X1 U195 ( .A1(A[14]), .A2(n378), .ZN(n562) );
  INV_X1 U196 ( .A(A[13]), .ZN(n461) );
  NAND2_X1 U197 ( .A1(A[13]), .A2(n378), .ZN(n569) );
  INV_X1 U198 ( .A(A[11]), .ZN(n478) );
  NAND2_X1 U199 ( .A1(A[11]), .A2(n377), .ZN(n579) );
  INV_X1 U200 ( .A(A[12]), .ZN(n470) );
  NAND2_X1 U201 ( .A1(A[12]), .A2(n378), .ZN(n574) );
  INV_X1 U202 ( .A(A[29]), .ZN(n460) );
  INV_X1 U203 ( .A(A[5]), .ZN(n523) );
  NAND2_X1 U204 ( .A1(A[5]), .A2(n377), .ZN(n592) );
  INV_X1 U205 ( .A(A[26]), .ZN(n485) );
  INV_X1 U206 ( .A(A[24]), .ZN(n501) );
  INV_X1 U207 ( .A(A[6]), .ZN(n516) );
  NAND2_X1 U208 ( .A1(A[6]), .A2(n377), .ZN(n584) );
  INV_X1 U209 ( .A(A[4]), .ZN(n530) );
  NAND2_X1 U210 ( .A1(A[4]), .A2(n377), .ZN(n585) );
  NAND2_X1 U211 ( .A1(A[3]), .A2(n377), .ZN(n593) );
  INV_X1 U212 ( .A(A[3]), .ZN(n543) );
  INV_X1 U213 ( .A(A[2]), .ZN(n550) );
  NAND2_X1 U214 ( .A1(A[2]), .A2(n377), .ZN(n586) );
  INV_X1 U215 ( .A(A[0]), .ZN(n564) );
  NAND2_X1 U216 ( .A1(A[0]), .A2(n377), .ZN(n601) );
  NAND2_X1 U217 ( .A1(A[1]), .A2(n377), .ZN(n594) );
  INV_X1 U218 ( .A(A[1]), .ZN(n557) );
  INV_X1 U219 ( .A(SH[4]), .ZN(n377) );
  INV_X1 U220 ( .A(SH[4]), .ZN(n378) );
  INV_X1 U221 ( .A(n385), .ZN(n379) );
  INV_X1 U222 ( .A(n385), .ZN(n380) );
  INV_X1 U223 ( .A(SH[3]), .ZN(n381) );
  INV_X1 U224 ( .A(SH[3]), .ZN(n382) );
  INV_X1 U225 ( .A(SH[3]), .ZN(n383) );
  INV_X1 U226 ( .A(SH[3]), .ZN(n384) );
  INV_X1 U227 ( .A(SH[3]), .ZN(n385) );
  INV_X1 U228 ( .A(n391), .ZN(n386) );
  INV_X1 U229 ( .A(n391), .ZN(n387) );
  INV_X1 U230 ( .A(n391), .ZN(n388) );
  INV_X1 U231 ( .A(SH[2]), .ZN(n389) );
  INV_X1 U232 ( .A(SH[2]), .ZN(n390) );
  INV_X1 U233 ( .A(SH[2]), .ZN(n391) );
  INV_X1 U234 ( .A(n396), .ZN(n392) );
  INV_X1 U235 ( .A(n396), .ZN(n393) );
  INV_X1 U236 ( .A(n396), .ZN(n394) );
  INV_X1 U237 ( .A(SH[1]), .ZN(n395) );
  INV_X1 U238 ( .A(SH[1]), .ZN(n396) );
  BUF_X1 U239 ( .A(SH[0]), .Z(n397) );
  BUF_X1 U240 ( .A(SH[0]), .Z(n398) );
  MUX2_X1 U241 ( .A(n399), .B(n400), .S(n398), .Z(B[9]) );
  MUX2_X1 U242 ( .A(n400), .B(n401), .S(n398), .Z(B[8]) );
  INV_X2 U243 ( .A(n402), .ZN(n400) );
  MUX2_X1 U244 ( .A(n403), .B(n404), .S(n386), .Z(n402) );
  MUX2_X1 U245 ( .A(n401), .B(n405), .S(n398), .Z(B[7]) );
  INV_X2 U246 ( .A(n406), .ZN(n401) );
  MUX2_X1 U247 ( .A(n407), .B(n408), .S(n386), .Z(n406) );
  MUX2_X1 U248 ( .A(n405), .B(n409), .S(n398), .Z(B[6]) );
  INV_X2 U249 ( .A(n410), .ZN(n405) );
  MUX2_X1 U250 ( .A(n411), .B(n412), .S(n386), .Z(n410) );
  MUX2_X1 U251 ( .A(n409), .B(n413), .S(n398), .Z(B[5]) );
  INV_X2 U252 ( .A(n414), .ZN(n409) );
  MUX2_X1 U253 ( .A(n415), .B(n416), .S(n386), .Z(n414) );
  MUX2_X1 U254 ( .A(n413), .B(n417), .S(n398), .Z(B[4]) );
  INV_X2 U255 ( .A(n418), .ZN(n413) );
  MUX2_X1 U256 ( .A(n404), .B(n419), .S(n386), .Z(n418) );
  NAND2_X2 U257 ( .A1(n420), .A2(n381), .ZN(n404) );
  INV_X2 U258 ( .A(n421), .ZN(n420) );
  MUX2_X1 U259 ( .A(n417), .B(n422), .S(n398), .Z(B[3]) );
  INV_X2 U260 ( .A(n423), .ZN(n417) );
  NAND2_X2 U261 ( .A1(n424), .A2(n389), .ZN(n423) );
  INV_X2 U262 ( .A(n408), .ZN(n424) );
  NAND2_X2 U263 ( .A1(n425), .A2(n381), .ZN(n408) );
  INV_X2 U264 ( .A(n426), .ZN(n425) );
  MUX2_X1 U265 ( .A(n427), .B(n428), .S(n398), .Z(B[31]) );
  MUX2_X1 U266 ( .A(n429), .B(n430), .S(n386), .Z(n427) );
  INV_X2 U267 ( .A(n431), .ZN(n430) );
  MUX2_X1 U268 ( .A(n432), .B(n433), .S(n379), .Z(n429) );
  INV_X2 U269 ( .A(n434), .ZN(n433) );
  MUX2_X1 U270 ( .A(n435), .B(n436), .S(n392), .Z(n432) );
  INV_X2 U271 ( .A(n437), .ZN(n436) );
  MUX2_X1 U272 ( .A(A[31]), .B(A[15]), .S(SH[4]), .Z(n435) );
  MUX2_X1 U273 ( .A(n428), .B(n438), .S(n398), .Z(B[30]) );
  INV_X2 U274 ( .A(n439), .ZN(n428) );
  MUX2_X1 U275 ( .A(n440), .B(n441), .S(n386), .Z(n439) );
  MUX2_X1 U276 ( .A(n442), .B(n443), .S(n379), .Z(n440) );
  MUX2_X1 U277 ( .A(n444), .B(n445), .S(n392), .Z(n442) );
  MUX2_X1 U278 ( .A(n446), .B(n447), .S(SH[4]), .Z(n444) );
  MUX2_X1 U279 ( .A(n422), .B(n448), .S(n398), .Z(B[2]) );
  INV_X2 U280 ( .A(n449), .ZN(n422) );
  NAND2_X2 U281 ( .A1(n450), .A2(n389), .ZN(n449) );
  INV_X2 U282 ( .A(n412), .ZN(n450) );
  NAND2_X2 U283 ( .A1(n451), .A2(n382), .ZN(n412) );
  INV_X2 U284 ( .A(n452), .ZN(n451) );
  MUX2_X1 U285 ( .A(n438), .B(n453), .S(n398), .Z(B[29]) );
  INV_X2 U286 ( .A(n454), .ZN(n438) );
  MUX2_X1 U287 ( .A(n455), .B(n456), .S(n386), .Z(n454) );
  MUX2_X1 U288 ( .A(n457), .B(n458), .S(n379), .Z(n455) );
  MUX2_X1 U289 ( .A(n437), .B(n459), .S(n392), .Z(n457) );
  MUX2_X1 U290 ( .A(n460), .B(n461), .S(SH[4]), .Z(n437) );
  MUX2_X1 U291 ( .A(n453), .B(n462), .S(n398), .Z(B[28]) );
  INV_X2 U292 ( .A(n463), .ZN(n453) );
  MUX2_X1 U293 ( .A(n464), .B(n465), .S(n386), .Z(n463) );
  MUX2_X1 U294 ( .A(n466), .B(n467), .S(n379), .Z(n464) );
  MUX2_X1 U295 ( .A(n445), .B(n468), .S(n392), .Z(n466) );
  MUX2_X1 U296 ( .A(n469), .B(n470), .S(SH[4]), .Z(n445) );
  MUX2_X1 U297 ( .A(n462), .B(n471), .S(n398), .Z(B[27]) );
  INV_X2 U298 ( .A(n472), .ZN(n462) );
  MUX2_X1 U299 ( .A(n431), .B(n473), .S(n386), .Z(n472) );
  MUX2_X1 U300 ( .A(n474), .B(n475), .S(n379), .Z(n431) );
  MUX2_X1 U301 ( .A(n459), .B(n476), .S(n392), .Z(n474) );
  MUX2_X1 U302 ( .A(n477), .B(n478), .S(SH[4]), .Z(n459) );
  MUX2_X1 U303 ( .A(n471), .B(n479), .S(n398), .Z(B[26]) );
  INV_X2 U304 ( .A(n480), .ZN(n471) );
  MUX2_X1 U305 ( .A(n441), .B(n481), .S(n386), .Z(n480) );
  MUX2_X1 U306 ( .A(n482), .B(n483), .S(n379), .Z(n441) );
  MUX2_X1 U307 ( .A(n468), .B(n484), .S(n392), .Z(n482) );
  MUX2_X1 U308 ( .A(n485), .B(n486), .S(SH[4]), .Z(n468) );
  MUX2_X1 U309 ( .A(n479), .B(n487), .S(n398), .Z(B[25]) );
  INV_X2 U310 ( .A(n488), .ZN(n479) );
  MUX2_X1 U311 ( .A(n456), .B(n489), .S(n386), .Z(n488) );
  MUX2_X1 U312 ( .A(n490), .B(n491), .S(n379), .Z(n456) );
  MUX2_X1 U313 ( .A(n476), .B(n492), .S(n392), .Z(n490) );
  MUX2_X1 U314 ( .A(n493), .B(n494), .S(SH[4]), .Z(n476) );
  MUX2_X1 U315 ( .A(n487), .B(n495), .S(n397), .Z(B[24]) );
  INV_X2 U316 ( .A(n496), .ZN(n487) );
  MUX2_X1 U317 ( .A(n465), .B(n497), .S(n387), .Z(n496) );
  MUX2_X1 U318 ( .A(n498), .B(n499), .S(n379), .Z(n465) );
  MUX2_X1 U319 ( .A(n484), .B(n500), .S(n392), .Z(n498) );
  MUX2_X1 U320 ( .A(n501), .B(n502), .S(SH[4]), .Z(n484) );
  MUX2_X1 U321 ( .A(n495), .B(n503), .S(n397), .Z(B[23]) );
  INV_X2 U322 ( .A(n504), .ZN(n495) );
  MUX2_X1 U323 ( .A(n473), .B(n505), .S(n387), .Z(n504) );
  MUX2_X1 U324 ( .A(n434), .B(n506), .S(n379), .Z(n473) );
  MUX2_X1 U325 ( .A(n492), .B(n507), .S(n392), .Z(n434) );
  MUX2_X1 U326 ( .A(n508), .B(n509), .S(SH[4]), .Z(n492) );
  MUX2_X1 U327 ( .A(n503), .B(n510), .S(n397), .Z(B[22]) );
  INV_X2 U328 ( .A(n511), .ZN(n503) );
  MUX2_X1 U329 ( .A(n481), .B(n512), .S(n387), .Z(n511) );
  MUX2_X1 U330 ( .A(n443), .B(n513), .S(n379), .Z(n481) );
  MUX2_X1 U331 ( .A(n500), .B(n514), .S(n392), .Z(n443) );
  MUX2_X1 U332 ( .A(n515), .B(n516), .S(SH[4]), .Z(n500) );
  MUX2_X1 U333 ( .A(n510), .B(n517), .S(n397), .Z(B[21]) );
  INV_X2 U334 ( .A(n518), .ZN(n510) );
  MUX2_X1 U335 ( .A(n489), .B(n519), .S(n387), .Z(n518) );
  MUX2_X1 U336 ( .A(n458), .B(n520), .S(n379), .Z(n489) );
  MUX2_X1 U337 ( .A(n507), .B(n521), .S(n392), .Z(n458) );
  MUX2_X1 U338 ( .A(n522), .B(n523), .S(SH[4]), .Z(n507) );
  MUX2_X1 U339 ( .A(n517), .B(n524), .S(n397), .Z(B[20]) );
  INV_X2 U340 ( .A(n525), .ZN(n517) );
  MUX2_X1 U341 ( .A(n497), .B(n526), .S(n387), .Z(n525) );
  MUX2_X1 U342 ( .A(n467), .B(n527), .S(n379), .Z(n497) );
  MUX2_X1 U343 ( .A(n514), .B(n528), .S(n392), .Z(n467) );
  MUX2_X1 U344 ( .A(n529), .B(n530), .S(SH[4]), .Z(n514) );
  MUX2_X1 U345 ( .A(n448), .B(n531), .S(n397), .Z(B[1]) );
  INV_X2 U346 ( .A(n532), .ZN(n531) );
  INV_X2 U347 ( .A(n533), .ZN(n448) );
  NAND2_X2 U348 ( .A1(n534), .A2(n390), .ZN(n533) );
  INV_X2 U349 ( .A(n416), .ZN(n534) );
  NAND2_X2 U350 ( .A1(n535), .A2(n382), .ZN(n416) );
  INV_X2 U351 ( .A(n536), .ZN(n535) );
  MUX2_X1 U352 ( .A(n524), .B(n537), .S(n397), .Z(B[19]) );
  INV_X2 U353 ( .A(n538), .ZN(n524) );
  MUX2_X1 U354 ( .A(n505), .B(n539), .S(n387), .Z(n538) );
  MUX2_X1 U355 ( .A(n475), .B(n540), .S(n380), .Z(n505) );
  MUX2_X1 U356 ( .A(n521), .B(n541), .S(n393), .Z(n475) );
  MUX2_X1 U357 ( .A(n542), .B(n543), .S(SH[4]), .Z(n521) );
  MUX2_X1 U358 ( .A(n537), .B(n544), .S(n397), .Z(B[18]) );
  INV_X2 U359 ( .A(n545), .ZN(n537) );
  MUX2_X1 U360 ( .A(n512), .B(n546), .S(n387), .Z(n545) );
  MUX2_X1 U361 ( .A(n483), .B(n547), .S(n380), .Z(n512) );
  MUX2_X1 U362 ( .A(n528), .B(n548), .S(n393), .Z(n483) );
  MUX2_X1 U363 ( .A(n549), .B(n550), .S(SH[4]), .Z(n528) );
  MUX2_X1 U364 ( .A(n544), .B(n551), .S(n397), .Z(B[17]) );
  INV_X2 U365 ( .A(n552), .ZN(n544) );
  MUX2_X1 U366 ( .A(n519), .B(n553), .S(n387), .Z(n552) );
  MUX2_X1 U367 ( .A(n491), .B(n554), .S(n380), .Z(n519) );
  MUX2_X1 U368 ( .A(n541), .B(n555), .S(n393), .Z(n491) );
  MUX2_X1 U369 ( .A(n556), .B(n557), .S(SH[4]), .Z(n541) );
  MUX2_X1 U370 ( .A(n551), .B(n558), .S(n397), .Z(B[16]) );
  INV_X2 U371 ( .A(n559), .ZN(n551) );
  MUX2_X1 U372 ( .A(n526), .B(n560), .S(n387), .Z(n559) );
  MUX2_X1 U373 ( .A(n499), .B(n561), .S(n380), .Z(n526) );
  MUX2_X1 U374 ( .A(n548), .B(n562), .S(n393), .Z(n499) );
  MUX2_X1 U375 ( .A(n563), .B(n564), .S(SH[4]), .Z(n548) );
  MUX2_X1 U376 ( .A(n558), .B(n565), .S(n397), .Z(B[15]) );
  INV_X2 U377 ( .A(n566), .ZN(n558) );
  MUX2_X1 U378 ( .A(n539), .B(n567), .S(n387), .Z(n566) );
  MUX2_X1 U379 ( .A(n506), .B(n568), .S(n380), .Z(n539) );
  MUX2_X1 U380 ( .A(n555), .B(n569), .S(n393), .Z(n506) );
  MUX2_X1 U381 ( .A(n565), .B(n570), .S(n397), .Z(B[14]) );
  INV_X2 U382 ( .A(n571), .ZN(n565) );
  MUX2_X1 U383 ( .A(n546), .B(n572), .S(n387), .Z(n571) );
  MUX2_X1 U384 ( .A(n513), .B(n573), .S(n380), .Z(n546) );
  MUX2_X1 U385 ( .A(n562), .B(n574), .S(n393), .Z(n513) );
  MUX2_X1 U386 ( .A(n570), .B(n575), .S(n397), .Z(B[13]) );
  INV_X2 U387 ( .A(n576), .ZN(n570) );
  MUX2_X1 U388 ( .A(n553), .B(n577), .S(n387), .Z(n576) );
  MUX2_X1 U389 ( .A(n520), .B(n578), .S(n380), .Z(n553) );
  MUX2_X1 U390 ( .A(n569), .B(n579), .S(n393), .Z(n520) );
  MUX2_X1 U391 ( .A(n575), .B(n580), .S(n397), .Z(B[12]) );
  INV_X2 U392 ( .A(n581), .ZN(n575) );
  MUX2_X1 U393 ( .A(n560), .B(n403), .S(n388), .Z(n581) );
  MUX2_X1 U394 ( .A(n561), .B(n582), .S(n380), .Z(n403) );
  MUX2_X1 U395 ( .A(n583), .B(n584), .S(n393), .Z(n561) );
  MUX2_X1 U396 ( .A(n527), .B(n421), .S(n380), .Z(n560) );
  MUX2_X1 U397 ( .A(n585), .B(n586), .S(n393), .Z(n421) );
  MUX2_X1 U398 ( .A(n574), .B(n587), .S(n393), .Z(n527) );
  MUX2_X1 U399 ( .A(n580), .B(n588), .S(n397), .Z(B[11]) );
  INV_X2 U400 ( .A(n589), .ZN(n580) );
  MUX2_X1 U401 ( .A(n567), .B(n407), .S(n388), .Z(n589) );
  NAND2_X2 U402 ( .A1(n590), .A2(n383), .ZN(n407) );
  INV_X2 U403 ( .A(n568), .ZN(n590) );
  MUX2_X1 U404 ( .A(n591), .B(n592), .S(n393), .Z(n568) );
  MUX2_X1 U405 ( .A(n540), .B(n426), .S(n380), .Z(n567) );
  MUX2_X1 U406 ( .A(n593), .B(n594), .S(n393), .Z(n426) );
  MUX2_X1 U407 ( .A(n579), .B(n595), .S(n394), .Z(n540) );
  MUX2_X1 U408 ( .A(n588), .B(n399), .S(n397), .Z(B[10]) );
  INV_X2 U409 ( .A(n596), .ZN(n399) );
  MUX2_X1 U410 ( .A(n577), .B(n415), .S(n388), .Z(n596) );
  NAND2_X2 U411 ( .A1(n597), .A2(n383), .ZN(n415) );
  INV_X2 U412 ( .A(n578), .ZN(n597) );
  MUX2_X1 U413 ( .A(n592), .B(n593), .S(n394), .Z(n578) );
  MUX2_X1 U414 ( .A(n554), .B(n536), .S(n380), .Z(n577) );
  NAND2_X2 U415 ( .A1(n598), .A2(n395), .ZN(n536) );
  INV_X2 U416 ( .A(n594), .ZN(n598) );
  MUX2_X1 U417 ( .A(n595), .B(n591), .S(n394), .Z(n554) );
  INV_X2 U418 ( .A(n599), .ZN(n588) );
  MUX2_X1 U419 ( .A(n572), .B(n411), .S(n388), .Z(n599) );
  NAND2_X2 U420 ( .A1(n600), .A2(n384), .ZN(n411) );
  INV_X2 U421 ( .A(n573), .ZN(n600) );
  MUX2_X1 U422 ( .A(n584), .B(n585), .S(n394), .Z(n573) );
  MUX2_X1 U423 ( .A(n547), .B(n452), .S(n380), .Z(n572) );
  MUX2_X1 U424 ( .A(n586), .B(n601), .S(n394), .Z(n452) );
  MUX2_X1 U425 ( .A(n587), .B(n583), .S(n394), .Z(n547) );
  NOR2_X2 U426 ( .A1(n397), .A2(n532), .ZN(B[0]) );
  NAND2_X2 U427 ( .A1(n602), .A2(n390), .ZN(n532) );
  INV_X2 U428 ( .A(n419), .ZN(n602) );
  NAND2_X2 U429 ( .A1(n603), .A2(n384), .ZN(n419) );
  INV_X2 U430 ( .A(n582), .ZN(n603) );
  NAND2_X2 U431 ( .A1(n604), .A2(n395), .ZN(n582) );
  INV_X2 U432 ( .A(n601), .ZN(n604) );
endmodule


module up_island_DW01_bsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408;

  INV_X1 U163 ( .A(A[18]), .ZN(n402) );
  INV_X1 U164 ( .A(A[15]), .ZN(n343) );
  INV_X1 U165 ( .A(A[19]), .ZN(n383) );
  INV_X1 U166 ( .A(A[20]), .ZN(n397) );
  INV_X1 U167 ( .A(A[21]), .ZN(n385) );
  INV_X1 U168 ( .A(A[9]), .ZN(n391) );
  INV_X1 U169 ( .A(A[10]), .ZN(n405) );
  INV_X1 U170 ( .A(A[22]), .ZN(n399) );
  INV_X1 U171 ( .A(A[23]), .ZN(n390) );
  INV_X1 U172 ( .A(A[8]), .ZN(n403) );
  INV_X1 U173 ( .A(A[16]), .ZN(n336) );
  INV_X1 U174 ( .A(A[17]), .ZN(n388) );
  INV_X1 U175 ( .A(A[28]), .ZN(n368) );
  INV_X1 U176 ( .A(A[27]), .ZN(n378) );
  INV_X1 U177 ( .A(A[25]), .ZN(n392) );
  INV_X1 U178 ( .A(A[30]), .ZN(n351) );
  INV_X1 U179 ( .A(A[7]), .ZN(n389) );
  INV_X1 U180 ( .A(A[14]), .ZN(n350) );
  INV_X1 U181 ( .A(A[13]), .ZN(n357) );
  INV_X1 U182 ( .A(A[11]), .ZN(n377) );
  INV_X1 U183 ( .A(A[12]), .ZN(n367) );
  INV_X1 U184 ( .A(A[29]), .ZN(n358) );
  INV_X1 U185 ( .A(A[5]), .ZN(n384) );
  INV_X1 U186 ( .A(A[26]), .ZN(n406) );
  INV_X1 U187 ( .A(A[24]), .ZN(n404) );
  INV_X1 U188 ( .A(A[6]), .ZN(n398) );
  INV_X1 U189 ( .A(A[4]), .ZN(n396) );
  INV_X1 U190 ( .A(A[3]), .ZN(n382) );
  INV_X1 U191 ( .A(A[2]), .ZN(n401) );
  INV_X1 U192 ( .A(A[0]), .ZN(n337) );
  INV_X1 U193 ( .A(A[1]), .ZN(n387) );
  BUF_X1 U194 ( .A(SH[4]), .Z(n202) );
  BUF_X1 U195 ( .A(SH[4]), .Z(n203) );
  BUF_X1 U196 ( .A(SH[4]), .Z(n204) );
  BUF_X1 U197 ( .A(SH[3]), .Z(n205) );
  BUF_X1 U198 ( .A(SH[3]), .Z(n206) );
  BUF_X1 U199 ( .A(SH[3]), .Z(n207) );
  BUF_X1 U200 ( .A(SH[2]), .Z(n208) );
  BUF_X1 U201 ( .A(SH[2]), .Z(n209) );
  BUF_X1 U202 ( .A(SH[2]), .Z(n210) );
  BUF_X1 U203 ( .A(SH[1]), .Z(n211) );
  BUF_X1 U204 ( .A(SH[1]), .Z(n212) );
  BUF_X1 U205 ( .A(SH[1]), .Z(n213) );
  BUF_X1 U206 ( .A(SH[0]), .Z(n214) );
  BUF_X1 U207 ( .A(SH[0]), .Z(n215) );
  BUF_X1 U208 ( .A(SH[0]), .Z(n216) );
  MUX2_X1 U209 ( .A(n217), .B(n218), .S(n214), .Z(B[9]) );
  MUX2_X1 U210 ( .A(n218), .B(n219), .S(n214), .Z(B[8]) );
  INV_X2 U211 ( .A(n220), .ZN(n218) );
  MUX2_X1 U212 ( .A(n221), .B(n222), .S(n208), .Z(n220) );
  MUX2_X1 U213 ( .A(n219), .B(n223), .S(n214), .Z(B[7]) );
  INV_X2 U214 ( .A(n224), .ZN(n219) );
  MUX2_X1 U215 ( .A(n225), .B(n226), .S(n208), .Z(n224) );
  MUX2_X1 U216 ( .A(n223), .B(n227), .S(n214), .Z(B[6]) );
  INV_X2 U217 ( .A(n228), .ZN(n223) );
  MUX2_X1 U218 ( .A(n229), .B(n230), .S(n208), .Z(n228) );
  MUX2_X1 U219 ( .A(n227), .B(n231), .S(n214), .Z(B[5]) );
  INV_X2 U220 ( .A(n232), .ZN(n227) );
  MUX2_X1 U221 ( .A(n233), .B(n234), .S(n208), .Z(n232) );
  MUX2_X1 U222 ( .A(n231), .B(n235), .S(n214), .Z(B[4]) );
  INV_X2 U223 ( .A(n236), .ZN(n231) );
  MUX2_X1 U224 ( .A(n222), .B(n237), .S(n208), .Z(n236) );
  MUX2_X1 U225 ( .A(n238), .B(n239), .S(n205), .Z(n222) );
  MUX2_X1 U226 ( .A(n235), .B(n240), .S(n214), .Z(B[3]) );
  INV_X2 U227 ( .A(n241), .ZN(n235) );
  MUX2_X1 U228 ( .A(n226), .B(n242), .S(n208), .Z(n241) );
  MUX2_X1 U229 ( .A(n243), .B(n244), .S(n205), .Z(n226) );
  MUX2_X1 U230 ( .A(n245), .B(n246), .S(n214), .Z(B[31]) );
  MUX2_X1 U231 ( .A(n246), .B(n247), .S(n214), .Z(B[30]) );
  INV_X2 U232 ( .A(n248), .ZN(n246) );
  MUX2_X1 U233 ( .A(n249), .B(n250), .S(n208), .Z(n248) );
  MUX2_X1 U234 ( .A(n240), .B(n251), .S(n214), .Z(B[2]) );
  INV_X2 U235 ( .A(n252), .ZN(n240) );
  MUX2_X1 U236 ( .A(n230), .B(n249), .S(n208), .Z(n252) );
  MUX2_X1 U237 ( .A(n253), .B(n254), .S(n205), .Z(n249) );
  MUX2_X1 U238 ( .A(n255), .B(n256), .S(n205), .Z(n230) );
  MUX2_X1 U239 ( .A(n247), .B(n257), .S(n214), .Z(B[29]) );
  INV_X2 U240 ( .A(n258), .ZN(n247) );
  MUX2_X1 U241 ( .A(n259), .B(n260), .S(n208), .Z(n258) );
  MUX2_X1 U242 ( .A(n257), .B(n261), .S(n214), .Z(B[28]) );
  INV_X2 U243 ( .A(n262), .ZN(n257) );
  MUX2_X1 U244 ( .A(n263), .B(n264), .S(n208), .Z(n262) );
  MUX2_X1 U245 ( .A(n261), .B(n265), .S(n215), .Z(B[27]) );
  INV_X2 U246 ( .A(n266), .ZN(n261) );
  MUX2_X1 U247 ( .A(n267), .B(n268), .S(n208), .Z(n266) );
  MUX2_X1 U248 ( .A(n265), .B(n269), .S(n215), .Z(B[26]) );
  INV_X2 U249 ( .A(n270), .ZN(n265) );
  MUX2_X1 U250 ( .A(n250), .B(n271), .S(n208), .Z(n270) );
  MUX2_X1 U251 ( .A(n256), .B(n272), .S(n205), .Z(n250) );
  MUX2_X1 U252 ( .A(n273), .B(n274), .S(n211), .Z(n256) );
  MUX2_X1 U253 ( .A(n269), .B(n275), .S(n215), .Z(B[25]) );
  INV_X2 U254 ( .A(n276), .ZN(n269) );
  MUX2_X1 U255 ( .A(n260), .B(n277), .S(n209), .Z(n276) );
  MUX2_X1 U256 ( .A(n278), .B(n279), .S(n205), .Z(n260) );
  MUX2_X1 U257 ( .A(n275), .B(n280), .S(n215), .Z(B[24]) );
  INV_X2 U258 ( .A(n281), .ZN(n275) );
  MUX2_X1 U259 ( .A(n264), .B(n282), .S(n209), .Z(n281) );
  MUX2_X1 U260 ( .A(n283), .B(n284), .S(n205), .Z(n264) );
  MUX2_X1 U261 ( .A(n280), .B(n285), .S(n215), .Z(B[23]) );
  INV_X2 U262 ( .A(n286), .ZN(n280) );
  MUX2_X1 U263 ( .A(n268), .B(n287), .S(n209), .Z(n286) );
  MUX2_X1 U264 ( .A(n288), .B(n289), .S(n205), .Z(n268) );
  MUX2_X1 U265 ( .A(n285), .B(n290), .S(n215), .Z(B[22]) );
  INV_X2 U266 ( .A(n291), .ZN(n285) );
  MUX2_X1 U267 ( .A(n271), .B(n292), .S(n209), .Z(n291) );
  MUX2_X1 U268 ( .A(n254), .B(n293), .S(n205), .Z(n271) );
  MUX2_X1 U269 ( .A(n294), .B(n295), .S(n211), .Z(n254) );
  MUX2_X1 U270 ( .A(n290), .B(n296), .S(n215), .Z(B[21]) );
  INV_X2 U271 ( .A(n297), .ZN(n290) );
  MUX2_X1 U272 ( .A(n277), .B(n298), .S(n209), .Z(n297) );
  MUX2_X1 U273 ( .A(n299), .B(n300), .S(n205), .Z(n277) );
  MUX2_X1 U274 ( .A(n296), .B(n301), .S(n215), .Z(B[20]) );
  INV_X2 U275 ( .A(n302), .ZN(n296) );
  MUX2_X1 U276 ( .A(n282), .B(n303), .S(n209), .Z(n302) );
  MUX2_X1 U277 ( .A(n304), .B(n305), .S(n205), .Z(n282) );
  MUX2_X1 U278 ( .A(n251), .B(n306), .S(n215), .Z(B[1]) );
  INV_X2 U279 ( .A(n307), .ZN(n251) );
  MUX2_X1 U280 ( .A(n234), .B(n259), .S(n209), .Z(n307) );
  MUX2_X1 U281 ( .A(n308), .B(n299), .S(n205), .Z(n259) );
  MUX2_X1 U282 ( .A(n309), .B(n310), .S(n211), .Z(n299) );
  MUX2_X1 U283 ( .A(n311), .B(n278), .S(n206), .Z(n234) );
  MUX2_X1 U284 ( .A(n312), .B(n313), .S(n211), .Z(n278) );
  MUX2_X1 U285 ( .A(n301), .B(n314), .S(n215), .Z(B[19]) );
  INV_X2 U286 ( .A(n315), .ZN(n301) );
  MUX2_X1 U287 ( .A(n287), .B(n316), .S(n209), .Z(n315) );
  MUX2_X1 U288 ( .A(n317), .B(n318), .S(n206), .Z(n287) );
  MUX2_X1 U289 ( .A(n314), .B(n319), .S(n215), .Z(B[18]) );
  INV_X2 U290 ( .A(n320), .ZN(n314) );
  MUX2_X1 U291 ( .A(n292), .B(n321), .S(n209), .Z(n320) );
  MUX2_X1 U292 ( .A(n272), .B(n322), .S(n206), .Z(n292) );
  MUX2_X1 U293 ( .A(n323), .B(n324), .S(n211), .Z(n272) );
  MUX2_X1 U294 ( .A(n319), .B(n325), .S(n215), .Z(B[17]) );
  INV_X2 U295 ( .A(n326), .ZN(n319) );
  MUX2_X1 U296 ( .A(n298), .B(n327), .S(n209), .Z(n326) );
  MUX2_X1 U297 ( .A(n279), .B(n328), .S(n206), .Z(n298) );
  MUX2_X1 U298 ( .A(n329), .B(n330), .S(n211), .Z(n279) );
  MUX2_X1 U299 ( .A(n325), .B(n331), .S(n216), .Z(B[16]) );
  INV_X2 U300 ( .A(n332), .ZN(n325) );
  MUX2_X1 U301 ( .A(n303), .B(n333), .S(n209), .Z(n332) );
  MUX2_X1 U302 ( .A(n284), .B(n334), .S(n206), .Z(n303) );
  MUX2_X1 U303 ( .A(n324), .B(n335), .S(n211), .Z(n284) );
  MUX2_X1 U304 ( .A(n336), .B(n337), .S(n202), .Z(n324) );
  MUX2_X1 U305 ( .A(n331), .B(n338), .S(n216), .Z(B[15]) );
  INV_X2 U306 ( .A(n339), .ZN(n331) );
  MUX2_X1 U307 ( .A(n316), .B(n340), .S(n209), .Z(n339) );
  MUX2_X1 U308 ( .A(n289), .B(n341), .S(n206), .Z(n316) );
  MUX2_X1 U309 ( .A(n330), .B(n342), .S(n211), .Z(n289) );
  MUX2_X1 U310 ( .A(n343), .B(n344), .S(n202), .Z(n330) );
  MUX2_X1 U311 ( .A(n338), .B(n345), .S(n216), .Z(B[14]) );
  INV_X2 U312 ( .A(n346), .ZN(n338) );
  MUX2_X1 U313 ( .A(n321), .B(n347), .S(n210), .Z(n346) );
  MUX2_X1 U314 ( .A(n293), .B(n348), .S(n206), .Z(n321) );
  MUX2_X1 U315 ( .A(n335), .B(n349), .S(n211), .Z(n293) );
  MUX2_X1 U316 ( .A(n350), .B(n351), .S(n202), .Z(n335) );
  MUX2_X1 U317 ( .A(n345), .B(n352), .S(n216), .Z(B[13]) );
  INV_X2 U318 ( .A(n353), .ZN(n345) );
  MUX2_X1 U319 ( .A(n327), .B(n354), .S(n210), .Z(n353) );
  MUX2_X1 U320 ( .A(n300), .B(n355), .S(n206), .Z(n327) );
  MUX2_X1 U321 ( .A(n342), .B(n356), .S(n211), .Z(n300) );
  MUX2_X1 U322 ( .A(n357), .B(n358), .S(n202), .Z(n342) );
  MUX2_X1 U323 ( .A(n352), .B(n359), .S(n216), .Z(B[12]) );
  INV_X2 U324 ( .A(n360), .ZN(n352) );
  MUX2_X1 U325 ( .A(n333), .B(n221), .S(n210), .Z(n360) );
  MUX2_X1 U326 ( .A(n334), .B(n361), .S(n206), .Z(n221) );
  MUX2_X1 U327 ( .A(n362), .B(n363), .S(n211), .Z(n334) );
  MUX2_X1 U328 ( .A(n305), .B(n238), .S(n206), .Z(n333) );
  MUX2_X1 U329 ( .A(n364), .B(n365), .S(n211), .Z(n238) );
  MUX2_X1 U330 ( .A(n349), .B(n366), .S(n212), .Z(n305) );
  MUX2_X1 U331 ( .A(n367), .B(n368), .S(n202), .Z(n349) );
  MUX2_X1 U332 ( .A(n359), .B(n369), .S(n216), .Z(B[11]) );
  INV_X2 U333 ( .A(n370), .ZN(n359) );
  MUX2_X1 U334 ( .A(n340), .B(n225), .S(n210), .Z(n370) );
  MUX2_X1 U335 ( .A(n341), .B(n371), .S(n206), .Z(n225) );
  MUX2_X1 U336 ( .A(n372), .B(n373), .S(n212), .Z(n341) );
  MUX2_X1 U337 ( .A(n318), .B(n243), .S(n206), .Z(n340) );
  MUX2_X1 U338 ( .A(n374), .B(n375), .S(n212), .Z(n243) );
  MUX2_X1 U339 ( .A(n356), .B(n376), .S(n212), .Z(n318) );
  MUX2_X1 U340 ( .A(n377), .B(n378), .S(n202), .Z(n356) );
  MUX2_X1 U341 ( .A(n369), .B(n217), .S(n216), .Z(B[10]) );
  INV_X2 U342 ( .A(n379), .ZN(n217) );
  MUX2_X1 U343 ( .A(n354), .B(n233), .S(n210), .Z(n379) );
  MUX2_X1 U344 ( .A(n355), .B(n308), .S(n207), .Z(n233) );
  MUX2_X1 U345 ( .A(n380), .B(n381), .S(n212), .Z(n308) );
  MUX2_X1 U346 ( .A(n373), .B(n374), .S(n212), .Z(n355) );
  MUX2_X1 U347 ( .A(n382), .B(n383), .S(n202), .Z(n374) );
  MUX2_X1 U348 ( .A(n384), .B(n385), .S(n202), .Z(n373) );
  MUX2_X1 U349 ( .A(n328), .B(n311), .S(n207), .Z(n354) );
  MUX2_X1 U350 ( .A(n375), .B(n386), .S(n212), .Z(n311) );
  MUX2_X1 U351 ( .A(n387), .B(n388), .S(n202), .Z(n375) );
  MUX2_X1 U352 ( .A(n376), .B(n372), .S(n212), .Z(n328) );
  MUX2_X1 U353 ( .A(n389), .B(n390), .S(n202), .Z(n372) );
  MUX2_X1 U354 ( .A(n391), .B(n392), .S(n202), .Z(n376) );
  INV_X2 U355 ( .A(n393), .ZN(n369) );
  MUX2_X1 U356 ( .A(n347), .B(n229), .S(n210), .Z(n393) );
  MUX2_X1 U357 ( .A(n348), .B(n253), .S(n207), .Z(n229) );
  MUX2_X1 U358 ( .A(n394), .B(n395), .S(n212), .Z(n253) );
  MUX2_X1 U359 ( .A(n363), .B(n364), .S(n212), .Z(n348) );
  MUX2_X1 U360 ( .A(n396), .B(n397), .S(n202), .Z(n364) );
  MUX2_X1 U361 ( .A(n398), .B(n399), .S(n203), .Z(n363) );
  MUX2_X1 U362 ( .A(n322), .B(n255), .S(n207), .Z(n347) );
  MUX2_X1 U363 ( .A(n365), .B(n400), .S(n212), .Z(n255) );
  MUX2_X1 U364 ( .A(n401), .B(n402), .S(n203), .Z(n365) );
  MUX2_X1 U365 ( .A(n366), .B(n362), .S(n212), .Z(n322) );
  MUX2_X1 U366 ( .A(n403), .B(n404), .S(n203), .Z(n362) );
  MUX2_X1 U367 ( .A(n405), .B(n406), .S(n203), .Z(n366) );
  MUX2_X1 U368 ( .A(n306), .B(n245), .S(n216), .Z(B[0]) );
  INV_X2 U369 ( .A(n407), .ZN(n245) );
  MUX2_X1 U370 ( .A(n242), .B(n267), .S(n210), .Z(n407) );
  MUX2_X1 U371 ( .A(n244), .B(n317), .S(n207), .Z(n267) );
  MUX2_X1 U372 ( .A(n310), .B(n329), .S(n213), .Z(n317) );
  MUX2_X1 U373 ( .A(n388), .B(n387), .S(n203), .Z(n329) );
  MUX2_X1 U374 ( .A(n383), .B(n382), .S(n203), .Z(n310) );
  MUX2_X1 U375 ( .A(n381), .B(n312), .S(n213), .Z(n244) );
  MUX2_X1 U376 ( .A(n392), .B(n391), .S(n203), .Z(n312) );
  MUX2_X1 U377 ( .A(n378), .B(n377), .S(n203), .Z(n381) );
  MUX2_X1 U378 ( .A(n371), .B(n288), .S(n207), .Z(n242) );
  MUX2_X1 U379 ( .A(n313), .B(n309), .S(n213), .Z(n288) );
  MUX2_X1 U380 ( .A(n385), .B(n384), .S(n203), .Z(n309) );
  MUX2_X1 U381 ( .A(n390), .B(n389), .S(n203), .Z(n313) );
  MUX2_X1 U382 ( .A(n386), .B(n380), .S(n213), .Z(n371) );
  MUX2_X1 U383 ( .A(n358), .B(n357), .S(n203), .Z(n380) );
  MUX2_X1 U384 ( .A(n344), .B(n343), .S(n203), .Z(n386) );
  INV_X2 U385 ( .A(A[31]), .ZN(n344) );
  INV_X2 U386 ( .A(n408), .ZN(n306) );
  MUX2_X1 U387 ( .A(n237), .B(n263), .S(n210), .Z(n408) );
  MUX2_X1 U388 ( .A(n239), .B(n304), .S(n207), .Z(n263) );
  MUX2_X1 U389 ( .A(n295), .B(n323), .S(n213), .Z(n304) );
  MUX2_X1 U390 ( .A(n402), .B(n401), .S(n204), .Z(n323) );
  MUX2_X1 U391 ( .A(n397), .B(n396), .S(n204), .Z(n295) );
  MUX2_X1 U392 ( .A(n395), .B(n273), .S(n213), .Z(n239) );
  MUX2_X1 U393 ( .A(n406), .B(n405), .S(n204), .Z(n273) );
  MUX2_X1 U394 ( .A(n368), .B(n367), .S(n204), .Z(n395) );
  MUX2_X1 U395 ( .A(n361), .B(n283), .S(n207), .Z(n237) );
  MUX2_X1 U396 ( .A(n274), .B(n294), .S(n213), .Z(n283) );
  MUX2_X1 U397 ( .A(n399), .B(n398), .S(n204), .Z(n294) );
  MUX2_X1 U398 ( .A(n404), .B(n403), .S(n204), .Z(n274) );
  MUX2_X1 U399 ( .A(n400), .B(n394), .S(n213), .Z(n361) );
  MUX2_X1 U400 ( .A(n351), .B(n350), .S(n204), .Z(n394) );
  MUX2_X1 U401 ( .A(n337), .B(n336), .S(n204), .Z(n400) );
endmodule


module up_island_DW_rbsh_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409;

  INV_X1 U164 ( .A(A[18]), .ZN(n404) );
  INV_X1 U165 ( .A(A[15]), .ZN(n338) );
  INV_X1 U166 ( .A(A[19]), .ZN(n390) );
  INV_X1 U167 ( .A(A[20]), .ZN(n402) );
  INV_X1 U168 ( .A(A[21]), .ZN(n388) );
  INV_X1 U169 ( .A(A[9]), .ZN(n382) );
  INV_X1 U170 ( .A(A[10]), .ZN(n374) );
  INV_X1 U171 ( .A(A[22]), .ZN(n397) );
  INV_X1 U172 ( .A(A[23]), .ZN(n383) );
  INV_X1 U173 ( .A(A[8]), .ZN(n396) );
  INV_X1 U174 ( .A(A[16]), .ZN(n400) );
  INV_X1 U175 ( .A(A[17]), .ZN(n386) );
  INV_X1 U176 ( .A(A[28]), .ZN(n358) );
  INV_X1 U177 ( .A(A[27]), .ZN(n363) );
  INV_X1 U178 ( .A(A[25]), .ZN(n381) );
  INV_X1 U179 ( .A(A[30]), .ZN(n344) );
  INV_X1 U180 ( .A(A[7]), .ZN(n384) );
  INV_X1 U181 ( .A(A[14]), .ZN(n345) );
  INV_X1 U182 ( .A(A[13]), .ZN(n352) );
  INV_X1 U183 ( .A(A[11]), .ZN(n364) );
  INV_X1 U184 ( .A(A[12]), .ZN(n359) );
  INV_X1 U185 ( .A(A[29]), .ZN(n351) );
  INV_X1 U186 ( .A(A[5]), .ZN(n389) );
  INV_X1 U187 ( .A(A[26]), .ZN(n373) );
  INV_X1 U188 ( .A(A[24]), .ZN(n395) );
  INV_X1 U189 ( .A(A[6]), .ZN(n398) );
  INV_X1 U190 ( .A(A[4]), .ZN(n403) );
  INV_X1 U191 ( .A(A[3]), .ZN(n391) );
  INV_X1 U192 ( .A(A[2]), .ZN(n405) );
  INV_X1 U193 ( .A(A[0]), .ZN(n401) );
  INV_X1 U194 ( .A(A[1]), .ZN(n387) );
  BUF_X1 U195 ( .A(SH[4]), .Z(n203) );
  BUF_X1 U196 ( .A(SH[4]), .Z(n204) );
  BUF_X1 U197 ( .A(SH[4]), .Z(n205) );
  BUF_X1 U198 ( .A(SH[3]), .Z(n206) );
  BUF_X1 U199 ( .A(SH[3]), .Z(n207) );
  BUF_X1 U200 ( .A(SH[3]), .Z(n208) );
  BUF_X1 U201 ( .A(SH[2]), .Z(n209) );
  BUF_X1 U202 ( .A(SH[2]), .Z(n210) );
  BUF_X1 U203 ( .A(SH[2]), .Z(n211) );
  BUF_X1 U204 ( .A(SH[1]), .Z(n212) );
  BUF_X1 U205 ( .A(SH[1]), .Z(n213) );
  BUF_X1 U206 ( .A(SH[1]), .Z(n214) );
  BUF_X1 U207 ( .A(SH[0]), .Z(n215) );
  BUF_X1 U208 ( .A(SH[0]), .Z(n216) );
  BUF_X1 U209 ( .A(SH[0]), .Z(n217) );
  MUX2_X1 U210 ( .A(n218), .B(n219), .S(n215), .Z(B[9]) );
  MUX2_X1 U211 ( .A(n220), .B(n218), .S(n215), .Z(B[8]) );
  INV_X2 U212 ( .A(n221), .ZN(n218) );
  MUX2_X1 U213 ( .A(n222), .B(n223), .S(n209), .Z(n221) );
  MUX2_X1 U214 ( .A(n224), .B(n220), .S(n215), .Z(B[7]) );
  INV_X2 U215 ( .A(n225), .ZN(n220) );
  MUX2_X1 U216 ( .A(n226), .B(n227), .S(n209), .Z(n225) );
  MUX2_X1 U217 ( .A(n228), .B(n224), .S(n215), .Z(B[6]) );
  INV_X2 U218 ( .A(n229), .ZN(n224) );
  MUX2_X1 U219 ( .A(n230), .B(n231), .S(n209), .Z(n229) );
  MUX2_X1 U220 ( .A(n232), .B(n228), .S(n215), .Z(B[5]) );
  INV_X2 U221 ( .A(n233), .ZN(n228) );
  MUX2_X1 U222 ( .A(n234), .B(n235), .S(n209), .Z(n233) );
  MUX2_X1 U223 ( .A(n236), .B(n232), .S(n215), .Z(B[4]) );
  INV_X2 U224 ( .A(n237), .ZN(n232) );
  MUX2_X1 U225 ( .A(n238), .B(n222), .S(n209), .Z(n237) );
  MUX2_X1 U226 ( .A(n239), .B(n240), .S(n206), .Z(n222) );
  MUX2_X1 U227 ( .A(n241), .B(n236), .S(n215), .Z(B[3]) );
  INV_X2 U228 ( .A(n242), .ZN(n236) );
  MUX2_X1 U229 ( .A(n243), .B(n226), .S(n209), .Z(n242) );
  MUX2_X1 U230 ( .A(n244), .B(n245), .S(n206), .Z(n226) );
  MUX2_X1 U231 ( .A(n246), .B(n247), .S(n215), .Z(B[31]) );
  MUX2_X1 U232 ( .A(n248), .B(n246), .S(n215), .Z(B[30]) );
  INV_X2 U233 ( .A(n249), .ZN(n246) );
  MUX2_X1 U234 ( .A(n250), .B(n251), .S(n209), .Z(n249) );
  MUX2_X1 U235 ( .A(n252), .B(n241), .S(n215), .Z(B[2]) );
  INV_X2 U236 ( .A(n253), .ZN(n241) );
  MUX2_X1 U237 ( .A(n251), .B(n230), .S(n209), .Z(n253) );
  MUX2_X1 U238 ( .A(n254), .B(n255), .S(n206), .Z(n230) );
  MUX2_X1 U239 ( .A(n256), .B(n257), .S(n206), .Z(n251) );
  MUX2_X1 U240 ( .A(n258), .B(n248), .S(n215), .Z(B[29]) );
  INV_X2 U241 ( .A(n259), .ZN(n248) );
  MUX2_X1 U242 ( .A(n260), .B(n261), .S(n209), .Z(n259) );
  MUX2_X1 U243 ( .A(n262), .B(n258), .S(n215), .Z(B[28]) );
  INV_X2 U244 ( .A(n263), .ZN(n258) );
  MUX2_X1 U245 ( .A(n264), .B(n265), .S(n209), .Z(n263) );
  MUX2_X1 U246 ( .A(n266), .B(n262), .S(n216), .Z(B[27]) );
  INV_X2 U247 ( .A(n267), .ZN(n262) );
  MUX2_X1 U248 ( .A(n268), .B(n269), .S(n209), .Z(n267) );
  MUX2_X1 U249 ( .A(n270), .B(n266), .S(n216), .Z(B[26]) );
  INV_X2 U250 ( .A(n271), .ZN(n266) );
  MUX2_X1 U251 ( .A(n272), .B(n250), .S(n209), .Z(n271) );
  MUX2_X1 U252 ( .A(n273), .B(n254), .S(n206), .Z(n250) );
  MUX2_X1 U253 ( .A(n274), .B(n275), .S(n212), .Z(n254) );
  MUX2_X1 U254 ( .A(n276), .B(n270), .S(n216), .Z(B[25]) );
  INV_X2 U255 ( .A(n277), .ZN(n270) );
  MUX2_X1 U256 ( .A(n278), .B(n260), .S(n210), .Z(n277) );
  MUX2_X1 U257 ( .A(n279), .B(n280), .S(n206), .Z(n260) );
  MUX2_X1 U258 ( .A(n281), .B(n276), .S(n216), .Z(B[24]) );
  INV_X2 U259 ( .A(n282), .ZN(n276) );
  MUX2_X1 U260 ( .A(n283), .B(n264), .S(n210), .Z(n282) );
  MUX2_X1 U261 ( .A(n284), .B(n285), .S(n206), .Z(n264) );
  MUX2_X1 U262 ( .A(n286), .B(n281), .S(n216), .Z(B[23]) );
  INV_X2 U263 ( .A(n287), .ZN(n281) );
  MUX2_X1 U264 ( .A(n288), .B(n268), .S(n210), .Z(n287) );
  MUX2_X1 U265 ( .A(n289), .B(n290), .S(n206), .Z(n268) );
  MUX2_X1 U266 ( .A(n291), .B(n286), .S(n216), .Z(B[22]) );
  INV_X2 U267 ( .A(n292), .ZN(n286) );
  MUX2_X1 U268 ( .A(n293), .B(n272), .S(n210), .Z(n292) );
  MUX2_X1 U269 ( .A(n294), .B(n256), .S(n206), .Z(n272) );
  MUX2_X1 U270 ( .A(n295), .B(n296), .S(n212), .Z(n256) );
  MUX2_X1 U271 ( .A(n297), .B(n291), .S(n216), .Z(B[21]) );
  INV_X2 U272 ( .A(n298), .ZN(n291) );
  MUX2_X1 U273 ( .A(n299), .B(n278), .S(n210), .Z(n298) );
  MUX2_X1 U274 ( .A(n300), .B(n301), .S(n206), .Z(n278) );
  MUX2_X1 U275 ( .A(n302), .B(n297), .S(n216), .Z(B[20]) );
  INV_X2 U276 ( .A(n303), .ZN(n297) );
  MUX2_X1 U277 ( .A(n304), .B(n283), .S(n210), .Z(n303) );
  MUX2_X1 U278 ( .A(n305), .B(n306), .S(n206), .Z(n283) );
  MUX2_X1 U279 ( .A(n307), .B(n252), .S(n216), .Z(B[1]) );
  INV_X2 U280 ( .A(n308), .ZN(n252) );
  MUX2_X1 U281 ( .A(n261), .B(n234), .S(n210), .Z(n308) );
  MUX2_X1 U282 ( .A(n280), .B(n309), .S(n206), .Z(n234) );
  MUX2_X1 U283 ( .A(n310), .B(n311), .S(n212), .Z(n280) );
  MUX2_X1 U284 ( .A(n301), .B(n312), .S(n207), .Z(n261) );
  MUX2_X1 U285 ( .A(n313), .B(n314), .S(n212), .Z(n301) );
  MUX2_X1 U286 ( .A(n315), .B(n302), .S(n216), .Z(B[19]) );
  INV_X2 U287 ( .A(n316), .ZN(n302) );
  MUX2_X1 U288 ( .A(n317), .B(n288), .S(n210), .Z(n316) );
  MUX2_X1 U289 ( .A(n318), .B(n319), .S(n207), .Z(n288) );
  MUX2_X1 U290 ( .A(n320), .B(n315), .S(n216), .Z(B[18]) );
  INV_X2 U291 ( .A(n321), .ZN(n315) );
  MUX2_X1 U292 ( .A(n322), .B(n293), .S(n210), .Z(n321) );
  MUX2_X1 U293 ( .A(n323), .B(n273), .S(n207), .Z(n293) );
  MUX2_X1 U294 ( .A(n324), .B(n325), .S(n212), .Z(n273) );
  MUX2_X1 U295 ( .A(n326), .B(n320), .S(n216), .Z(B[17]) );
  INV_X2 U296 ( .A(n327), .ZN(n320) );
  MUX2_X1 U297 ( .A(n328), .B(n299), .S(n210), .Z(n327) );
  MUX2_X1 U298 ( .A(n329), .B(n279), .S(n207), .Z(n299) );
  MUX2_X1 U299 ( .A(n330), .B(n331), .S(n212), .Z(n279) );
  MUX2_X1 U300 ( .A(n332), .B(n326), .S(n217), .Z(B[16]) );
  INV_X2 U301 ( .A(n333), .ZN(n326) );
  MUX2_X1 U302 ( .A(n334), .B(n304), .S(n210), .Z(n333) );
  MUX2_X1 U303 ( .A(n335), .B(n284), .S(n207), .Z(n304) );
  MUX2_X1 U304 ( .A(n336), .B(n324), .S(n212), .Z(n284) );
  MUX2_X1 U305 ( .A(n337), .B(n338), .S(n203), .Z(n324) );
  MUX2_X1 U306 ( .A(n339), .B(n332), .S(n217), .Z(B[15]) );
  INV_X2 U307 ( .A(n340), .ZN(n332) );
  MUX2_X1 U308 ( .A(n341), .B(n317), .S(n210), .Z(n340) );
  MUX2_X1 U309 ( .A(n342), .B(n289), .S(n207), .Z(n317) );
  MUX2_X1 U310 ( .A(n343), .B(n330), .S(n212), .Z(n289) );
  MUX2_X1 U311 ( .A(n344), .B(n345), .S(n203), .Z(n330) );
  MUX2_X1 U312 ( .A(n346), .B(n339), .S(n217), .Z(B[14]) );
  INV_X2 U313 ( .A(n347), .ZN(n339) );
  MUX2_X1 U314 ( .A(n348), .B(n322), .S(n211), .Z(n347) );
  MUX2_X1 U315 ( .A(n349), .B(n294), .S(n207), .Z(n322) );
  MUX2_X1 U316 ( .A(n350), .B(n336), .S(n212), .Z(n294) );
  MUX2_X1 U317 ( .A(n351), .B(n352), .S(n203), .Z(n336) );
  MUX2_X1 U318 ( .A(n353), .B(n346), .S(n217), .Z(B[13]) );
  INV_X2 U319 ( .A(n354), .ZN(n346) );
  MUX2_X1 U320 ( .A(n355), .B(n328), .S(n211), .Z(n354) );
  MUX2_X1 U321 ( .A(n356), .B(n300), .S(n207), .Z(n328) );
  MUX2_X1 U322 ( .A(n357), .B(n343), .S(n212), .Z(n300) );
  MUX2_X1 U323 ( .A(n358), .B(n359), .S(n203), .Z(n343) );
  MUX2_X1 U324 ( .A(n360), .B(n353), .S(n217), .Z(B[12]) );
  INV_X2 U325 ( .A(n361), .ZN(n353) );
  MUX2_X1 U326 ( .A(n223), .B(n334), .S(n211), .Z(n361) );
  MUX2_X1 U327 ( .A(n240), .B(n305), .S(n207), .Z(n334) );
  MUX2_X1 U328 ( .A(n362), .B(n350), .S(n212), .Z(n305) );
  MUX2_X1 U329 ( .A(n363), .B(n364), .S(n203), .Z(n350) );
  MUX2_X1 U330 ( .A(n365), .B(n366), .S(n212), .Z(n240) );
  MUX2_X1 U331 ( .A(n367), .B(n335), .S(n207), .Z(n223) );
  MUX2_X1 U332 ( .A(n368), .B(n369), .S(n213), .Z(n335) );
  MUX2_X1 U333 ( .A(n370), .B(n360), .S(n217), .Z(B[11]) );
  INV_X2 U334 ( .A(n371), .ZN(n360) );
  MUX2_X1 U335 ( .A(n227), .B(n341), .S(n211), .Z(n371) );
  MUX2_X1 U336 ( .A(n245), .B(n318), .S(n207), .Z(n341) );
  MUX2_X1 U337 ( .A(n372), .B(n357), .S(n213), .Z(n318) );
  MUX2_X1 U338 ( .A(n373), .B(n374), .S(n203), .Z(n357) );
  MUX2_X1 U339 ( .A(n375), .B(n376), .S(n213), .Z(n245) );
  MUX2_X1 U340 ( .A(n377), .B(n342), .S(n207), .Z(n227) );
  MUX2_X1 U341 ( .A(n378), .B(n379), .S(n213), .Z(n342) );
  MUX2_X1 U342 ( .A(n219), .B(n370), .S(n217), .Z(B[10]) );
  INV_X2 U343 ( .A(n380), .ZN(n370) );
  MUX2_X1 U344 ( .A(n231), .B(n348), .S(n211), .Z(n380) );
  MUX2_X1 U345 ( .A(n255), .B(n323), .S(n208), .Z(n348) );
  MUX2_X1 U346 ( .A(n369), .B(n362), .S(n213), .Z(n323) );
  MUX2_X1 U347 ( .A(n381), .B(n382), .S(n203), .Z(n362) );
  MUX2_X1 U348 ( .A(n383), .B(n384), .S(n203), .Z(n369) );
  MUX2_X1 U349 ( .A(n385), .B(n365), .S(n213), .Z(n255) );
  MUX2_X1 U350 ( .A(n386), .B(n387), .S(n203), .Z(n365) );
  MUX2_X1 U351 ( .A(n257), .B(n349), .S(n208), .Z(n231) );
  MUX2_X1 U352 ( .A(n366), .B(n368), .S(n213), .Z(n349) );
  MUX2_X1 U353 ( .A(n388), .B(n389), .S(n203), .Z(n368) );
  MUX2_X1 U354 ( .A(n390), .B(n391), .S(n203), .Z(n366) );
  MUX2_X1 U355 ( .A(n392), .B(n393), .S(n213), .Z(n257) );
  INV_X2 U356 ( .A(n394), .ZN(n219) );
  MUX2_X1 U357 ( .A(n235), .B(n355), .S(n211), .Z(n394) );
  MUX2_X1 U358 ( .A(n309), .B(n329), .S(n208), .Z(n355) );
  MUX2_X1 U359 ( .A(n379), .B(n372), .S(n213), .Z(n329) );
  MUX2_X1 U360 ( .A(n395), .B(n396), .S(n203), .Z(n372) );
  MUX2_X1 U361 ( .A(n397), .B(n398), .S(n204), .Z(n379) );
  MUX2_X1 U362 ( .A(n399), .B(n375), .S(n213), .Z(n309) );
  MUX2_X1 U363 ( .A(n400), .B(n401), .S(n204), .Z(n375) );
  MUX2_X1 U364 ( .A(n312), .B(n356), .S(n208), .Z(n235) );
  MUX2_X1 U365 ( .A(n376), .B(n378), .S(n213), .Z(n356) );
  MUX2_X1 U366 ( .A(n402), .B(n403), .S(n204), .Z(n378) );
  MUX2_X1 U367 ( .A(n404), .B(n405), .S(n204), .Z(n376) );
  MUX2_X1 U368 ( .A(n406), .B(n407), .S(n213), .Z(n312) );
  MUX2_X1 U369 ( .A(n247), .B(n307), .S(n217), .Z(B[0]) );
  INV_X2 U370 ( .A(n408), .ZN(n307) );
  MUX2_X1 U371 ( .A(n265), .B(n238), .S(n211), .Z(n408) );
  MUX2_X1 U372 ( .A(n285), .B(n367), .S(n208), .Z(n238) );
  MUX2_X1 U373 ( .A(n393), .B(n385), .S(n214), .Z(n367) );
  MUX2_X1 U374 ( .A(n338), .B(n337), .S(n204), .Z(n385) );
  INV_X2 U375 ( .A(A[31]), .ZN(n337) );
  MUX2_X1 U376 ( .A(n352), .B(n351), .S(n204), .Z(n393) );
  MUX2_X1 U377 ( .A(n296), .B(n274), .S(n214), .Z(n285) );
  MUX2_X1 U378 ( .A(n384), .B(n383), .S(n204), .Z(n274) );
  MUX2_X1 U379 ( .A(n389), .B(n388), .S(n204), .Z(n296) );
  MUX2_X1 U380 ( .A(n306), .B(n239), .S(n208), .Z(n265) );
  MUX2_X1 U381 ( .A(n275), .B(n392), .S(n214), .Z(n239) );
  MUX2_X1 U382 ( .A(n364), .B(n363), .S(n204), .Z(n392) );
  MUX2_X1 U383 ( .A(n382), .B(n381), .S(n204), .Z(n275) );
  MUX2_X1 U384 ( .A(n325), .B(n295), .S(n214), .Z(n306) );
  MUX2_X1 U385 ( .A(n391), .B(n390), .S(n204), .Z(n295) );
  MUX2_X1 U386 ( .A(n387), .B(n386), .S(n204), .Z(n325) );
  INV_X2 U387 ( .A(n409), .ZN(n247) );
  MUX2_X1 U388 ( .A(n269), .B(n243), .S(n211), .Z(n409) );
  MUX2_X1 U389 ( .A(n290), .B(n377), .S(n208), .Z(n243) );
  MUX2_X1 U390 ( .A(n407), .B(n399), .S(n214), .Z(n377) );
  MUX2_X1 U391 ( .A(n345), .B(n344), .S(n205), .Z(n399) );
  MUX2_X1 U392 ( .A(n359), .B(n358), .S(n205), .Z(n407) );
  MUX2_X1 U393 ( .A(n314), .B(n310), .S(n214), .Z(n290) );
  MUX2_X1 U394 ( .A(n398), .B(n397), .S(n205), .Z(n310) );
  MUX2_X1 U395 ( .A(n403), .B(n402), .S(n205), .Z(n314) );
  MUX2_X1 U396 ( .A(n319), .B(n244), .S(n208), .Z(n269) );
  MUX2_X1 U397 ( .A(n311), .B(n406), .S(n214), .Z(n244) );
  MUX2_X1 U398 ( .A(n374), .B(n373), .S(n205), .Z(n406) );
  MUX2_X1 U399 ( .A(n396), .B(n395), .S(n205), .Z(n311) );
  MUX2_X1 U400 ( .A(n331), .B(n313), .S(n214), .Z(n319) );
  MUX2_X1 U401 ( .A(n405), .B(n404), .S(n205), .Z(n313) );
  MUX2_X1 U402 ( .A(n401), .B(n400), .S(n205), .Z(n331) );
endmodule


module up_island_DW_sra_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  INV_X1 U170 ( .A(A[18]), .ZN(n1580) );
  INV_X1 U171 ( .A(A[15]), .ZN(n1592) );
  INV_X1 U172 ( .A(A[19]), .ZN(n1556) );
  INV_X1 U173 ( .A(A[20]), .ZN(n1578) );
  INV_X1 U174 ( .A(A[21]), .ZN(n1554) );
  INV_X1 U175 ( .A(A[9]), .ZN(n1608) );
  INV_X1 U176 ( .A(A[10]), .ZN(n1640) );
  INV_X1 U177 ( .A(A[22]), .ZN(n1568) );
  INV_X1 U178 ( .A(A[23]), .ZN(n1544) );
  INV_X1 U179 ( .A(A[8]), .ZN(n1642) );
  INV_X1 U180 ( .A(A[16]), .ZN(n1572) );
  INV_X1 U181 ( .A(A[17]), .ZN(n1548) );
  INV_X1 U182 ( .A(A[28]), .ZN(n1488) );
  INV_X1 U183 ( .A(A[27]), .ZN(n1502) );
  INV_X1 U184 ( .A(A[25]), .ZN(n1542) );
  INV_X1 U185 ( .A(A[30]), .ZN(n1458) );
  INV_X1 U186 ( .A(A[7]), .ZN(n1598) );
  INV_X1 U187 ( .A(A[14]), .ZN(n1621) );
  INV_X1 U188 ( .A(A[13]), .ZN(n1594) );
  INV_X1 U189 ( .A(A[11]), .ZN(n1606) );
  INV_X1 U190 ( .A(A[12]), .ZN(n1623) );
  INV_X1 U191 ( .A(A[29]), .ZN(n1474) );
  INV_X1 U192 ( .A(A[5]), .ZN(n1600) );
  INV_X1 U193 ( .A(A[26]), .ZN(n1522) );
  INV_X1 U194 ( .A(A[24]), .ZN(n1566) );
  INV_X1 U195 ( .A(A[6]), .ZN(n1627) );
  INV_X1 U196 ( .A(A[4]), .ZN(n1629) );
  INV_X1 U197 ( .A(A[3]), .ZN(n1612) );
  INV_X1 U198 ( .A(A[2]), .ZN(n1635) );
  INV_X1 U199 ( .A(SH[1]), .ZN(n1150) );
  INV_X1 U200 ( .A(SH[1]), .ZN(n1152) );
  INV_X1 U201 ( .A(SH[1]), .ZN(n1151) );
  BUF_X1 U202 ( .A(SH[4]), .Z(n1106) );
  BUF_X1 U203 ( .A(SH[4]), .Z(n1107) );
  BUF_X1 U204 ( .A(SH[4]), .Z(n1108) );
  INV_X1 U205 ( .A(n1138), .ZN(n1109) );
  INV_X1 U206 ( .A(n1139), .ZN(n1110) );
  INV_X1 U207 ( .A(n1139), .ZN(n1111) );
  INV_X1 U208 ( .A(n1139), .ZN(n1112) );
  INV_X1 U209 ( .A(n1140), .ZN(n1113) );
  BUF_X1 U210 ( .A(SH[3]), .Z(n1114) );
  BUF_X1 U211 ( .A(SH[3]), .Z(n1115) );
  BUF_X1 U212 ( .A(SH[3]), .Z(n1116) );
  BUF_X1 U213 ( .A(SH[3]), .Z(n1117) );
  BUF_X1 U214 ( .A(SH[3]), .Z(n1118) );
  BUF_X1 U215 ( .A(SH[3]), .Z(n1119) );
  BUF_X1 U216 ( .A(SH[3]), .Z(n1120) );
  BUF_X1 U217 ( .A(SH[3]), .Z(n1121) );
  BUF_X1 U218 ( .A(SH[3]), .Z(n1122) );
  BUF_X1 U219 ( .A(SH[3]), .Z(n1123) );
  BUF_X1 U220 ( .A(SH[3]), .Z(n1124) );
  BUF_X1 U221 ( .A(SH[3]), .Z(n1125) );
  BUF_X1 U222 ( .A(SH[3]), .Z(n1126) );
  BUF_X1 U223 ( .A(SH[3]), .Z(n1127) );
  BUF_X1 U224 ( .A(SH[3]), .Z(n1128) );
  BUF_X1 U225 ( .A(SH[3]), .Z(n1129) );
  BUF_X1 U226 ( .A(SH[3]), .Z(n1130) );
  BUF_X1 U227 ( .A(SH[3]), .Z(n1131) );
  BUF_X1 U228 ( .A(SH[3]), .Z(n1132) );
  BUF_X1 U229 ( .A(SH[3]), .Z(n1133) );
  BUF_X1 U230 ( .A(SH[3]), .Z(n1134) );
  BUF_X1 U231 ( .A(SH[3]), .Z(n1135) );
  BUF_X1 U232 ( .A(SH[3]), .Z(n1136) );
  BUF_X1 U233 ( .A(SH[3]), .Z(n1137) );
  BUF_X1 U234 ( .A(SH[3]), .Z(n1138) );
  BUF_X1 U235 ( .A(SH[3]), .Z(n1139) );
  BUF_X1 U236 ( .A(SH[3]), .Z(n1140) );
  INV_X1 U237 ( .A(n1145), .ZN(n1141) );
  INV_X1 U238 ( .A(n1145), .ZN(n1142) );
  INV_X1 U239 ( .A(n1145), .ZN(n1143) );
  INV_X1 U240 ( .A(n1145), .ZN(n1144) );
  INV_X4 U241 ( .A(SH[2]), .ZN(n1145) );
  INV_X1 U242 ( .A(n1151), .ZN(n1146) );
  INV_X1 U243 ( .A(n1151), .ZN(n1147) );
  INV_X1 U244 ( .A(n1151), .ZN(n1148) );
  INV_X1 U245 ( .A(n1151), .ZN(n1149) );
  INV_X1 U246 ( .A(n1186), .ZN(n1153) );
  INV_X1 U247 ( .A(n1187), .ZN(n1154) );
  INV_X1 U248 ( .A(n1187), .ZN(n1155) );
  INV_X1 U249 ( .A(n1187), .ZN(n1156) );
  INV_X1 U250 ( .A(n1188), .ZN(n1157) );
  BUF_X1 U251 ( .A(SH[0]), .Z(n1158) );
  BUF_X1 U252 ( .A(SH[0]), .Z(n1159) );
  BUF_X1 U253 ( .A(SH[0]), .Z(n1160) );
  BUF_X1 U254 ( .A(SH[0]), .Z(n1161) );
  BUF_X1 U255 ( .A(SH[0]), .Z(n1162) );
  BUF_X1 U256 ( .A(SH[0]), .Z(n1163) );
  BUF_X1 U257 ( .A(SH[0]), .Z(n1164) );
  BUF_X1 U258 ( .A(SH[0]), .Z(n1165) );
  BUF_X1 U259 ( .A(SH[0]), .Z(n1166) );
  BUF_X1 U260 ( .A(SH[0]), .Z(n1167) );
  BUF_X1 U261 ( .A(SH[0]), .Z(n1168) );
  BUF_X1 U262 ( .A(SH[0]), .Z(n1169) );
  BUF_X1 U263 ( .A(SH[0]), .Z(n1170) );
  BUF_X1 U264 ( .A(SH[0]), .Z(n1171) );
  BUF_X1 U265 ( .A(SH[0]), .Z(n1172) );
  BUF_X1 U266 ( .A(SH[0]), .Z(n1173) );
  BUF_X1 U267 ( .A(SH[0]), .Z(n1174) );
  BUF_X1 U268 ( .A(SH[0]), .Z(n1175) );
  BUF_X1 U269 ( .A(SH[0]), .Z(n1176) );
  BUF_X1 U270 ( .A(SH[0]), .Z(n1177) );
  BUF_X1 U271 ( .A(SH[0]), .Z(n1178) );
  BUF_X1 U272 ( .A(SH[0]), .Z(n1179) );
  BUF_X1 U273 ( .A(SH[0]), .Z(n1180) );
  BUF_X1 U274 ( .A(SH[0]), .Z(n1181) );
  BUF_X1 U275 ( .A(SH[0]), .Z(n1182) );
  BUF_X1 U276 ( .A(SH[0]), .Z(n1183) );
  BUF_X1 U277 ( .A(SH[0]), .Z(n1184) );
  BUF_X1 U278 ( .A(SH[0]), .Z(n1185) );
  BUF_X1 U279 ( .A(SH[0]), .Z(n1186) );
  BUF_X1 U280 ( .A(SH[0]), .Z(n1187) );
  BUF_X1 U281 ( .A(SH[0]), .Z(n1188) );
  NAND2_X2 U282 ( .A1(n1189), .A2(n1190), .ZN(B[9]) );
  MUX2_X1 U283 ( .A(n1191), .B(n1192), .S(n1141), .Z(n1190) );
  NAND2_X2 U284 ( .A1(n1186), .A2(n1193), .ZN(n1192) );
  NAND2_X2 U285 ( .A1(n1185), .A2(n1194), .ZN(n1191) );
  MUX2_X1 U286 ( .A(n1195), .B(n1196), .S(n1144), .Z(n1189) );
  NAND2_X2 U287 ( .A1(n1197), .A2(n1155), .ZN(n1196) );
  NAND2_X2 U288 ( .A1(n1198), .A2(n1153), .ZN(n1195) );
  NAND2_X2 U289 ( .A1(n1199), .A2(n1200), .ZN(B[8]) );
  MUX2_X1 U290 ( .A(n1201), .B(n1202), .S(n1144), .Z(n1200) );
  NAND2_X2 U291 ( .A1(n1185), .A2(n1197), .ZN(n1202) );
  NAND2_X2 U292 ( .A1(n1184), .A2(n1198), .ZN(n1201) );
  MUX2_X1 U293 ( .A(n1203), .B(n1204), .S(n1144), .Z(n1199) );
  NAND2_X2 U294 ( .A1(n1205), .A2(n1153), .ZN(n1204) );
  NAND2_X2 U295 ( .A1(n1206), .A2(n1153), .ZN(n1203) );
  NAND2_X2 U296 ( .A1(n1207), .A2(n1208), .ZN(B[7]) );
  MUX2_X1 U297 ( .A(n1209), .B(n1210), .S(n1144), .Z(n1208) );
  NAND2_X2 U298 ( .A1(n1184), .A2(n1205), .ZN(n1210) );
  NAND2_X2 U299 ( .A1(n1183), .A2(n1206), .ZN(n1209) );
  MUX2_X1 U300 ( .A(n1211), .B(n1212), .S(n1144), .Z(n1207) );
  NAND2_X2 U301 ( .A1(n1213), .A2(n1153), .ZN(n1212) );
  NAND2_X2 U302 ( .A1(n1214), .A2(n1153), .ZN(n1211) );
  NAND2_X2 U303 ( .A1(n1215), .A2(n1216), .ZN(B[6]) );
  MUX2_X1 U304 ( .A(n1217), .B(n1218), .S(n1144), .Z(n1216) );
  NAND2_X2 U305 ( .A1(n1183), .A2(n1213), .ZN(n1218) );
  NAND2_X2 U306 ( .A1(n1182), .A2(n1214), .ZN(n1217) );
  MUX2_X1 U307 ( .A(n1219), .B(n1220), .S(n1144), .Z(n1215) );
  NAND2_X2 U308 ( .A1(n1194), .A2(n1153), .ZN(n1220) );
  NAND2_X2 U309 ( .A1(n1221), .A2(n1153), .ZN(n1219) );
  NAND2_X2 U310 ( .A1(n1222), .A2(n1223), .ZN(B[5]) );
  MUX2_X1 U311 ( .A(n1224), .B(n1225), .S(n1144), .Z(n1223) );
  NAND2_X2 U312 ( .A1(n1182), .A2(n1194), .ZN(n1225) );
  NAND2_X2 U313 ( .A1(n1181), .A2(n1221), .ZN(n1224) );
  MUX2_X1 U314 ( .A(n1226), .B(n1227), .S(n1143), .Z(n1222) );
  NAND2_X2 U315 ( .A1(n1198), .A2(n1153), .ZN(n1227) );
  NAND2_X2 U316 ( .A1(n1228), .A2(n1153), .ZN(n1226) );
  NAND2_X2 U317 ( .A1(n1229), .A2(n1230), .ZN(B[4]) );
  MUX2_X1 U318 ( .A(n1231), .B(n1232), .S(n1143), .Z(n1230) );
  NAND2_X2 U319 ( .A1(n1181), .A2(n1198), .ZN(n1232) );
  NAND2_X2 U320 ( .A1(n1233), .A2(n1234), .ZN(n1198) );
  MUX2_X1 U321 ( .A(n1235), .B(n1236), .S(n1146), .Z(n1234) );
  NAND2_X2 U322 ( .A1(n1133), .A2(n1237), .ZN(n1236) );
  NAND2_X2 U323 ( .A1(n1135), .A2(n1238), .ZN(n1235) );
  MUX2_X1 U324 ( .A(n1239), .B(n1240), .S(n1149), .Z(n1233) );
  NAND2_X2 U325 ( .A1(n1241), .A2(n1110), .ZN(n1240) );
  NAND2_X2 U326 ( .A1(n1242), .A2(n1109), .ZN(n1239) );
  NAND2_X2 U327 ( .A1(n1180), .A2(n1228), .ZN(n1231) );
  MUX2_X1 U328 ( .A(n1243), .B(n1244), .S(n1143), .Z(n1229) );
  NAND2_X2 U329 ( .A1(n1206), .A2(n1153), .ZN(n1244) );
  NAND2_X2 U330 ( .A1(n1245), .A2(n1153), .ZN(n1243) );
  NAND2_X2 U331 ( .A1(n1246), .A2(n1247), .ZN(B[3]) );
  MUX2_X1 U332 ( .A(n1248), .B(n1249), .S(n1143), .Z(n1247) );
  NAND2_X2 U333 ( .A1(n1180), .A2(n1206), .ZN(n1249) );
  NAND2_X2 U334 ( .A1(n1250), .A2(n1251), .ZN(n1206) );
  MUX2_X1 U335 ( .A(n1252), .B(n1253), .S(n1149), .Z(n1251) );
  NAND2_X2 U336 ( .A1(n1133), .A2(n1254), .ZN(n1253) );
  NAND2_X2 U337 ( .A1(n1135), .A2(n1255), .ZN(n1252) );
  MUX2_X1 U338 ( .A(n1256), .B(n1257), .S(n1149), .Z(n1250) );
  NAND2_X2 U339 ( .A1(n1258), .A2(n1109), .ZN(n1257) );
  NAND2_X2 U340 ( .A1(n1259), .A2(n1109), .ZN(n1256) );
  NAND2_X2 U341 ( .A1(n1179), .A2(n1245), .ZN(n1248) );
  MUX2_X1 U342 ( .A(n1260), .B(n1261), .S(n1143), .Z(n1246) );
  NAND2_X2 U343 ( .A1(n1214), .A2(n1153), .ZN(n1261) );
  NAND2_X2 U344 ( .A1(n1262), .A2(n1154), .ZN(n1260) );
  NAND2_X2 U345 ( .A1(n1263), .A2(n1264), .ZN(B[30]) );
  NAND2_X2 U346 ( .A1(n1141), .A2(\A[31] ), .ZN(n1264) );
  MUX2_X1 U347 ( .A(n1265), .B(n1266), .S(n1186), .Z(n1263) );
  NAND2_X2 U348 ( .A1(n1267), .A2(n1145), .ZN(n1265) );
  NAND2_X2 U349 ( .A1(n1268), .A2(n1269), .ZN(B[2]) );
  MUX2_X1 U350 ( .A(n1270), .B(n1271), .S(n1143), .Z(n1269) );
  NAND2_X2 U351 ( .A1(n1179), .A2(n1214), .ZN(n1271) );
  NAND2_X2 U352 ( .A1(n1272), .A2(n1273), .ZN(n1214) );
  MUX2_X1 U353 ( .A(n1274), .B(n1275), .S(n1149), .Z(n1273) );
  NAND2_X2 U354 ( .A1(n1131), .A2(n1238), .ZN(n1275) );
  NAND2_X2 U355 ( .A1(n1134), .A2(n1276), .ZN(n1274) );
  MUX2_X1 U356 ( .A(n1277), .B(n1278), .S(n1148), .Z(n1272) );
  NAND2_X2 U357 ( .A1(n1242), .A2(n1109), .ZN(n1278) );
  NAND2_X2 U358 ( .A1(n1279), .A2(n1109), .ZN(n1277) );
  NAND2_X2 U359 ( .A1(n1178), .A2(n1262), .ZN(n1270) );
  NAND2_X2 U360 ( .A1(n1280), .A2(n1281), .ZN(n1262) );
  MUX2_X1 U361 ( .A(n1282), .B(n1283), .S(n1148), .Z(n1281) );
  NAND2_X2 U362 ( .A1(n1132), .A2(n1284), .ZN(n1283) );
  NAND2_X2 U363 ( .A1(n1134), .A2(n1241), .ZN(n1282) );
  MUX2_X1 U364 ( .A(n1285), .B(n1286), .S(n1148), .Z(n1280) );
  NAND2_X2 U365 ( .A1(n1287), .A2(n1109), .ZN(n1286) );
  NAND2_X2 U366 ( .A1(n1288), .A2(n1109), .ZN(n1285) );
  MUX2_X1 U367 ( .A(n1289), .B(n1290), .S(n1143), .Z(n1268) );
  NAND2_X2 U368 ( .A1(n1221), .A2(n1154), .ZN(n1290) );
  NAND2_X2 U369 ( .A1(n1291), .A2(n1154), .ZN(n1289) );
  NAND2_X2 U370 ( .A1(n1292), .A2(n1293), .ZN(B[29]) );
  NAND3_X1 U371 ( .A1(n1157), .A2(n1145), .A3(n1294), .ZN(n1293) );
  MUX2_X1 U372 ( .A(n1295), .B(n1266), .S(n1143), .Z(n1292) );
  NAND2_X2 U373 ( .A1(n1178), .A2(n1267), .ZN(n1295) );
  NAND2_X2 U374 ( .A1(n1296), .A2(n1297), .ZN(B[28]) );
  NAND3_X1 U375 ( .A1(n1157), .A2(n1145), .A3(n1298), .ZN(n1297) );
  MUX2_X1 U376 ( .A(n1299), .B(n1266), .S(n1143), .Z(n1296) );
  NAND2_X2 U377 ( .A1(n1177), .A2(n1294), .ZN(n1299) );
  NAND2_X2 U378 ( .A1(n1300), .A2(n1301), .ZN(B[27]) );
  NAND3_X1 U379 ( .A1(n1157), .A2(n1145), .A3(n1302), .ZN(n1301) );
  MUX2_X1 U380 ( .A(n1303), .B(n1266), .S(n1143), .Z(n1300) );
  NAND2_X2 U381 ( .A1(n1177), .A2(n1298), .ZN(n1303) );
  NAND2_X2 U382 ( .A1(n1304), .A2(n1305), .ZN(B[26]) );
  MUX2_X1 U383 ( .A(n1306), .B(n1307), .S(n1143), .Z(n1305) );
  NAND2_X2 U384 ( .A1(n1176), .A2(\A[31] ), .ZN(n1307) );
  NAND2_X2 U385 ( .A1(n1176), .A2(n1302), .ZN(n1306) );
  MUX2_X1 U386 ( .A(n1308), .B(n1309), .S(n1143), .Z(n1304) );
  NAND2_X2 U387 ( .A1(n1267), .A2(n1154), .ZN(n1309) );
  NAND2_X2 U388 ( .A1(n1310), .A2(n1154), .ZN(n1308) );
  NAND2_X2 U389 ( .A1(n1311), .A2(n1312), .ZN(B[25]) );
  MUX2_X1 U390 ( .A(n1313), .B(n1314), .S(n1143), .Z(n1312) );
  NAND2_X2 U391 ( .A1(n1175), .A2(n1267), .ZN(n1314) );
  OAI21_X2 U392 ( .B1(n1266), .B2(n1150), .A(n1315), .ZN(n1267) );
  MUX2_X1 U393 ( .A(n1316), .B(n1266), .S(n1138), .Z(n1315) );
  NAND2_X2 U394 ( .A1(n1317), .A2(n1150), .ZN(n1316) );
  NAND2_X2 U395 ( .A1(n1175), .A2(n1310), .ZN(n1313) );
  MUX2_X1 U396 ( .A(n1318), .B(n1319), .S(n1143), .Z(n1311) );
  NAND2_X2 U397 ( .A1(n1294), .A2(n1154), .ZN(n1319) );
  NAND2_X2 U398 ( .A1(n1320), .A2(n1154), .ZN(n1318) );
  NAND2_X2 U399 ( .A1(n1321), .A2(n1322), .ZN(B[24]) );
  MUX2_X1 U400 ( .A(n1323), .B(n1324), .S(n1143), .Z(n1322) );
  NAND2_X2 U401 ( .A1(n1174), .A2(n1294), .ZN(n1324) );
  OAI21_X2 U402 ( .B1(n1266), .B2(n1151), .A(n1325), .ZN(n1294) );
  MUX2_X1 U403 ( .A(n1326), .B(n1266), .S(n1138), .Z(n1325) );
  NAND2_X2 U404 ( .A1(n1327), .A2(n1150), .ZN(n1326) );
  NAND2_X2 U405 ( .A1(n1174), .A2(n1320), .ZN(n1323) );
  MUX2_X1 U406 ( .A(n1328), .B(n1329), .S(n1143), .Z(n1321) );
  NAND2_X2 U407 ( .A1(n1298), .A2(n1154), .ZN(n1329) );
  NAND2_X2 U408 ( .A1(n1330), .A2(n1154), .ZN(n1328) );
  NAND2_X2 U409 ( .A1(n1331), .A2(n1332), .ZN(B[23]) );
  MUX2_X1 U410 ( .A(n1333), .B(n1334), .S(n1143), .Z(n1332) );
  NAND2_X2 U411 ( .A1(n1173), .A2(n1298), .ZN(n1334) );
  NAND2_X2 U412 ( .A1(n1335), .A2(n1336), .ZN(n1298) );
  NAND3_X1 U413 ( .A1(n1152), .A2(n1113), .A3(n1337), .ZN(n1336) );
  MUX2_X1 U414 ( .A(n1338), .B(n1266), .S(n1137), .Z(n1335) );
  NAND2_X2 U415 ( .A1(n1146), .A2(n1317), .ZN(n1338) );
  NAND2_X2 U416 ( .A1(n1172), .A2(n1330), .ZN(n1333) );
  MUX2_X1 U417 ( .A(n1339), .B(n1340), .S(n1142), .Z(n1331) );
  NAND2_X2 U418 ( .A1(n1302), .A2(n1154), .ZN(n1340) );
  NAND2_X2 U419 ( .A1(n1341), .A2(n1154), .ZN(n1339) );
  NAND2_X2 U420 ( .A1(n1342), .A2(n1343), .ZN(B[22]) );
  MUX2_X1 U421 ( .A(n1344), .B(n1345), .S(n1142), .Z(n1343) );
  NAND2_X2 U422 ( .A1(n1172), .A2(n1302), .ZN(n1345) );
  NAND2_X2 U423 ( .A1(n1346), .A2(n1347), .ZN(n1302) );
  NAND3_X1 U424 ( .A1(n1152), .A2(n1112), .A3(n1348), .ZN(n1347) );
  MUX2_X1 U425 ( .A(n1349), .B(n1266), .S(n1136), .Z(n1346) );
  NAND2_X2 U426 ( .A1(n1146), .A2(n1327), .ZN(n1349) );
  NAND2_X2 U427 ( .A1(n1171), .A2(n1341), .ZN(n1344) );
  MUX2_X1 U428 ( .A(n1350), .B(n1351), .S(n1142), .Z(n1342) );
  NAND2_X2 U429 ( .A1(n1310), .A2(n1154), .ZN(n1351) );
  NAND2_X2 U430 ( .A1(n1352), .A2(n1155), .ZN(n1350) );
  NAND2_X2 U431 ( .A1(n1353), .A2(n1354), .ZN(B[21]) );
  MUX2_X1 U432 ( .A(n1355), .B(n1356), .S(n1142), .Z(n1354) );
  NAND2_X2 U433 ( .A1(n1171), .A2(n1310), .ZN(n1356) );
  NAND2_X2 U434 ( .A1(n1357), .A2(n1358), .ZN(n1310) );
  NAND3_X1 U435 ( .A1(n1152), .A2(n1113), .A3(n1359), .ZN(n1358) );
  MUX2_X1 U436 ( .A(n1360), .B(n1266), .S(n1137), .Z(n1357) );
  NAND2_X2 U437 ( .A1(n1146), .A2(n1337), .ZN(n1360) );
  NAND2_X2 U438 ( .A1(n1170), .A2(n1352), .ZN(n1355) );
  MUX2_X1 U439 ( .A(n1361), .B(n1362), .S(n1142), .Z(n1353) );
  NAND2_X2 U440 ( .A1(n1320), .A2(n1155), .ZN(n1362) );
  NAND2_X2 U441 ( .A1(n1363), .A2(n1155), .ZN(n1361) );
  NAND2_X2 U442 ( .A1(n1364), .A2(n1365), .ZN(B[20]) );
  MUX2_X1 U443 ( .A(n1366), .B(n1367), .S(n1142), .Z(n1365) );
  NAND2_X2 U444 ( .A1(n1170), .A2(n1320), .ZN(n1367) );
  NAND2_X2 U445 ( .A1(n1368), .A2(n1369), .ZN(n1320) );
  NAND3_X1 U446 ( .A1(n1152), .A2(n1112), .A3(n1370), .ZN(n1369) );
  MUX2_X1 U447 ( .A(n1371), .B(n1266), .S(n1136), .Z(n1368) );
  NAND2_X2 U448 ( .A1(n1146), .A2(n1348), .ZN(n1371) );
  NAND2_X2 U449 ( .A1(n1169), .A2(n1363), .ZN(n1366) );
  MUX2_X1 U450 ( .A(n1372), .B(n1373), .S(n1142), .Z(n1364) );
  NAND2_X2 U451 ( .A1(n1330), .A2(n1155), .ZN(n1373) );
  NAND2_X2 U452 ( .A1(n1374), .A2(n1155), .ZN(n1372) );
  NAND2_X2 U453 ( .A1(n1375), .A2(n1376), .ZN(B[1]) );
  MUX2_X1 U454 ( .A(n1377), .B(n1378), .S(n1142), .Z(n1376) );
  NAND2_X2 U455 ( .A1(n1169), .A2(n1221), .ZN(n1378) );
  NAND2_X2 U456 ( .A1(n1379), .A2(n1380), .ZN(n1221) );
  MUX2_X1 U457 ( .A(n1381), .B(n1382), .S(n1148), .Z(n1380) );
  NAND2_X2 U458 ( .A1(n1130), .A2(n1255), .ZN(n1382) );
  NAND2_X2 U459 ( .A1(n1132), .A2(n1383), .ZN(n1381) );
  MUX2_X1 U460 ( .A(n1384), .B(n1385), .S(n1148), .Z(n1379) );
  NAND2_X2 U461 ( .A1(n1259), .A2(n1109), .ZN(n1385) );
  NAND2_X2 U462 ( .A1(n1386), .A2(n1109), .ZN(n1384) );
  NAND2_X2 U463 ( .A1(n1168), .A2(n1291), .ZN(n1377) );
  NAND2_X2 U464 ( .A1(n1387), .A2(n1388), .ZN(n1291) );
  MUX2_X1 U465 ( .A(n1389), .B(n1390), .S(n1148), .Z(n1388) );
  NAND2_X2 U466 ( .A1(n1130), .A2(n1391), .ZN(n1390) );
  NAND2_X2 U467 ( .A1(n1131), .A2(n1258), .ZN(n1389) );
  MUX2_X1 U468 ( .A(n1392), .B(n1393), .S(n1148), .Z(n1387) );
  NAND2_X2 U469 ( .A1(n1394), .A2(n1109), .ZN(n1393) );
  NAND2_X2 U470 ( .A1(n1395), .A2(n1109), .ZN(n1392) );
  MUX2_X1 U471 ( .A(n1396), .B(n1397), .S(n1142), .Z(n1375) );
  NAND2_X2 U472 ( .A1(n1228), .A2(n1155), .ZN(n1397) );
  NAND2_X2 U473 ( .A1(n1398), .A2(n1155), .ZN(n1396) );
  NAND2_X2 U474 ( .A1(n1399), .A2(n1400), .ZN(B[19]) );
  MUX2_X1 U475 ( .A(n1401), .B(n1402), .S(n1142), .Z(n1400) );
  NAND2_X2 U476 ( .A1(n1168), .A2(n1330), .ZN(n1402) );
  NAND2_X2 U477 ( .A1(n1403), .A2(n1404), .ZN(n1330) );
  NAND3_X1 U478 ( .A1(n1152), .A2(n1112), .A3(n1405), .ZN(n1404) );
  MUX2_X1 U479 ( .A(n1406), .B(n1266), .S(n1137), .Z(n1403) );
  NAND2_X2 U480 ( .A1(n1146), .A2(n1359), .ZN(n1406) );
  NAND2_X2 U481 ( .A1(n1167), .A2(n1374), .ZN(n1401) );
  MUX2_X1 U482 ( .A(n1407), .B(n1408), .S(n1142), .Z(n1399) );
  NAND2_X2 U483 ( .A1(n1341), .A2(n1155), .ZN(n1408) );
  NAND2_X2 U484 ( .A1(n1409), .A2(n1155), .ZN(n1407) );
  NAND2_X2 U485 ( .A1(n1410), .A2(n1411), .ZN(B[18]) );
  MUX2_X1 U486 ( .A(n1412), .B(n1413), .S(n1142), .Z(n1411) );
  NAND2_X2 U487 ( .A1(n1167), .A2(n1341), .ZN(n1413) );
  NAND2_X2 U488 ( .A1(n1414), .A2(n1415), .ZN(n1341) );
  NAND3_X1 U489 ( .A1(n1152), .A2(n1112), .A3(n1416), .ZN(n1415) );
  MUX2_X1 U490 ( .A(n1417), .B(n1266), .S(n1136), .Z(n1414) );
  NAND2_X2 U491 ( .A1(n1146), .A2(n1370), .ZN(n1417) );
  NAND2_X2 U492 ( .A1(n1166), .A2(n1409), .ZN(n1412) );
  MUX2_X1 U493 ( .A(n1418), .B(n1419), .S(n1142), .Z(n1410) );
  NAND2_X2 U494 ( .A1(n1352), .A2(n1155), .ZN(n1419) );
  NAND2_X2 U495 ( .A1(n1420), .A2(n1155), .ZN(n1418) );
  NAND2_X2 U496 ( .A1(n1421), .A2(n1422), .ZN(B[17]) );
  MUX2_X1 U497 ( .A(n1423), .B(n1424), .S(n1142), .Z(n1422) );
  NAND2_X2 U498 ( .A1(n1166), .A2(n1352), .ZN(n1424) );
  NAND2_X2 U499 ( .A1(n1425), .A2(n1426), .ZN(n1352) );
  MUX2_X1 U500 ( .A(n1427), .B(n1428), .S(n1148), .Z(n1426) );
  NAND2_X2 U501 ( .A1(n1129), .A2(\A[31] ), .ZN(n1428) );
  NAND2_X2 U502 ( .A1(n1129), .A2(n1317), .ZN(n1427) );
  MUX2_X1 U503 ( .A(n1429), .B(n1430), .S(n1148), .Z(n1425) );
  NAND2_X2 U504 ( .A1(n1405), .A2(n1109), .ZN(n1430) );
  NAND2_X2 U505 ( .A1(n1431), .A2(n1110), .ZN(n1429) );
  NAND2_X2 U506 ( .A1(n1165), .A2(n1420), .ZN(n1423) );
  MUX2_X1 U507 ( .A(n1432), .B(n1433), .S(n1142), .Z(n1421) );
  NAND2_X2 U508 ( .A1(n1363), .A2(n1156), .ZN(n1433) );
  NAND2_X2 U509 ( .A1(n1434), .A2(n1156), .ZN(n1432) );
  NAND2_X2 U510 ( .A1(n1435), .A2(n1436), .ZN(B[16]) );
  MUX2_X1 U511 ( .A(n1437), .B(n1438), .S(n1142), .Z(n1436) );
  NAND2_X2 U512 ( .A1(n1165), .A2(n1363), .ZN(n1438) );
  NAND2_X2 U513 ( .A1(n1439), .A2(n1440), .ZN(n1363) );
  MUX2_X1 U514 ( .A(n1441), .B(n1442), .S(n1148), .Z(n1440) );
  NAND2_X2 U515 ( .A1(n1128), .A2(\A[31] ), .ZN(n1442) );
  NAND2_X2 U516 ( .A1(n1127), .A2(n1327), .ZN(n1441) );
  MUX2_X1 U517 ( .A(n1443), .B(n1444), .S(n1148), .Z(n1439) );
  NAND2_X2 U518 ( .A1(n1416), .A2(n1110), .ZN(n1444) );
  NAND2_X2 U519 ( .A1(n1445), .A2(n1110), .ZN(n1443) );
  NAND2_X2 U520 ( .A1(n1164), .A2(n1434), .ZN(n1437) );
  MUX2_X1 U521 ( .A(n1446), .B(n1447), .S(n1141), .Z(n1435) );
  NAND2_X2 U522 ( .A1(n1374), .A2(n1156), .ZN(n1447) );
  NAND2_X2 U523 ( .A1(n1448), .A2(n1156), .ZN(n1446) );
  NAND2_X2 U524 ( .A1(n1449), .A2(n1450), .ZN(B[15]) );
  MUX2_X1 U525 ( .A(n1451), .B(n1452), .S(n1141), .Z(n1450) );
  NAND2_X2 U526 ( .A1(n1164), .A2(n1374), .ZN(n1452) );
  NAND2_X2 U527 ( .A1(n1453), .A2(n1454), .ZN(n1374) );
  MUX2_X1 U528 ( .A(n1455), .B(n1456), .S(n1148), .Z(n1454) );
  NAND2_X2 U529 ( .A1(n1128), .A2(n1317), .ZN(n1456) );
  INV_X2 U530 ( .A(n1457), .ZN(n1317) );
  MUX2_X1 U531 ( .A(n1458), .B(n1266), .S(n1106), .Z(n1457) );
  NAND2_X2 U532 ( .A1(n1127), .A2(n1337), .ZN(n1455) );
  MUX2_X1 U533 ( .A(n1459), .B(n1460), .S(n1148), .Z(n1453) );
  NAND2_X2 U534 ( .A1(n1431), .A2(n1110), .ZN(n1460) );
  NAND2_X2 U535 ( .A1(n1461), .A2(n1110), .ZN(n1459) );
  NAND2_X2 U536 ( .A1(n1163), .A2(n1448), .ZN(n1451) );
  MUX2_X1 U537 ( .A(n1462), .B(n1463), .S(n1141), .Z(n1449) );
  NAND2_X2 U538 ( .A1(n1409), .A2(n1156), .ZN(n1463) );
  NAND2_X2 U539 ( .A1(n1464), .A2(n1156), .ZN(n1462) );
  NAND2_X2 U540 ( .A1(n1465), .A2(n1466), .ZN(B[14]) );
  MUX2_X1 U541 ( .A(n1467), .B(n1468), .S(n1141), .Z(n1466) );
  NAND2_X2 U542 ( .A1(n1163), .A2(n1409), .ZN(n1468) );
  NAND2_X2 U543 ( .A1(n1469), .A2(n1470), .ZN(n1409) );
  MUX2_X1 U544 ( .A(n1471), .B(n1472), .S(n1148), .Z(n1470) );
  NAND2_X2 U545 ( .A1(n1126), .A2(n1327), .ZN(n1472) );
  INV_X2 U546 ( .A(n1473), .ZN(n1327) );
  MUX2_X1 U547 ( .A(n1474), .B(n1266), .S(n1106), .Z(n1473) );
  NAND2_X2 U548 ( .A1(n1126), .A2(n1348), .ZN(n1471) );
  MUX2_X1 U549 ( .A(n1475), .B(n1476), .S(n1148), .Z(n1469) );
  NAND2_X2 U550 ( .A1(n1445), .A2(n1110), .ZN(n1476) );
  NAND2_X2 U551 ( .A1(n1237), .A2(n1110), .ZN(n1475) );
  NAND2_X2 U552 ( .A1(n1162), .A2(n1464), .ZN(n1467) );
  MUX2_X1 U553 ( .A(n1477), .B(n1478), .S(n1141), .Z(n1465) );
  NAND2_X2 U554 ( .A1(n1420), .A2(n1156), .ZN(n1478) );
  NAND2_X2 U555 ( .A1(n1193), .A2(n1156), .ZN(n1477) );
  NAND2_X2 U556 ( .A1(n1479), .A2(n1480), .ZN(B[13]) );
  MUX2_X1 U557 ( .A(n1481), .B(n1482), .S(n1141), .Z(n1480) );
  NAND2_X2 U558 ( .A1(n1162), .A2(n1420), .ZN(n1482) );
  NAND2_X2 U559 ( .A1(n1483), .A2(n1484), .ZN(n1420) );
  MUX2_X1 U560 ( .A(n1485), .B(n1486), .S(n1148), .Z(n1484) );
  NAND2_X2 U561 ( .A1(n1125), .A2(n1337), .ZN(n1486) );
  INV_X2 U562 ( .A(n1487), .ZN(n1337) );
  MUX2_X1 U563 ( .A(n1488), .B(n1266), .S(n1106), .Z(n1487) );
  NAND2_X2 U564 ( .A1(n1125), .A2(n1359), .ZN(n1485) );
  MUX2_X1 U565 ( .A(n1489), .B(n1490), .S(n1148), .Z(n1483) );
  NAND2_X2 U566 ( .A1(n1461), .A2(n1110), .ZN(n1490) );
  NAND2_X2 U567 ( .A1(n1254), .A2(n1110), .ZN(n1489) );
  NAND2_X2 U568 ( .A1(n1161), .A2(n1193), .ZN(n1481) );
  MUX2_X1 U569 ( .A(n1491), .B(n1492), .S(n1141), .Z(n1479) );
  NAND2_X2 U570 ( .A1(n1434), .A2(n1156), .ZN(n1492) );
  NAND2_X2 U571 ( .A1(n1197), .A2(n1156), .ZN(n1491) );
  NAND2_X2 U572 ( .A1(n1493), .A2(n1494), .ZN(B[12]) );
  MUX2_X1 U573 ( .A(n1495), .B(n1496), .S(n1141), .Z(n1494) );
  NAND2_X2 U574 ( .A1(n1161), .A2(n1434), .ZN(n1496) );
  NAND2_X2 U575 ( .A1(n1497), .A2(n1498), .ZN(n1434) );
  MUX2_X1 U576 ( .A(n1499), .B(n1500), .S(n1147), .Z(n1498) );
  NAND2_X2 U577 ( .A1(n1124), .A2(n1348), .ZN(n1500) );
  INV_X2 U578 ( .A(n1501), .ZN(n1348) );
  MUX2_X1 U579 ( .A(n1502), .B(n1266), .S(n1106), .Z(n1501) );
  NAND2_X2 U580 ( .A1(n1124), .A2(n1370), .ZN(n1499) );
  MUX2_X1 U581 ( .A(n1503), .B(n1504), .S(n1147), .Z(n1497) );
  NAND2_X2 U582 ( .A1(n1237), .A2(n1110), .ZN(n1504) );
  NAND2_X2 U583 ( .A1(n1238), .A2(n1110), .ZN(n1503) );
  NAND2_X2 U584 ( .A1(n1160), .A2(n1197), .ZN(n1495) );
  NAND2_X2 U585 ( .A1(n1505), .A2(n1506), .ZN(n1197) );
  MUX2_X1 U586 ( .A(n1507), .B(n1508), .S(n1147), .Z(n1506) );
  NAND2_X2 U587 ( .A1(n1123), .A2(n1416), .ZN(n1508) );
  NAND2_X2 U588 ( .A1(n1123), .A2(n1445), .ZN(n1507) );
  MUX2_X1 U589 ( .A(n1509), .B(n1510), .S(n1147), .Z(n1505) );
  NAND2_X2 U590 ( .A1(n1276), .A2(n1111), .ZN(n1510) );
  NAND2_X2 U591 ( .A1(n1284), .A2(n1111), .ZN(n1509) );
  MUX2_X1 U592 ( .A(n1511), .B(n1512), .S(n1141), .Z(n1493) );
  NAND2_X2 U593 ( .A1(n1448), .A2(n1157), .ZN(n1512) );
  NAND2_X2 U594 ( .A1(n1205), .A2(n1156), .ZN(n1511) );
  NAND2_X2 U595 ( .A1(n1513), .A2(n1514), .ZN(B[11]) );
  MUX2_X1 U596 ( .A(n1515), .B(n1516), .S(n1141), .Z(n1514) );
  NAND2_X2 U597 ( .A1(n1160), .A2(n1448), .ZN(n1516) );
  NAND2_X2 U598 ( .A1(n1517), .A2(n1518), .ZN(n1448) );
  MUX2_X1 U599 ( .A(n1519), .B(n1520), .S(n1147), .Z(n1518) );
  NAND2_X2 U600 ( .A1(n1122), .A2(n1359), .ZN(n1520) );
  INV_X2 U601 ( .A(n1521), .ZN(n1359) );
  MUX2_X1 U602 ( .A(n1522), .B(n1266), .S(n1106), .Z(n1521) );
  NAND2_X2 U603 ( .A1(n1122), .A2(n1405), .ZN(n1519) );
  MUX2_X1 U604 ( .A(n1523), .B(n1524), .S(n1147), .Z(n1517) );
  NAND2_X2 U605 ( .A1(n1254), .A2(n1111), .ZN(n1524) );
  NAND2_X2 U606 ( .A1(n1255), .A2(n1111), .ZN(n1523) );
  NAND2_X2 U607 ( .A1(n1159), .A2(n1205), .ZN(n1515) );
  NAND2_X2 U608 ( .A1(n1525), .A2(n1526), .ZN(n1205) );
  MUX2_X1 U609 ( .A(n1527), .B(n1528), .S(n1147), .Z(n1526) );
  NAND2_X2 U610 ( .A1(n1121), .A2(n1431), .ZN(n1528) );
  NAND2_X2 U611 ( .A1(n1121), .A2(n1461), .ZN(n1527) );
  MUX2_X1 U612 ( .A(n1529), .B(n1530), .S(n1147), .Z(n1525) );
  NAND2_X2 U613 ( .A1(n1383), .A2(n1111), .ZN(n1530) );
  NAND2_X2 U614 ( .A1(n1391), .A2(n1111), .ZN(n1529) );
  MUX2_X1 U615 ( .A(n1531), .B(n1532), .S(n1141), .Z(n1513) );
  NAND2_X2 U616 ( .A1(n1464), .A2(n1157), .ZN(n1532) );
  NAND2_X2 U617 ( .A1(n1213), .A2(n1156), .ZN(n1531) );
  NAND2_X2 U618 ( .A1(n1533), .A2(n1534), .ZN(B[10]) );
  MUX2_X1 U619 ( .A(n1535), .B(n1536), .S(n1141), .Z(n1534) );
  NAND2_X2 U620 ( .A1(n1159), .A2(n1464), .ZN(n1536) );
  NAND2_X2 U621 ( .A1(n1537), .A2(n1538), .ZN(n1464) );
  MUX2_X1 U622 ( .A(n1539), .B(n1540), .S(n1147), .Z(n1538) );
  NAND2_X2 U623 ( .A1(n1120), .A2(n1370), .ZN(n1540) );
  INV_X2 U624 ( .A(n1541), .ZN(n1370) );
  MUX2_X1 U625 ( .A(n1542), .B(n1266), .S(n1106), .Z(n1541) );
  NAND2_X2 U626 ( .A1(n1120), .A2(n1416), .ZN(n1539) );
  INV_X2 U627 ( .A(n1543), .ZN(n1416) );
  MUX2_X1 U628 ( .A(n1544), .B(n1266), .S(n1106), .Z(n1543) );
  MUX2_X1 U629 ( .A(n1545), .B(n1546), .S(n1147), .Z(n1537) );
  NAND2_X2 U630 ( .A1(n1238), .A2(n1111), .ZN(n1546) );
  INV_X2 U631 ( .A(n1547), .ZN(n1238) );
  MUX2_X1 U632 ( .A(n1548), .B(n1266), .S(n1106), .Z(n1547) );
  NAND2_X2 U633 ( .A1(n1276), .A2(n1111), .ZN(n1545) );
  NAND2_X2 U634 ( .A1(n1158), .A2(n1213), .ZN(n1535) );
  NAND2_X2 U635 ( .A1(n1549), .A2(n1550), .ZN(n1213) );
  MUX2_X1 U636 ( .A(n1551), .B(n1552), .S(n1147), .Z(n1550) );
  NAND2_X2 U637 ( .A1(n1119), .A2(n1445), .ZN(n1552) );
  INV_X2 U638 ( .A(n1553), .ZN(n1445) );
  MUX2_X1 U639 ( .A(n1554), .B(n1266), .S(n1106), .Z(n1553) );
  NAND2_X2 U640 ( .A1(n1119), .A2(n1237), .ZN(n1551) );
  INV_X2 U641 ( .A(n1555), .ZN(n1237) );
  MUX2_X1 U642 ( .A(n1556), .B(n1266), .S(n1106), .Z(n1555) );
  MUX2_X1 U643 ( .A(n1557), .B(n1558), .S(n1147), .Z(n1549) );
  NAND2_X2 U644 ( .A1(n1284), .A2(n1111), .ZN(n1558) );
  NAND2_X2 U645 ( .A1(n1241), .A2(n1111), .ZN(n1557) );
  MUX2_X1 U646 ( .A(n1559), .B(n1560), .S(n1141), .Z(n1533) );
  NAND2_X2 U647 ( .A1(n1193), .A2(n1157), .ZN(n1560) );
  NAND2_X2 U648 ( .A1(n1561), .A2(n1562), .ZN(n1193) );
  MUX2_X1 U649 ( .A(n1563), .B(n1564), .S(n1147), .Z(n1562) );
  NAND2_X2 U650 ( .A1(n1118), .A2(n1405), .ZN(n1564) );
  INV_X2 U651 ( .A(n1565), .ZN(n1405) );
  MUX2_X1 U652 ( .A(n1566), .B(n1266), .S(n1106), .Z(n1565) );
  NAND2_X2 U653 ( .A1(n1118), .A2(n1431), .ZN(n1563) );
  INV_X2 U654 ( .A(n1567), .ZN(n1431) );
  MUX2_X1 U655 ( .A(n1568), .B(n1266), .S(n1106), .Z(n1567) );
  MUX2_X1 U656 ( .A(n1569), .B(n1570), .S(n1147), .Z(n1561) );
  NAND2_X2 U657 ( .A1(n1255), .A2(n1111), .ZN(n1570) );
  INV_X2 U658 ( .A(n1571), .ZN(n1255) );
  MUX2_X1 U659 ( .A(n1572), .B(n1266), .S(n1107), .Z(n1571) );
  NAND2_X2 U660 ( .A1(n1383), .A2(n1111), .ZN(n1569) );
  NAND2_X2 U661 ( .A1(n1194), .A2(n1157), .ZN(n1559) );
  NAND2_X2 U662 ( .A1(n1573), .A2(n1574), .ZN(n1194) );
  MUX2_X1 U663 ( .A(n1575), .B(n1576), .S(n1147), .Z(n1574) );
  NAND2_X2 U664 ( .A1(n1117), .A2(n1461), .ZN(n1576) );
  INV_X2 U665 ( .A(n1577), .ZN(n1461) );
  MUX2_X1 U666 ( .A(n1578), .B(n1266), .S(n1107), .Z(n1577) );
  NAND2_X2 U667 ( .A1(n1117), .A2(n1254), .ZN(n1575) );
  INV_X2 U668 ( .A(n1579), .ZN(n1254) );
  MUX2_X1 U669 ( .A(n1580), .B(n1266), .S(n1107), .Z(n1579) );
  MUX2_X1 U670 ( .A(n1581), .B(n1582), .S(n1146), .Z(n1573) );
  NAND2_X2 U671 ( .A1(n1391), .A2(n1112), .ZN(n1582) );
  NAND2_X2 U672 ( .A1(n1258), .A2(n1112), .ZN(n1581) );
  NAND2_X2 U673 ( .A1(n1583), .A2(n1584), .ZN(B[0]) );
  MUX2_X1 U674 ( .A(n1585), .B(n1586), .S(n1141), .Z(n1584) );
  NAND2_X2 U675 ( .A1(n1158), .A2(n1228), .ZN(n1586) );
  NAND2_X2 U676 ( .A1(n1587), .A2(n1588), .ZN(n1228) );
  MUX2_X1 U677 ( .A(n1589), .B(n1590), .S(n1146), .Z(n1588) );
  NAND2_X2 U678 ( .A1(n1116), .A2(n1276), .ZN(n1590) );
  INV_X2 U679 ( .A(n1591), .ZN(n1276) );
  MUX2_X1 U680 ( .A(n1592), .B(n1266), .S(n1107), .Z(n1591) );
  INV_X2 U681 ( .A(\A[31] ), .ZN(n1266) );
  NAND2_X2 U682 ( .A1(n1116), .A2(n1284), .ZN(n1589) );
  INV_X2 U683 ( .A(n1593), .ZN(n1284) );
  MUX2_X1 U684 ( .A(n1594), .B(n1474), .S(n1107), .Z(n1593) );
  MUX2_X1 U685 ( .A(n1595), .B(n1596), .S(n1146), .Z(n1587) );
  NAND2_X2 U686 ( .A1(n1279), .A2(n1112), .ZN(n1596) );
  INV_X2 U687 ( .A(n1597), .ZN(n1279) );
  MUX2_X1 U688 ( .A(n1598), .B(n1544), .S(n1107), .Z(n1597) );
  NAND2_X2 U689 ( .A1(n1287), .A2(n1112), .ZN(n1595) );
  INV_X2 U690 ( .A(n1599), .ZN(n1287) );
  MUX2_X1 U691 ( .A(n1600), .B(n1554), .S(n1107), .Z(n1599) );
  NAND2_X2 U692 ( .A1(n1173), .A2(n1398), .ZN(n1585) );
  NAND2_X2 U693 ( .A1(n1601), .A2(n1602), .ZN(n1398) );
  MUX2_X1 U694 ( .A(n1603), .B(n1604), .S(n1146), .Z(n1602) );
  NAND2_X2 U695 ( .A1(n1115), .A2(n1241), .ZN(n1604) );
  INV_X2 U696 ( .A(n1605), .ZN(n1241) );
  MUX2_X1 U697 ( .A(n1606), .B(n1502), .S(n1107), .Z(n1605) );
  NAND2_X2 U698 ( .A1(n1115), .A2(n1242), .ZN(n1603) );
  INV_X2 U699 ( .A(n1607), .ZN(n1242) );
  MUX2_X1 U700 ( .A(n1608), .B(n1542), .S(n1107), .Z(n1607) );
  MUX2_X1 U701 ( .A(n1609), .B(n1610), .S(n1147), .Z(n1601) );
  NAND2_X2 U702 ( .A1(n1288), .A2(n1112), .ZN(n1610) );
  INV_X2 U703 ( .A(n1611), .ZN(n1288) );
  MUX2_X1 U704 ( .A(n1612), .B(n1556), .S(n1107), .Z(n1611) );
  NAND2_X2 U705 ( .A1(n1613), .A2(n1112), .ZN(n1609) );
  MUX2_X1 U706 ( .A(A[1]), .B(A[17]), .S(n1107), .Z(n1613) );
  MUX2_X1 U707 ( .A(n1614), .B(n1615), .S(n1142), .Z(n1583) );
  NAND2_X2 U708 ( .A1(n1245), .A2(n1157), .ZN(n1615) );
  NAND2_X2 U709 ( .A1(n1616), .A2(n1617), .ZN(n1245) );
  MUX2_X1 U710 ( .A(n1618), .B(n1619), .S(n1146), .Z(n1617) );
  NAND2_X2 U711 ( .A1(n1114), .A2(n1383), .ZN(n1619) );
  INV_X2 U712 ( .A(n1620), .ZN(n1383) );
  MUX2_X1 U713 ( .A(n1621), .B(n1458), .S(n1107), .Z(n1620) );
  NAND2_X2 U714 ( .A1(n1114), .A2(n1391), .ZN(n1618) );
  INV_X2 U715 ( .A(n1622), .ZN(n1391) );
  MUX2_X1 U716 ( .A(n1623), .B(n1488), .S(n1108), .Z(n1622) );
  MUX2_X1 U717 ( .A(n1624), .B(n1625), .S(n1146), .Z(n1616) );
  NAND2_X2 U718 ( .A1(n1386), .A2(n1112), .ZN(n1625) );
  INV_X2 U719 ( .A(n1626), .ZN(n1386) );
  MUX2_X1 U720 ( .A(n1627), .B(n1568), .S(n1108), .Z(n1626) );
  NAND2_X2 U721 ( .A1(n1394), .A2(n1112), .ZN(n1624) );
  INV_X2 U722 ( .A(n1628), .ZN(n1394) );
  MUX2_X1 U723 ( .A(n1629), .B(n1578), .S(n1108), .Z(n1628) );
  OAI21_X2 U724 ( .B1(n1630), .B2(n1631), .A(n1157), .ZN(n1614) );
  MUX2_X1 U725 ( .A(n1632), .B(n1633), .S(n1146), .Z(n1631) );
  AND2_X2 U726 ( .A1(n1395), .A2(n1112), .ZN(n1633) );
  INV_X2 U727 ( .A(n1634), .ZN(n1395) );
  MUX2_X1 U728 ( .A(n1635), .B(n1580), .S(n1108), .Z(n1634) );
  AND2_X2 U729 ( .A1(n1636), .A2(n1112), .ZN(n1632) );
  MUX2_X1 U730 ( .A(A[0]), .B(A[16]), .S(n1108), .Z(n1636) );
  MUX2_X1 U731 ( .A(n1637), .B(n1638), .S(n1147), .Z(n1630) );
  AND2_X2 U732 ( .A1(n1140), .A2(n1258), .ZN(n1638) );
  INV_X2 U733 ( .A(n1639), .ZN(n1258) );
  MUX2_X1 U734 ( .A(n1640), .B(n1522), .S(n1108), .Z(n1639) );
  AND2_X2 U735 ( .A1(n1140), .A2(n1259), .ZN(n1637) );
  INV_X2 U736 ( .A(n1641), .ZN(n1259) );
  MUX2_X1 U737 ( .A(n1642), .B(n1566), .S(n1108), .Z(n1641) );
endmodule


module up_island_DW_rightsh_1 ( A, SH, B, DATA_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609;

  INV_X1 U174 ( .A(A[18]), .ZN(n585) );
  INV_X1 U175 ( .A(A[15]), .ZN(n572) );
  INV_X1 U176 ( .A(A[19]), .ZN(n583) );
  INV_X1 U177 ( .A(A[20]), .ZN(n581) );
  INV_X1 U178 ( .A(A[21]), .ZN(n579) );
  INV_X1 U179 ( .A(A[9]), .ZN(n438) );
  INV_X1 U180 ( .A(A[10]), .ZN(n584) );
  INV_X1 U181 ( .A(A[22]), .ZN(n575) );
  INV_X1 U182 ( .A(A[23]), .ZN(n573) );
  INV_X1 U183 ( .A(A[8]), .ZN(n486) );
  INV_X1 U184 ( .A(A[16]), .ZN(n487) );
  INV_X1 U185 ( .A(A[17]), .ZN(n439) );
  NAND2_X1 U186 ( .A1(A[28]), .A2(n384), .ZN(n563) );
  INV_X1 U187 ( .A(A[28]), .ZN(n592) );
  NAND2_X1 U188 ( .A1(A[27]), .A2(n385), .ZN(n562) );
  INV_X1 U189 ( .A(A[27]), .ZN(n599) );
  NAND2_X1 U190 ( .A1(A[25]), .A2(n382), .ZN(n503) );
  INV_X1 U191 ( .A(A[25]), .ZN(n601) );
  NAND2_X1 U192 ( .A1(A[30]), .A2(n383), .ZN(n561) );
  INV_X1 U193 ( .A(A[30]), .ZN(n590) );
  INV_X1 U194 ( .A(A[7]), .ZN(n593) );
  INV_X1 U195 ( .A(A[14]), .ZN(n574) );
  INV_X1 U196 ( .A(A[13]), .ZN(n578) );
  INV_X1 U197 ( .A(A[11]), .ZN(n582) );
  INV_X1 U198 ( .A(A[12]), .ZN(n580) );
  NAND2_X1 U199 ( .A1(A[29]), .A2(n384), .ZN(n560) );
  INV_X1 U200 ( .A(A[29]), .ZN(n591) );
  INV_X1 U201 ( .A(A[5]), .ZN(n595) );
  NAND2_X1 U202 ( .A1(A[26]), .A2(n385), .ZN(n504) );
  INV_X1 U203 ( .A(A[26]), .ZN(n600) );
  NAND2_X1 U204 ( .A1(A[24]), .A2(n382), .ZN(n509) );
  INV_X1 U205 ( .A(A[24]), .ZN(n602) );
  INV_X1 U206 ( .A(A[6]), .ZN(n594) );
  INV_X1 U207 ( .A(A[4]), .ZN(n596) );
  INV_X1 U208 ( .A(A[3]), .ZN(n605) );
  INV_X1 U209 ( .A(A[2]), .ZN(n606) );
  INV_X1 U210 ( .A(SH[0]), .ZN(n397) );
  INV_X1 U211 ( .A(A[1]), .ZN(n609) );
  INV_X1 U212 ( .A(SH[4]), .ZN(n378) );
  INV_X1 U213 ( .A(SH[4]), .ZN(n379) );
  INV_X1 U214 ( .A(n386), .ZN(n380) );
  INV_X1 U215 ( .A(n386), .ZN(n381) );
  INV_X1 U216 ( .A(SH[3]), .ZN(n382) );
  INV_X1 U217 ( .A(SH[3]), .ZN(n383) );
  INV_X1 U218 ( .A(SH[3]), .ZN(n384) );
  INV_X1 U219 ( .A(SH[3]), .ZN(n385) );
  INV_X1 U220 ( .A(SH[3]), .ZN(n386) );
  BUF_X1 U221 ( .A(SH[2]), .Z(n387) );
  BUF_X1 U222 ( .A(SH[2]), .Z(n388) );
  INV_X1 U223 ( .A(n393), .ZN(n389) );
  INV_X1 U224 ( .A(n393), .ZN(n390) );
  INV_X1 U225 ( .A(n393), .ZN(n391) );
  INV_X1 U226 ( .A(SH[1]), .ZN(n392) );
  INV_X1 U227 ( .A(SH[1]), .ZN(n393) );
  INV_X1 U228 ( .A(n397), .ZN(n394) );
  INV_X1 U229 ( .A(n397), .ZN(n395) );
  INV_X1 U230 ( .A(n397), .ZN(n396) );
  MUX2_X1 U231 ( .A(n398), .B(n399), .S(n387), .Z(B[9]) );
  MUX2_X1 U232 ( .A(n400), .B(n401), .S(n388), .Z(B[8]) );
  MUX2_X1 U233 ( .A(n402), .B(n403), .S(n388), .Z(B[7]) );
  MUX2_X1 U234 ( .A(n404), .B(n405), .S(n388), .Z(B[6]) );
  MUX2_X1 U235 ( .A(n406), .B(n398), .S(n388), .Z(B[5]) );
  INV_X2 U236 ( .A(n407), .ZN(n398) );
  MUX2_X1 U237 ( .A(n408), .B(n409), .S(SH[4]), .Z(n407) );
  MUX2_X1 U238 ( .A(n410), .B(n411), .S(n389), .Z(n408) );
  MUX2_X1 U239 ( .A(n412), .B(n400), .S(n388), .Z(B[4]) );
  INV_X2 U240 ( .A(n413), .ZN(n400) );
  MUX2_X1 U241 ( .A(n414), .B(n415), .S(SH[4]), .Z(n413) );
  MUX2_X1 U242 ( .A(n416), .B(n417), .S(n389), .Z(n414) );
  MUX2_X1 U243 ( .A(n418), .B(n402), .S(n388), .Z(B[3]) );
  INV_X2 U244 ( .A(n419), .ZN(n402) );
  MUX2_X1 U245 ( .A(n420), .B(n421), .S(SH[4]), .Z(n419) );
  MUX2_X1 U246 ( .A(n422), .B(n410), .S(n389), .Z(n420) );
  MUX2_X1 U247 ( .A(n423), .B(n424), .S(n394), .Z(n410) );
  MUX2_X1 U248 ( .A(n425), .B(n426), .S(SH[4]), .Z(n418) );
  MUX2_X1 U249 ( .A(n427), .B(n428), .S(n389), .Z(n425) );
  INV_X2 U250 ( .A(n429), .ZN(n428) );
  NOR2_X2 U251 ( .A1(n387), .A2(n430), .ZN(B[31]) );
  NOR2_X2 U252 ( .A1(n387), .A2(n431), .ZN(B[30]) );
  MUX2_X1 U253 ( .A(n432), .B(n404), .S(n388), .Z(B[2]) );
  INV_X2 U254 ( .A(n433), .ZN(n404) );
  MUX2_X1 U255 ( .A(n434), .B(n435), .S(SH[4]), .Z(n433) );
  MUX2_X1 U256 ( .A(n436), .B(n416), .S(n389), .Z(n434) );
  MUX2_X1 U257 ( .A(n437), .B(n423), .S(n394), .Z(n416) );
  MUX2_X1 U258 ( .A(n438), .B(n439), .S(n380), .Z(n423) );
  MUX2_X1 U259 ( .A(n440), .B(n441), .S(SH[4]), .Z(n432) );
  MUX2_X1 U260 ( .A(n442), .B(n443), .S(n389), .Z(n440) );
  INV_X2 U261 ( .A(n444), .ZN(n443) );
  NOR2_X2 U262 ( .A1(n387), .A2(n445), .ZN(B[29]) );
  NOR2_X2 U263 ( .A1(n387), .A2(n446), .ZN(B[28]) );
  MUX2_X1 U264 ( .A(n447), .B(n448), .S(n388), .Z(B[27]) );
  INV_X2 U265 ( .A(n430), .ZN(n448) );
  NAND2_X2 U266 ( .A1(n449), .A2(n379), .ZN(n430) );
  INV_X2 U267 ( .A(n450), .ZN(n449) );
  MUX2_X1 U268 ( .A(n451), .B(n452), .S(n388), .Z(B[26]) );
  INV_X2 U269 ( .A(n431), .ZN(n452) );
  NAND2_X2 U270 ( .A1(n453), .A2(n379), .ZN(n431) );
  INV_X2 U271 ( .A(n454), .ZN(n453) );
  MUX2_X1 U272 ( .A(n455), .B(n456), .S(n388), .Z(B[25]) );
  INV_X2 U273 ( .A(n445), .ZN(n456) );
  NAND2_X2 U274 ( .A1(n457), .A2(n379), .ZN(n445) );
  INV_X2 U275 ( .A(n458), .ZN(n457) );
  MUX2_X1 U276 ( .A(n459), .B(n460), .S(n388), .Z(B[24]) );
  INV_X2 U277 ( .A(n446), .ZN(n460) );
  NAND2_X2 U278 ( .A1(n461), .A2(n379), .ZN(n446) );
  INV_X2 U279 ( .A(n462), .ZN(n461) );
  MUX2_X1 U280 ( .A(n463), .B(n447), .S(n388), .Z(B[23]) );
  INV_X2 U281 ( .A(n464), .ZN(n447) );
  NAND2_X2 U282 ( .A1(n465), .A2(n378), .ZN(n464) );
  INV_X2 U283 ( .A(n466), .ZN(n465) );
  MUX2_X1 U284 ( .A(n467), .B(n451), .S(n388), .Z(B[22]) );
  INV_X2 U285 ( .A(n468), .ZN(n451) );
  NAND2_X2 U286 ( .A1(n469), .A2(n378), .ZN(n468) );
  INV_X2 U287 ( .A(n470), .ZN(n469) );
  MUX2_X1 U288 ( .A(n471), .B(n455), .S(n388), .Z(B[21]) );
  INV_X2 U289 ( .A(n472), .ZN(n455) );
  NAND2_X2 U290 ( .A1(n473), .A2(n378), .ZN(n472) );
  INV_X2 U291 ( .A(n409), .ZN(n473) );
  MUX2_X1 U292 ( .A(n474), .B(n475), .S(n389), .Z(n409) );
  MUX2_X1 U293 ( .A(n476), .B(n459), .S(n388), .Z(B[20]) );
  INV_X2 U294 ( .A(n477), .ZN(n459) );
  NAND2_X2 U295 ( .A1(n478), .A2(n378), .ZN(n477) );
  INV_X2 U296 ( .A(n415), .ZN(n478) );
  MUX2_X1 U297 ( .A(n479), .B(n480), .S(n389), .Z(n415) );
  MUX2_X1 U298 ( .A(n481), .B(n406), .S(n388), .Z(B[1]) );
  INV_X2 U299 ( .A(n482), .ZN(n406) );
  MUX2_X1 U300 ( .A(n483), .B(n484), .S(SH[4]), .Z(n482) );
  MUX2_X1 U301 ( .A(n429), .B(n422), .S(n389), .Z(n483) );
  MUX2_X1 U302 ( .A(n485), .B(n437), .S(n394), .Z(n422) );
  MUX2_X1 U303 ( .A(n486), .B(n487), .S(n380), .Z(n437) );
  MUX2_X1 U304 ( .A(n488), .B(n489), .S(n394), .Z(n429) );
  MUX2_X1 U305 ( .A(n490), .B(n491), .S(SH[4]), .Z(n481) );
  MUX2_X1 U306 ( .A(n492), .B(n427), .S(n389), .Z(n490) );
  INV_X2 U307 ( .A(n493), .ZN(n427) );
  MUX2_X1 U308 ( .A(n494), .B(n495), .S(n394), .Z(n493) );
  MUX2_X1 U309 ( .A(n496), .B(n497), .S(n394), .Z(n492) );
  INV_X2 U310 ( .A(n498), .ZN(n497) );
  MUX2_X1 U311 ( .A(n499), .B(n463), .S(n387), .Z(B[19]) );
  INV_X2 U312 ( .A(n500), .ZN(n463) );
  NAND2_X2 U313 ( .A1(n501), .A2(n378), .ZN(n500) );
  INV_X2 U314 ( .A(n421), .ZN(n501) );
  MUX2_X1 U315 ( .A(n502), .B(n474), .S(n389), .Z(n421) );
  MUX2_X1 U316 ( .A(n503), .B(n504), .S(n394), .Z(n474) );
  MUX2_X1 U317 ( .A(n505), .B(n467), .S(n387), .Z(B[18]) );
  INV_X2 U318 ( .A(n506), .ZN(n467) );
  NAND2_X2 U319 ( .A1(n507), .A2(n378), .ZN(n506) );
  INV_X2 U320 ( .A(n435), .ZN(n507) );
  MUX2_X1 U321 ( .A(n508), .B(n479), .S(n389), .Z(n435) );
  MUX2_X1 U322 ( .A(n509), .B(n503), .S(n394), .Z(n479) );
  MUX2_X1 U323 ( .A(n510), .B(n471), .S(n387), .Z(B[17]) );
  INV_X2 U324 ( .A(n511), .ZN(n471) );
  NAND2_X2 U325 ( .A1(n512), .A2(n378), .ZN(n511) );
  INV_X2 U326 ( .A(n484), .ZN(n512) );
  MUX2_X1 U327 ( .A(n513), .B(n502), .S(n390), .Z(n484) );
  MUX2_X1 U328 ( .A(n514), .B(n509), .S(n394), .Z(n502) );
  MUX2_X1 U329 ( .A(n515), .B(n476), .S(n387), .Z(B[16]) );
  INV_X2 U330 ( .A(n516), .ZN(n476) );
  NAND2_X2 U331 ( .A1(n517), .A2(n378), .ZN(n516) );
  INV_X2 U332 ( .A(n518), .ZN(n517) );
  MUX2_X1 U333 ( .A(n519), .B(n499), .S(n387), .Z(B[15]) );
  INV_X2 U334 ( .A(n520), .ZN(n499) );
  NAND2_X2 U335 ( .A1(n426), .A2(n378), .ZN(n520) );
  INV_X2 U336 ( .A(n521), .ZN(n426) );
  MUX2_X1 U337 ( .A(n522), .B(n513), .S(n390), .Z(n521) );
  MUX2_X1 U338 ( .A(n523), .B(n524), .S(n394), .Z(n513) );
  MUX2_X1 U339 ( .A(n525), .B(n505), .S(n387), .Z(B[14]) );
  INV_X2 U340 ( .A(n526), .ZN(n505) );
  NAND2_X2 U341 ( .A1(n441), .A2(n378), .ZN(n526) );
  INV_X2 U342 ( .A(n527), .ZN(n441) );
  MUX2_X1 U343 ( .A(n528), .B(n529), .S(n390), .Z(n527) );
  MUX2_X1 U344 ( .A(n399), .B(n510), .S(n387), .Z(B[13]) );
  INV_X2 U345 ( .A(n530), .ZN(n510) );
  NAND2_X2 U346 ( .A1(n491), .A2(n378), .ZN(n530) );
  INV_X2 U347 ( .A(n531), .ZN(n491) );
  MUX2_X1 U348 ( .A(n532), .B(n522), .S(n390), .Z(n531) );
  MUX2_X1 U349 ( .A(n533), .B(n534), .S(n394), .Z(n522) );
  INV_X2 U350 ( .A(n535), .ZN(n399) );
  MUX2_X1 U351 ( .A(n536), .B(n458), .S(SH[4]), .Z(n535) );
  MUX2_X1 U352 ( .A(n537), .B(n538), .S(n390), .Z(n458) );
  MUX2_X1 U353 ( .A(n539), .B(n540), .S(n390), .Z(n536) );
  MUX2_X1 U354 ( .A(n401), .B(n515), .S(n387), .Z(B[12]) );
  INV_X2 U355 ( .A(n541), .ZN(n515) );
  NAND2_X2 U356 ( .A1(n542), .A2(n378), .ZN(n541) );
  INV_X2 U357 ( .A(n543), .ZN(n401) );
  MUX2_X1 U358 ( .A(n544), .B(n462), .S(SH[4]), .Z(n543) );
  MUX2_X1 U359 ( .A(n545), .B(n546), .S(n390), .Z(n462) );
  MUX2_X1 U360 ( .A(n547), .B(n548), .S(n390), .Z(n544) );
  MUX2_X1 U361 ( .A(n403), .B(n519), .S(n387), .Z(B[11]) );
  INV_X2 U362 ( .A(n549), .ZN(n519) );
  MUX2_X1 U363 ( .A(n550), .B(n450), .S(SH[4]), .Z(n549) );
  NAND2_X2 U364 ( .A1(n551), .A2(n392), .ZN(n450) );
  INV_X2 U365 ( .A(n538), .ZN(n551) );
  NAND2_X2 U366 ( .A1(n552), .A2(n397), .ZN(n538) );
  INV_X2 U367 ( .A(n553), .ZN(n552) );
  MUX2_X1 U368 ( .A(n540), .B(n532), .S(n390), .Z(n550) );
  MUX2_X1 U369 ( .A(n554), .B(n555), .S(n394), .Z(n532) );
  MUX2_X1 U370 ( .A(n556), .B(n557), .S(n395), .Z(n540) );
  INV_X2 U371 ( .A(n558), .ZN(n403) );
  MUX2_X1 U372 ( .A(n559), .B(n466), .S(SH[4]), .Z(n558) );
  MUX2_X1 U373 ( .A(n475), .B(n537), .S(n390), .Z(n466) );
  MUX2_X1 U374 ( .A(n560), .B(n561), .S(n395), .Z(n537) );
  MUX2_X1 U375 ( .A(n562), .B(n563), .S(n395), .Z(n475) );
  MUX2_X1 U376 ( .A(n411), .B(n539), .S(n390), .Z(n559) );
  MUX2_X1 U377 ( .A(n564), .B(n565), .S(n395), .Z(n539) );
  MUX2_X1 U378 ( .A(n566), .B(n567), .S(n395), .Z(n411) );
  MUX2_X1 U379 ( .A(n405), .B(n525), .S(n387), .Z(B[10]) );
  INV_X2 U380 ( .A(n568), .ZN(n525) );
  MUX2_X1 U381 ( .A(n569), .B(n454), .S(SH[4]), .Z(n568) );
  NAND2_X2 U382 ( .A1(n570), .A2(n392), .ZN(n454) );
  INV_X2 U383 ( .A(n546), .ZN(n570) );
  MUX2_X1 U384 ( .A(n561), .B(n553), .S(n395), .Z(n546) );
  NAND2_X2 U385 ( .A1(A[31]), .A2(n383), .ZN(n553) );
  MUX2_X1 U386 ( .A(n548), .B(n571), .S(n390), .Z(n569) );
  MUX2_X1 U387 ( .A(n565), .B(n556), .S(n395), .Z(n548) );
  MUX2_X1 U388 ( .A(n572), .B(n573), .S(n380), .Z(n556) );
  MUX2_X1 U389 ( .A(n574), .B(n575), .S(n380), .Z(n565) );
  INV_X2 U390 ( .A(n576), .ZN(n405) );
  MUX2_X1 U391 ( .A(n577), .B(n470), .S(SH[4]), .Z(n576) );
  MUX2_X1 U392 ( .A(n480), .B(n545), .S(n391), .Z(n470) );
  MUX2_X1 U393 ( .A(n563), .B(n560), .S(n395), .Z(n545) );
  MUX2_X1 U394 ( .A(n504), .B(n562), .S(n395), .Z(n480) );
  MUX2_X1 U395 ( .A(n417), .B(n547), .S(n391), .Z(n577) );
  MUX2_X1 U396 ( .A(n567), .B(n564), .S(n395), .Z(n547) );
  MUX2_X1 U397 ( .A(n578), .B(n579), .S(n380), .Z(n564) );
  MUX2_X1 U398 ( .A(n580), .B(n581), .S(n380), .Z(n567) );
  MUX2_X1 U399 ( .A(n424), .B(n566), .S(n395), .Z(n417) );
  MUX2_X1 U400 ( .A(n582), .B(n583), .S(n380), .Z(n566) );
  MUX2_X1 U401 ( .A(n584), .B(n585), .S(n380), .Z(n424) );
  MUX2_X1 U402 ( .A(n586), .B(n412), .S(n388), .Z(B[0]) );
  INV_X2 U403 ( .A(n587), .ZN(n412) );
  MUX2_X1 U404 ( .A(n588), .B(n518), .S(SH[4]), .Z(n587) );
  MUX2_X1 U405 ( .A(n529), .B(n508), .S(n391), .Z(n518) );
  MUX2_X1 U406 ( .A(n524), .B(n514), .S(n395), .Z(n508) );
  MUX2_X1 U407 ( .A(n573), .B(n589), .S(n380), .Z(n514) );
  INV_X2 U408 ( .A(A[31]), .ZN(n589) );
  MUX2_X1 U409 ( .A(n575), .B(n590), .S(n380), .Z(n524) );
  MUX2_X1 U410 ( .A(n534), .B(n523), .S(n396), .Z(n529) );
  MUX2_X1 U411 ( .A(n579), .B(n591), .S(n380), .Z(n523) );
  MUX2_X1 U412 ( .A(n581), .B(n592), .S(n380), .Z(n534) );
  MUX2_X1 U413 ( .A(n444), .B(n436), .S(n391), .Z(n588) );
  MUX2_X1 U414 ( .A(n489), .B(n485), .S(n396), .Z(n436) );
  MUX2_X1 U415 ( .A(n593), .B(n572), .S(n381), .Z(n485) );
  MUX2_X1 U416 ( .A(n594), .B(n574), .S(n381), .Z(n489) );
  MUX2_X1 U417 ( .A(n495), .B(n488), .S(n396), .Z(n444) );
  MUX2_X1 U418 ( .A(n595), .B(n578), .S(n381), .Z(n488) );
  MUX2_X1 U419 ( .A(n596), .B(n580), .S(n381), .Z(n495) );
  MUX2_X1 U420 ( .A(n597), .B(n542), .S(SH[4]), .Z(n586) );
  INV_X2 U421 ( .A(n598), .ZN(n542) );
  MUX2_X1 U422 ( .A(n571), .B(n528), .S(n391), .Z(n598) );
  MUX2_X1 U423 ( .A(n555), .B(n533), .S(n396), .Z(n528) );
  MUX2_X1 U424 ( .A(n583), .B(n599), .S(n381), .Z(n533) );
  MUX2_X1 U425 ( .A(n585), .B(n600), .S(n381), .Z(n555) );
  MUX2_X1 U426 ( .A(n557), .B(n554), .S(n396), .Z(n571) );
  MUX2_X1 U427 ( .A(n439), .B(n601), .S(n381), .Z(n554) );
  MUX2_X1 U428 ( .A(n487), .B(n602), .S(n381), .Z(n557) );
  MUX2_X1 U429 ( .A(n603), .B(n442), .S(n391), .Z(n597) );
  INV_X2 U430 ( .A(n604), .ZN(n442) );
  MUX2_X1 U431 ( .A(n498), .B(n494), .S(n396), .Z(n604) );
  MUX2_X1 U432 ( .A(n605), .B(n582), .S(n381), .Z(n494) );
  MUX2_X1 U433 ( .A(n606), .B(n584), .S(n381), .Z(n498) );
  MUX2_X1 U434 ( .A(n607), .B(n496), .S(n396), .Z(n603) );
  INV_X2 U435 ( .A(n608), .ZN(n496) );
  MUX2_X1 U436 ( .A(n609), .B(n438), .S(n381), .Z(n608) );
  MUX2_X1 U437 ( .A(A[0]), .B(A[8]), .S(n381), .Z(n607) );
endmodule


module up_island_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n8, n9, n10, n14, n15, n19, n24, n25, n26, n30, n31, n35, n40, n50,
         n60, n82, n83, n87, n92, n93, n94, n98, n99, n103, n108, n109, n110,
         n114, n115, n119, n124, n125, n126, n130, n131, n135, n140, n141,
         n142, n146, n147, n151, n156, n157, n158, n162, n163, n167, n172,
         n173, n174, n178, n179, n183, n188, n189, n190, n194, n195, n199,
         n204, n205, n206, n210, n211, n215, n220, n221, n222, n226, n227,
         n231, n236, n237, n238, n242, n243, n247, n252, n253, n254, n258,
         n259, n263, n268, n269, n270, n274, n275, n279, n284, n285, n286,
         n290, n291, n295, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170;

  NAND2_X2 OR_NOTi ( .A1(n295), .A2(n299), .ZN(n3058) );
  INV_X4 U1 ( .A(n441), .ZN(n295) );
  NAND2_X2 AND_NOTi ( .A1(n441), .A2(n290), .ZN(n291) );
  INV_X4 U2 ( .A(n291), .ZN(product[0]) );
  INV_X4 U11 ( .A(n347), .ZN(n290) );
  OAI21_X2 AO21i ( .B1(n284), .B2(n285), .A(n286), .ZN(n2499) );
  INV_X4 U3 ( .A(n3026), .ZN(n286) );
  INV_X4 U21 ( .A(n347), .ZN(n285) );
  INV_X4 U12 ( .A(n395), .ZN(n284) );
  NAND2_X2 OR_NOTi1 ( .A1(n279), .A2(n302), .ZN(n3025) );
  INV_X4 U13 ( .A(n441), .ZN(n279) );
  NAND2_X2 AND_NOTi1 ( .A1(n441), .A2(n274), .ZN(n275) );
  INV_X4 U22 ( .A(n275), .ZN(n2498) );
  INV_X4 U14 ( .A(n350), .ZN(n274) );
  OAI21_X2 AO21i1 ( .B1(n268), .B2(n269), .A(n270), .ZN(n2467) );
  INV_X4 U31 ( .A(n2993), .ZN(n270) );
  INV_X4 U23 ( .A(n350), .ZN(n269) );
  INV_X4 U15 ( .A(n398), .ZN(n268) );
  NAND2_X2 OR_NOTi2 ( .A1(n263), .A2(n305), .ZN(n2992) );
  INV_X4 U16 ( .A(n441), .ZN(n263) );
  NAND2_X2 AND_NOTi2 ( .A1(n441), .A2(n258), .ZN(n259) );
  INV_X4 U24 ( .A(n259), .ZN(n2466) );
  INV_X4 U17 ( .A(n353), .ZN(n258) );
  OAI21_X2 AO21i2 ( .B1(n252), .B2(n253), .A(n254), .ZN(n2435) );
  INV_X4 U32 ( .A(n2960), .ZN(n254) );
  INV_X4 U25 ( .A(n353), .ZN(n253) );
  INV_X4 U18 ( .A(n401), .ZN(n252) );
  NAND2_X2 OR_NOTi3 ( .A1(n247), .A2(n308), .ZN(n2959) );
  INV_X4 U19 ( .A(n441), .ZN(n247) );
  NAND2_X2 AND_NOTi3 ( .A1(n441), .A2(n242), .ZN(n243) );
  INV_X4 U26 ( .A(n243), .ZN(n2434) );
  INV_X4 U110 ( .A(n356), .ZN(n242) );
  OAI21_X2 AO21i3 ( .B1(n236), .B2(n237), .A(n238), .ZN(n2403) );
  INV_X4 U33 ( .A(n2927), .ZN(n238) );
  INV_X4 U27 ( .A(n356), .ZN(n237) );
  INV_X4 U111 ( .A(n404), .ZN(n236) );
  NAND2_X2 OR_NOTi4 ( .A1(n231), .A2(n311), .ZN(n2926) );
  INV_X4 U112 ( .A(n441), .ZN(n231) );
  NAND2_X2 AND_NOTi4 ( .A1(n441), .A2(n226), .ZN(n227) );
  INV_X4 U28 ( .A(n227), .ZN(n2402) );
  INV_X4 U113 ( .A(n359), .ZN(n226) );
  OAI21_X2 AO21i4 ( .B1(n220), .B2(n221), .A(n222), .ZN(n2371) );
  INV_X4 U34 ( .A(n2894), .ZN(n222) );
  INV_X4 U29 ( .A(n359), .ZN(n221) );
  INV_X4 U114 ( .A(n407), .ZN(n220) );
  NAND2_X2 OR_NOTi5 ( .A1(n215), .A2(n314), .ZN(n2893) );
  INV_X4 U115 ( .A(n441), .ZN(n215) );
  NAND2_X2 AND_NOTi5 ( .A1(n441), .A2(n210), .ZN(n211) );
  INV_X4 U210 ( .A(n211), .ZN(n2370) );
  INV_X4 U116 ( .A(n362), .ZN(n210) );
  OAI21_X2 AO21i5 ( .B1(n204), .B2(n205), .A(n206), .ZN(n2339) );
  INV_X4 U35 ( .A(n2861), .ZN(n206) );
  INV_X4 U211 ( .A(n362), .ZN(n205) );
  INV_X4 U117 ( .A(n410), .ZN(n204) );
  NAND2_X2 OR_NOTi6 ( .A1(n199), .A2(n317), .ZN(n2860) );
  INV_X4 U118 ( .A(n441), .ZN(n199) );
  NAND2_X2 AND_NOTi6 ( .A1(n441), .A2(n194), .ZN(n195) );
  INV_X4 U212 ( .A(n195), .ZN(n2338) );
  INV_X4 U119 ( .A(n365), .ZN(n194) );
  OAI21_X2 AO21i6 ( .B1(n188), .B2(n189), .A(n190), .ZN(n2307) );
  INV_X4 U36 ( .A(n2828), .ZN(n190) );
  INV_X4 U213 ( .A(n365), .ZN(n189) );
  INV_X4 U120 ( .A(n413), .ZN(n188) );
  NAND2_X2 OR_NOTi7 ( .A1(n183), .A2(n320), .ZN(n2827) );
  INV_X4 U121 ( .A(n441), .ZN(n183) );
  NAND2_X2 AND_NOTi7 ( .A1(n441), .A2(n178), .ZN(n179) );
  INV_X4 U214 ( .A(n179), .ZN(n2306) );
  INV_X4 U122 ( .A(n368), .ZN(n178) );
  OAI21_X2 AO21i7 ( .B1(n172), .B2(n173), .A(n174), .ZN(n2275) );
  INV_X4 U37 ( .A(n2795), .ZN(n174) );
  INV_X4 U215 ( .A(n368), .ZN(n173) );
  INV_X4 U123 ( .A(n416), .ZN(n172) );
  NAND2_X2 OR_NOTi8 ( .A1(n167), .A2(n323), .ZN(n2794) );
  INV_X4 U124 ( .A(n441), .ZN(n167) );
  NAND2_X2 AND_NOTi8 ( .A1(n441), .A2(n162), .ZN(n163) );
  INV_X4 U216 ( .A(n163), .ZN(n2274) );
  INV_X4 U125 ( .A(n371), .ZN(n162) );
  OAI21_X2 AO21i8 ( .B1(n156), .B2(n157), .A(n158), .ZN(n2243) );
  INV_X4 U38 ( .A(n2762), .ZN(n158) );
  INV_X4 U217 ( .A(n371), .ZN(n157) );
  INV_X4 U126 ( .A(n419), .ZN(n156) );
  NAND2_X2 OR_NOTi9 ( .A1(n151), .A2(n326), .ZN(n2761) );
  INV_X4 U127 ( .A(n441), .ZN(n151) );
  NAND2_X2 AND_NOTi9 ( .A1(n441), .A2(n146), .ZN(n147) );
  INV_X4 U218 ( .A(n147), .ZN(n2242) );
  INV_X4 U128 ( .A(n374), .ZN(n146) );
  OAI21_X2 AO21i9 ( .B1(n140), .B2(n141), .A(n142), .ZN(n2211) );
  INV_X4 U39 ( .A(n2729), .ZN(n142) );
  INV_X4 U219 ( .A(n374), .ZN(n141) );
  INV_X4 U129 ( .A(n422), .ZN(n140) );
  NAND2_X2 OR_NOTi10 ( .A1(n135), .A2(n329), .ZN(n2728) );
  INV_X4 U130 ( .A(n441), .ZN(n135) );
  NAND2_X2 AND_NOTi10 ( .A1(n441), .A2(n130), .ZN(n131) );
  INV_X4 U220 ( .A(n131), .ZN(n2210) );
  INV_X4 U131 ( .A(n377), .ZN(n130) );
  OAI21_X2 AO21i10 ( .B1(n124), .B2(n125), .A(n126), .ZN(n2179) );
  INV_X4 U310 ( .A(n2696), .ZN(n126) );
  INV_X4 U221 ( .A(n377), .ZN(n125) );
  INV_X4 U132 ( .A(n425), .ZN(n124) );
  NAND2_X2 OR_NOTi11 ( .A1(n119), .A2(n332), .ZN(n2695) );
  INV_X4 U133 ( .A(n441), .ZN(n119) );
  NAND2_X2 AND_NOTi11 ( .A1(n441), .A2(n114), .ZN(n115) );
  INV_X4 U222 ( .A(n115), .ZN(n2178) );
  INV_X4 U134 ( .A(n380), .ZN(n114) );
  OAI21_X2 AO21i11 ( .B1(n108), .B2(n109), .A(n110), .ZN(n2147) );
  INV_X4 U311 ( .A(n2663), .ZN(n110) );
  INV_X4 U223 ( .A(n380), .ZN(n109) );
  INV_X4 U135 ( .A(n428), .ZN(n108) );
  NAND2_X2 OR_NOTi12 ( .A1(n103), .A2(n335), .ZN(n2662) );
  INV_X4 U136 ( .A(n441), .ZN(n103) );
  NAND2_X2 AND_NOTi12 ( .A1(n441), .A2(n98), .ZN(n99) );
  INV_X4 U224 ( .A(n99), .ZN(n2146) );
  INV_X4 U137 ( .A(n383), .ZN(n98) );
  OAI21_X2 AO21i12 ( .B1(n92), .B2(n93), .A(n94), .ZN(n2115) );
  INV_X4 U312 ( .A(n2630), .ZN(n94) );
  INV_X4 U225 ( .A(n383), .ZN(n93) );
  INV_X4 U138 ( .A(n431), .ZN(n92) );
  NAND2_X2 OR_NOTi13 ( .A1(n87), .A2(n338), .ZN(n2629) );
  INV_X4 U139 ( .A(n441), .ZN(n87) );
  NAND2_X2 AND_NOTi13 ( .A1(n441), .A2(n82), .ZN(n83) );
  INV_X4 U226 ( .A(n83), .ZN(n2114) );
  INV_X4 U140 ( .A(n386), .ZN(n82) );
  OAI21_X2 AO21i13 ( .B1(n40), .B2(n50), .A(n60), .ZN(n2083) );
  INV_X4 U313 ( .A(n2597), .ZN(n60) );
  INV_X4 U227 ( .A(n386), .ZN(n50) );
  INV_X4 U141 ( .A(n434), .ZN(n40) );
  NAND2_X2 OR_NOTi14 ( .A1(n35), .A2(n341), .ZN(n2596) );
  INV_X4 U142 ( .A(n441), .ZN(n35) );
  NAND2_X2 AND_NOTi14 ( .A1(n441), .A2(n30), .ZN(n31) );
  INV_X4 U228 ( .A(n31), .ZN(n2082) );
  INV_X4 U143 ( .A(n389), .ZN(n30) );
  OAI21_X2 AO21i14 ( .B1(n24), .B2(n25), .A(n26), .ZN(n2051) );
  INV_X4 U314 ( .A(n2564), .ZN(n26) );
  INV_X4 U229 ( .A(n389), .ZN(n25) );
  INV_X4 U144 ( .A(n437), .ZN(n24) );
  NAND2_X2 OR_NOTi15 ( .A1(n19), .A2(n342), .ZN(n2563) );
  INV_X4 U145 ( .A(n441), .ZN(n19) );
  NAND2_X2 AND_NOTi15 ( .A1(n441), .A2(n14), .ZN(n15) );
  INV_X4 U230 ( .A(n15), .ZN(n2050) );
  INV_X4 U146 ( .A(n392), .ZN(n14) );
  OAI21_X2 AO21i15 ( .B1(n8), .B2(n9), .A(n10), .ZN(n2019) );
  INV_X4 U315 ( .A(n2531), .ZN(n10) );
  INV_X4 U231 ( .A(n392), .ZN(n9) );
  INV_X4 U147 ( .A(n440), .ZN(n8) );
  BUF_X32 U4 ( .A(n3170), .Z(n297) );
  BUF_X32 U5 ( .A(n3170), .Z(n298) );
  BUF_X32 U6 ( .A(n3170), .Z(n299) );
  BUF_X32 U7 ( .A(n3169), .Z(n300) );
  BUF_X32 U8 ( .A(n3169), .Z(n301) );
  BUF_X32 U9 ( .A(n3169), .Z(n302) );
  BUF_X32 U10 ( .A(n3168), .Z(n303) );
  BUF_X32 U20 ( .A(n3168), .Z(n304) );
  BUF_X32 U30 ( .A(n3168), .Z(n305) );
  BUF_X32 U40 ( .A(n3167), .Z(n306) );
  BUF_X32 U41 ( .A(n3167), .Z(n307) );
  BUF_X32 U42 ( .A(n3167), .Z(n308) );
  BUF_X32 U43 ( .A(n3166), .Z(n309) );
  BUF_X32 U44 ( .A(n3166), .Z(n310) );
  BUF_X32 U45 ( .A(n3166), .Z(n311) );
  BUF_X32 U46 ( .A(n3165), .Z(n312) );
  BUF_X32 U47 ( .A(n3165), .Z(n313) );
  BUF_X32 U48 ( .A(n3165), .Z(n314) );
  BUF_X32 U49 ( .A(n3164), .Z(n315) );
  BUF_X32 U50 ( .A(n3164), .Z(n316) );
  BUF_X32 U51 ( .A(n3164), .Z(n317) );
  BUF_X32 U52 ( .A(n3163), .Z(n318) );
  BUF_X32 U53 ( .A(n3163), .Z(n319) );
  BUF_X32 U54 ( .A(n3163), .Z(n320) );
  BUF_X32 U55 ( .A(n3162), .Z(n321) );
  BUF_X32 U56 ( .A(n3162), .Z(n322) );
  BUF_X32 U57 ( .A(n3162), .Z(n323) );
  BUF_X32 U58 ( .A(n3161), .Z(n324) );
  BUF_X32 U59 ( .A(n3161), .Z(n325) );
  BUF_X32 U60 ( .A(n3161), .Z(n326) );
  BUF_X32 U61 ( .A(n3160), .Z(n327) );
  BUF_X32 U62 ( .A(n3160), .Z(n328) );
  BUF_X32 U63 ( .A(n3160), .Z(n329) );
  BUF_X32 U64 ( .A(n3159), .Z(n330) );
  BUF_X32 U65 ( .A(n3159), .Z(n331) );
  BUF_X32 U66 ( .A(n3159), .Z(n332) );
  BUF_X32 U67 ( .A(n3158), .Z(n333) );
  BUF_X32 U68 ( .A(n3158), .Z(n334) );
  BUF_X32 U69 ( .A(n3158), .Z(n335) );
  BUF_X32 U70 ( .A(n3157), .Z(n336) );
  BUF_X32 U71 ( .A(n3157), .Z(n337) );
  BUF_X32 U72 ( .A(n3157), .Z(n338) );
  BUF_X32 U73 ( .A(n3156), .Z(n339) );
  BUF_X32 U74 ( .A(n3156), .Z(n340) );
  BUF_X32 U75 ( .A(n3156), .Z(n341) );
  BUF_X32 U76 ( .A(a[31]), .Z(n342) );
  BUF_X32 U79 ( .A(n3138), .Z(n345) );
  BUF_X32 U80 ( .A(n3138), .Z(n346) );
  BUF_X32 U81 ( .A(n3138), .Z(n347) );
  BUF_X32 U165 ( .A(n3122), .Z(n393) );
  BUF_X32 U166 ( .A(n3122), .Z(n394) );
  BUF_X32 U167 ( .A(n3122), .Z(n395) );
  BUF_X32 U168 ( .A(n3121), .Z(n396) );
  BUF_X32 U169 ( .A(n3121), .Z(n397) );
  BUF_X32 U171 ( .A(n3120), .Z(n399) );
  BUF_X32 U172 ( .A(n3120), .Z(n400) );
  BUF_X32 U174 ( .A(n3119), .Z(n402) );
  BUF_X32 U175 ( .A(n3119), .Z(n403) );
  BUF_X32 U177 ( .A(n3118), .Z(n405) );
  BUF_X32 U178 ( .A(n3118), .Z(n406) );
  BUF_X32 U180 ( .A(n3117), .Z(n408) );
  BUF_X32 U181 ( .A(n3117), .Z(n409) );
  BUF_X32 U183 ( .A(n3116), .Z(n411) );
  BUF_X32 U184 ( .A(n3116), .Z(n412) );
  BUF_X32 U186 ( .A(n3115), .Z(n414) );
  BUF_X32 U187 ( .A(n3115), .Z(n415) );
  BUF_X32 U189 ( .A(n3114), .Z(n417) );
  BUF_X32 U190 ( .A(n3114), .Z(n418) );
  BUF_X32 U192 ( .A(n3113), .Z(n420) );
  BUF_X32 U193 ( .A(n3113), .Z(n421) );
  BUF_X32 U195 ( .A(n3112), .Z(n423) );
  BUF_X32 U196 ( .A(n3112), .Z(n424) );
  BUF_X32 U198 ( .A(n3111), .Z(n426) );
  BUF_X32 U199 ( .A(n3111), .Z(n427) );
  BUF_X32 U201 ( .A(n3110), .Z(n429) );
  BUF_X32 U202 ( .A(n3110), .Z(n430) );
  BUF_X32 U204 ( .A(n3109), .Z(n432) );
  BUF_X32 U205 ( .A(n3109), .Z(n433) );
  BUF_X32 U207 ( .A(n3108), .Z(n435) );
  BUF_X32 U208 ( .A(n3108), .Z(n436) );
  BUF_X32 U232 ( .A(n3107), .Z(n438) );
  BUF_X32 U233 ( .A(n3107), .Z(n439) );
  BUF_X32 U235 ( .A(b[0]), .Z(n441) );
  BUF_X32 U238 ( .A(n765), .Z(n444) );
  BUF_X32 U239 ( .A(n765), .Z(n445) );
  BUF_X32 U240 ( .A(n683), .Z(n446) );
  BUF_X32 U241 ( .A(n682), .Z(n447) );
  INV_X32 U242 ( .A(n510), .ZN(product[63]) );
  XNOR2_X2 U243 ( .A(n517), .B(n448), .ZN(product[62]) );
  OAI21_X4 U244 ( .B1(n445), .B2(n511), .A(n512), .ZN(n510) );
  NAND2_X4 U245 ( .A1(n520), .A2(n513), .ZN(n511) );
  AOI21_X4 U246 ( .B1(n521), .B2(n513), .A(n514), .ZN(n512) );
  INV_X4 U247 ( .A(n515), .ZN(n513) );
  INV_X4 U248 ( .A(n516), .ZN(n514) );
  NAND2_X4 U249 ( .A1(n1011), .A2(n516), .ZN(n448) );
  INV_X32 U250 ( .A(n515), .ZN(n1011) );
  NOR2_X4 U251 ( .A1(n2019), .A2(n1073), .ZN(n515) );
  NAND2_X4 U252 ( .A1(n2019), .A2(n1073), .ZN(n516) );
  XNOR2_X2 U253 ( .A(n528), .B(n449), .ZN(product[61]) );
  OAI21_X4 U254 ( .B1(n445), .B2(n518), .A(n519), .ZN(n517) );
  INV_X4 U255 ( .A(n520), .ZN(n518) );
  INV_X4 U256 ( .A(n521), .ZN(n519) );
  NOR2_X4 U257 ( .A1(n447), .A2(n522), .ZN(n520) );
  OAI21_X4 U258 ( .B1(n446), .B2(n522), .A(n523), .ZN(n521) );
  NAND2_X4 U259 ( .A1(n533), .A2(n524), .ZN(n522) );
  AOI21_X4 U260 ( .B1(n534), .B2(n524), .A(n525), .ZN(n523) );
  INV_X4 U261 ( .A(n526), .ZN(n524) );
  INV_X4 U262 ( .A(n527), .ZN(n525) );
  NAND2_X4 U263 ( .A1(n1012), .A2(n527), .ZN(n449) );
  INV_X32 U264 ( .A(n526), .ZN(n1012) );
  NOR2_X4 U265 ( .A1(n1075), .A2(n1074), .ZN(n526) );
  NAND2_X4 U266 ( .A1(n1075), .A2(n1074), .ZN(n527) );
  XNOR2_X2 U267 ( .A(n537), .B(n450), .ZN(product[60]) );
  OAI21_X4 U268 ( .B1(n445), .B2(n529), .A(n530), .ZN(n528) );
  NAND2_X4 U269 ( .A1(n680), .A2(n531), .ZN(n529) );
  AOI21_X4 U270 ( .B1(n681), .B2(n531), .A(n534), .ZN(n530) );
  INV_X4 U271 ( .A(n532), .ZN(n531) );
  INV_X4 U272 ( .A(n533), .ZN(n532) );
  NOR2_X4 U273 ( .A1(n542), .A2(n535), .ZN(n533) );
  OAI21_X4 U274 ( .B1(n543), .B2(n535), .A(n536), .ZN(n534) );
  NAND2_X4 U275 ( .A1(n1013), .A2(n536), .ZN(n450) );
  INV_X32 U276 ( .A(n535), .ZN(n1013) );
  NOR2_X4 U277 ( .A1(n1077), .A2(n1076), .ZN(n535) );
  NAND2_X4 U278 ( .A1(n1077), .A2(n1076), .ZN(n536) );
  XNOR2_X2 U279 ( .A(n552), .B(n451), .ZN(product[59]) );
  OAI21_X4 U280 ( .B1(n445), .B2(n538), .A(n539), .ZN(n537) );
  NAND2_X4 U281 ( .A1(n680), .A2(n540), .ZN(n538) );
  AOI21_X4 U282 ( .B1(n681), .B2(n540), .A(n541), .ZN(n539) );
  INV_X4 U283 ( .A(n542), .ZN(n540) );
  INV_X4 U284 ( .A(n543), .ZN(n541) );
  NAND2_X4 U285 ( .A1(n651), .A2(n544), .ZN(n542) );
  AOI21_X4 U286 ( .B1(n544), .B2(n652), .A(n545), .ZN(n543) );
  NOR2_X4 U287 ( .A1(n616), .A2(n546), .ZN(n544) );
  OAI21_X4 U288 ( .B1(n617), .B2(n546), .A(n547), .ZN(n545) );
  NAND2_X4 U289 ( .A1(n557), .A2(n548), .ZN(n546) );
  AOI21_X4 U290 ( .B1(n558), .B2(n548), .A(n549), .ZN(n547) );
  INV_X4 U291 ( .A(n550), .ZN(n548) );
  INV_X4 U292 ( .A(n551), .ZN(n549) );
  NAND2_X4 U293 ( .A1(n1014), .A2(n551), .ZN(n451) );
  INV_X32 U294 ( .A(n550), .ZN(n1014) );
  NOR2_X4 U295 ( .A1(n1078), .A2(n1081), .ZN(n550) );
  NAND2_X4 U296 ( .A1(n1078), .A2(n1081), .ZN(n551) );
  XNOR2_X2 U297 ( .A(n565), .B(n452), .ZN(product[58]) );
  OAI21_X4 U298 ( .B1(n445), .B2(n553), .A(n554), .ZN(n552) );
  NAND2_X4 U299 ( .A1(n608), .A2(n555), .ZN(n553) );
  AOI21_X4 U300 ( .B1(n609), .B2(n555), .A(n558), .ZN(n554) );
  INV_X4 U301 ( .A(n556), .ZN(n555) );
  INV_X4 U302 ( .A(n557), .ZN(n556) );
  NOR2_X4 U303 ( .A1(n590), .A2(n559), .ZN(n557) );
  OAI21_X4 U304 ( .B1(n591), .B2(n559), .A(n560), .ZN(n558) );
  NAND2_X4 U305 ( .A1(n570), .A2(n561), .ZN(n559) );
  AOI21_X4 U306 ( .B1(n571), .B2(n561), .A(n562), .ZN(n560) );
  INV_X4 U307 ( .A(n563), .ZN(n561) );
  INV_X4 U308 ( .A(n564), .ZN(n562) );
  NAND2_X4 U309 ( .A1(n1015), .A2(n564), .ZN(n452) );
  INV_X32 U316 ( .A(n563), .ZN(n1015) );
  NOR2_X4 U317 ( .A1(n1085), .A2(n1082), .ZN(n563) );
  NAND2_X4 U318 ( .A1(n1085), .A2(n1082), .ZN(n564) );
  XNOR2_X2 U319 ( .A(n574), .B(n453), .ZN(product[57]) );
  OAI21_X4 U320 ( .B1(n445), .B2(n566), .A(n567), .ZN(n565) );
  NAND2_X4 U321 ( .A1(n584), .A2(n568), .ZN(n566) );
  AOI21_X4 U322 ( .B1(n585), .B2(n568), .A(n571), .ZN(n567) );
  INV_X4 U323 ( .A(n569), .ZN(n568) );
  INV_X4 U324 ( .A(n570), .ZN(n569) );
  NOR2_X4 U325 ( .A1(n579), .A2(n572), .ZN(n570) );
  OAI21_X4 U326 ( .B1(n580), .B2(n572), .A(n573), .ZN(n571) );
  NAND2_X4 U327 ( .A1(n1016), .A2(n573), .ZN(n453) );
  INV_X32 U328 ( .A(n572), .ZN(n1016) );
  NOR2_X4 U329 ( .A1(n1086), .A2(n1091), .ZN(n572) );
  NAND2_X4 U330 ( .A1(n1086), .A2(n1091), .ZN(n573) );
  XNOR2_X2 U331 ( .A(n581), .B(n454), .ZN(product[56]) );
  OAI21_X4 U332 ( .B1(n445), .B2(n575), .A(n576), .ZN(n574) );
  NAND2_X4 U333 ( .A1(n584), .A2(n577), .ZN(n575) );
  AOI21_X4 U334 ( .B1(n585), .B2(n577), .A(n578), .ZN(n576) );
  INV_X4 U335 ( .A(n579), .ZN(n577) );
  INV_X4 U336 ( .A(n580), .ZN(n578) );
  NAND2_X4 U337 ( .A1(n1017), .A2(n580), .ZN(n454) );
  INV_X32 U338 ( .A(n579), .ZN(n1017) );
  NOR2_X4 U339 ( .A1(n1092), .A2(n1097), .ZN(n579) );
  NAND2_X4 U340 ( .A1(n1092), .A2(n1097), .ZN(n580) );
  XNOR2_X2 U341 ( .A(n596), .B(n455), .ZN(product[55]) );
  OAI21_X4 U342 ( .B1(n445), .B2(n582), .A(n583), .ZN(n581) );
  INV_X4 U343 ( .A(n584), .ZN(n582) );
  INV_X4 U344 ( .A(n585), .ZN(n583) );
  NOR2_X4 U345 ( .A1(n447), .A2(n586), .ZN(n584) );
  OAI21_X4 U346 ( .B1(n446), .B2(n586), .A(n587), .ZN(n585) );
  NAND2_X4 U347 ( .A1(n612), .A2(n588), .ZN(n586) );
  AOI21_X4 U348 ( .B1(n613), .B2(n588), .A(n589), .ZN(n587) );
  INV_X4 U349 ( .A(n590), .ZN(n588) );
  INV_X4 U350 ( .A(n591), .ZN(n589) );
  NAND2_X4 U351 ( .A1(n601), .A2(n592), .ZN(n590) );
  AOI21_X4 U352 ( .B1(n602), .B2(n592), .A(n593), .ZN(n591) );
  INV_X4 U353 ( .A(n594), .ZN(n592) );
  INV_X4 U354 ( .A(n595), .ZN(n593) );
  NAND2_X4 U355 ( .A1(n1018), .A2(n595), .ZN(n455) );
  INV_X32 U356 ( .A(n594), .ZN(n1018) );
  NOR2_X4 U357 ( .A1(n1098), .A2(n1105), .ZN(n594) );
  NAND2_X4 U358 ( .A1(n1098), .A2(n1105), .ZN(n595) );
  XNOR2_X2 U359 ( .A(n605), .B(n456), .ZN(product[54]) );
  OAI21_X4 U360 ( .B1(n445), .B2(n597), .A(n598), .ZN(n596) );
  NAND2_X4 U361 ( .A1(n608), .A2(n599), .ZN(n597) );
  AOI21_X4 U362 ( .B1(n609), .B2(n599), .A(n602), .ZN(n598) );
  INV_X4 U363 ( .A(n600), .ZN(n599) );
  INV_X4 U364 ( .A(n601), .ZN(n600) );
  INV_X4 U365 ( .A(n603), .ZN(n601) );
  INV_X4 U366 ( .A(n604), .ZN(n602) );
  NAND2_X4 U367 ( .A1(n1019), .A2(n604), .ZN(n456) );
  INV_X32 U368 ( .A(n603), .ZN(n1019) );
  NOR2_X4 U369 ( .A1(n1106), .A2(n1113), .ZN(n603) );
  NAND2_X4 U370 ( .A1(n1106), .A2(n1113), .ZN(n604) );
  XNOR2_X2 U371 ( .A(n622), .B(n457), .ZN(product[53]) );
  OAI21_X4 U372 ( .B1(n445), .B2(n606), .A(n607), .ZN(n605) );
  INV_X4 U373 ( .A(n608), .ZN(n606) );
  INV_X4 U374 ( .A(n609), .ZN(n607) );
  NOR2_X4 U375 ( .A1(n447), .A2(n610), .ZN(n608) );
  OAI21_X4 U376 ( .B1(n446), .B2(n610), .A(n611), .ZN(n609) );
  INV_X4 U377 ( .A(n612), .ZN(n610) );
  INV_X4 U378 ( .A(n613), .ZN(n611) );
  NOR2_X4 U379 ( .A1(n649), .A2(n614), .ZN(n612) );
  OAI21_X4 U380 ( .B1(n650), .B2(n614), .A(n617), .ZN(n613) );
  INV_X4 U381 ( .A(n615), .ZN(n614) );
  INV_X4 U382 ( .A(n616), .ZN(n615) );
  NAND2_X4 U383 ( .A1(n618), .A2(n638), .ZN(n616) );
  AOI21_X4 U384 ( .B1(n618), .B2(n639), .A(n619), .ZN(n617) );
  NOR2_X4 U385 ( .A1(n627), .A2(n620), .ZN(n618) );
  OAI21_X4 U386 ( .B1(n628), .B2(n620), .A(n621), .ZN(n619) );
  NAND2_X4 U387 ( .A1(n1020), .A2(n621), .ZN(n457) );
  INV_X32 U388 ( .A(n620), .ZN(n1020) );
  NOR2_X4 U389 ( .A1(n1114), .A2(n1123), .ZN(n620) );
  NAND2_X4 U390 ( .A1(n1114), .A2(n1123), .ZN(n621) );
  XNOR2_X2 U391 ( .A(n629), .B(n458), .ZN(product[52]) );
  OAI21_X4 U392 ( .B1(n445), .B2(n623), .A(n624), .ZN(n622) );
  NAND2_X4 U393 ( .A1(n632), .A2(n625), .ZN(n623) );
  AOI21_X4 U394 ( .B1(n633), .B2(n625), .A(n626), .ZN(n624) );
  INV_X4 U395 ( .A(n627), .ZN(n625) );
  INV_X4 U396 ( .A(n628), .ZN(n626) );
  NAND2_X4 U397 ( .A1(n1021), .A2(n628), .ZN(n458) );
  INV_X32 U398 ( .A(n627), .ZN(n1021) );
  NOR2_X4 U399 ( .A1(n1124), .A2(n1133), .ZN(n627) );
  NAND2_X4 U400 ( .A1(n1124), .A2(n1133), .ZN(n628) );
  XNOR2_X2 U401 ( .A(n642), .B(n459), .ZN(product[51]) );
  OAI21_X4 U402 ( .B1(n445), .B2(n630), .A(n631), .ZN(n629) );
  INV_X4 U403 ( .A(n632), .ZN(n630) );
  INV_X4 U404 ( .A(n633), .ZN(n631) );
  NOR2_X4 U405 ( .A1(n447), .A2(n634), .ZN(n632) );
  OAI21_X4 U406 ( .B1(n446), .B2(n634), .A(n635), .ZN(n633) );
  NAND2_X4 U407 ( .A1(n647), .A2(n636), .ZN(n634) );
  AOI21_X4 U408 ( .B1(n648), .B2(n636), .A(n639), .ZN(n635) );
  INV_X4 U409 ( .A(n637), .ZN(n636) );
  INV_X4 U410 ( .A(n638), .ZN(n637) );
  INV_X4 U411 ( .A(n640), .ZN(n638) );
  INV_X4 U412 ( .A(n641), .ZN(n639) );
  NAND2_X4 U413 ( .A1(n1022), .A2(n641), .ZN(n459) );
  INV_X32 U414 ( .A(n640), .ZN(n1022) );
  NOR2_X4 U415 ( .A1(n1134), .A2(n1145), .ZN(n640) );
  NAND2_X4 U416 ( .A1(n1134), .A2(n1145), .ZN(n641) );
  XNOR2_X2 U417 ( .A(n659), .B(n460), .ZN(product[50]) );
  OAI21_X4 U418 ( .B1(n445), .B2(n643), .A(n644), .ZN(n642) );
  NAND2_X4 U419 ( .A1(n680), .A2(n645), .ZN(n643) );
  AOI21_X4 U420 ( .B1(n681), .B2(n645), .A(n648), .ZN(n644) );
  INV_X4 U421 ( .A(n646), .ZN(n645) );
  INV_X4 U422 ( .A(n647), .ZN(n646) );
  INV_X4 U423 ( .A(n649), .ZN(n647) );
  INV_X4 U424 ( .A(n650), .ZN(n648) );
  INV_X4 U425 ( .A(n651), .ZN(n649) );
  INV_X4 U426 ( .A(n652), .ZN(n650) );
  NOR2_X4 U427 ( .A1(n675), .A2(n653), .ZN(n651) );
  OAI21_X4 U428 ( .B1(n653), .B2(n676), .A(n654), .ZN(n652) );
  NAND2_X4 U429 ( .A1(n664), .A2(n655), .ZN(n653) );
  AOI21_X4 U430 ( .B1(n665), .B2(n655), .A(n656), .ZN(n654) );
  INV_X4 U431 ( .A(n657), .ZN(n655) );
  INV_X4 U432 ( .A(n658), .ZN(n656) );
  NAND2_X4 U433 ( .A1(n1023), .A2(n658), .ZN(n460) );
  INV_X32 U434 ( .A(n657), .ZN(n1023) );
  NOR2_X4 U435 ( .A1(n1157), .A2(n1146), .ZN(n657) );
  NAND2_X4 U436 ( .A1(n1157), .A2(n1146), .ZN(n658) );
  XNOR2_X2 U437 ( .A(n668), .B(n461), .ZN(product[49]) );
  OAI21_X4 U438 ( .B1(n444), .B2(n660), .A(n661), .ZN(n659) );
  NAND2_X4 U439 ( .A1(n671), .A2(n662), .ZN(n660) );
  AOI21_X4 U440 ( .B1(n672), .B2(n662), .A(n665), .ZN(n661) );
  INV_X4 U441 ( .A(n663), .ZN(n662) );
  INV_X4 U442 ( .A(n664), .ZN(n663) );
  INV_X4 U443 ( .A(n666), .ZN(n664) );
  INV_X4 U444 ( .A(n667), .ZN(n665) );
  NAND2_X4 U445 ( .A1(n1024), .A2(n667), .ZN(n461) );
  INV_X32 U446 ( .A(n666), .ZN(n1024) );
  NOR2_X4 U447 ( .A1(n1158), .A2(n1171), .ZN(n666) );
  NAND2_X4 U448 ( .A1(n1158), .A2(n1171), .ZN(n667) );
  XNOR2_X2 U449 ( .A(n677), .B(n462), .ZN(product[48]) );
  OAI21_X4 U450 ( .B1(n444), .B2(n669), .A(n670), .ZN(n668) );
  INV_X4 U451 ( .A(n671), .ZN(n669) );
  INV_X4 U452 ( .A(n672), .ZN(n670) );
  NOR2_X4 U453 ( .A1(n447), .A2(n673), .ZN(n671) );
  OAI21_X4 U454 ( .B1(n446), .B2(n673), .A(n676), .ZN(n672) );
  INV_X4 U455 ( .A(n674), .ZN(n673) );
  INV_X4 U456 ( .A(n675), .ZN(n674) );
  NAND2_X4 U457 ( .A1(n1025), .A2(n676), .ZN(n462) );
  INV_X32 U458 ( .A(n675), .ZN(n1025) );
  NOR2_X4 U459 ( .A1(n1172), .A2(n1185), .ZN(n675) );
  NAND2_X4 U460 ( .A1(n1172), .A2(n1185), .ZN(n676) );
  XNOR2_X2 U461 ( .A(n692), .B(n463), .ZN(product[47]) );
  OAI21_X4 U462 ( .B1(n444), .B2(n678), .A(n679), .ZN(n677) );
  INV_X4 U463 ( .A(n680), .ZN(n678) );
  INV_X4 U464 ( .A(n681), .ZN(n679) );
  INV_X4 U465 ( .A(n447), .ZN(n680) );
  INV_X4 U466 ( .A(n446), .ZN(n681) );
  NAND2_X4 U467 ( .A1(n741), .A2(n684), .ZN(n682) );
  AOI21_X4 U468 ( .B1(n684), .B2(n742), .A(n685), .ZN(n683) );
  NOR2_X4 U469 ( .A1(n686), .A2(n719), .ZN(n684) );
  OAI21_X4 U470 ( .B1(n686), .B2(n720), .A(n687), .ZN(n685) );
  NAND2_X4 U471 ( .A1(n688), .A2(n708), .ZN(n686) );
  AOI21_X4 U472 ( .B1(n688), .B2(n709), .A(n689), .ZN(n687) );
  NOR2_X4 U473 ( .A1(n697), .A2(n690), .ZN(n688) );
  OAI21_X4 U474 ( .B1(n690), .B2(n698), .A(n691), .ZN(n689) );
  NAND2_X4 U475 ( .A1(n1026), .A2(n691), .ZN(n463) );
  INV_X32 U476 ( .A(n690), .ZN(n1026) );
  NOR2_X4 U477 ( .A1(n1186), .A2(n1201), .ZN(n690) );
  NAND2_X4 U478 ( .A1(n1186), .A2(n1201), .ZN(n691) );
  XNOR2_X2 U479 ( .A(n699), .B(n464), .ZN(product[46]) );
  OAI21_X4 U480 ( .B1(n444), .B2(n693), .A(n694), .ZN(n692) );
  NAND2_X4 U481 ( .A1(n702), .A2(n695), .ZN(n693) );
  AOI21_X4 U482 ( .B1(n703), .B2(n695), .A(n696), .ZN(n694) );
  INV_X4 U483 ( .A(n697), .ZN(n695) );
  INV_X4 U484 ( .A(n698), .ZN(n696) );
  NAND2_X4 U485 ( .A1(n1027), .A2(n698), .ZN(n464) );
  INV_X32 U486 ( .A(n697), .ZN(n1027) );
  NOR2_X4 U487 ( .A1(n1202), .A2(n1217), .ZN(n697) );
  NAND2_X4 U488 ( .A1(n1202), .A2(n1217), .ZN(n698) );
  XNOR2_X2 U489 ( .A(n712), .B(n465), .ZN(product[45]) );
  OAI21_X4 U490 ( .B1(n444), .B2(n700), .A(n701), .ZN(n699) );
  INV_X4 U491 ( .A(n702), .ZN(n700) );
  INV_X4 U492 ( .A(n703), .ZN(n701) );
  NOR2_X4 U493 ( .A1(n739), .A2(n704), .ZN(n702) );
  OAI21_X4 U494 ( .B1(n740), .B2(n704), .A(n705), .ZN(n703) );
  NAND2_X4 U495 ( .A1(n717), .A2(n706), .ZN(n704) );
  AOI21_X4 U496 ( .B1(n718), .B2(n706), .A(n709), .ZN(n705) );
  INV_X4 U497 ( .A(n707), .ZN(n706) );
  INV_X4 U498 ( .A(n708), .ZN(n707) );
  INV_X4 U499 ( .A(n710), .ZN(n708) );
  INV_X4 U500 ( .A(n711), .ZN(n709) );
  NAND2_X4 U501 ( .A1(n1028), .A2(n711), .ZN(n465) );
  INV_X32 U502 ( .A(n710), .ZN(n1028) );
  NOR2_X4 U503 ( .A1(n1218), .A2(n1235), .ZN(n710) );
  NAND2_X4 U504 ( .A1(n1218), .A2(n1235), .ZN(n711) );
  XNOR2_X2 U505 ( .A(n725), .B(n466), .ZN(product[44]) );
  OAI21_X4 U506 ( .B1(n444), .B2(n713), .A(n714), .ZN(n712) );
  NAND2_X4 U507 ( .A1(n737), .A2(n715), .ZN(n713) );
  AOI21_X4 U508 ( .B1(n738), .B2(n715), .A(n718), .ZN(n714) );
  INV_X4 U509 ( .A(n716), .ZN(n715) );
  INV_X4 U510 ( .A(n717), .ZN(n716) );
  INV_X4 U511 ( .A(n719), .ZN(n717) );
  INV_X4 U512 ( .A(n720), .ZN(n718) );
  NAND2_X4 U513 ( .A1(n730), .A2(n721), .ZN(n719) );
  AOI21_X4 U514 ( .B1(n721), .B2(n731), .A(n722), .ZN(n720) );
  INV_X4 U515 ( .A(n723), .ZN(n721) );
  INV_X4 U516 ( .A(n724), .ZN(n722) );
  NAND2_X4 U517 ( .A1(n1029), .A2(n724), .ZN(n466) );
  INV_X32 U518 ( .A(n723), .ZN(n1029) );
  NOR2_X4 U519 ( .A1(n1236), .A2(n1253), .ZN(n723) );
  NAND2_X4 U520 ( .A1(n1236), .A2(n1253), .ZN(n724) );
  XNOR2_X2 U521 ( .A(n734), .B(n467), .ZN(product[43]) );
  OAI21_X4 U522 ( .B1(n444), .B2(n726), .A(n727), .ZN(n725) );
  NAND2_X4 U523 ( .A1(n737), .A2(n728), .ZN(n726) );
  AOI21_X4 U524 ( .B1(n738), .B2(n728), .A(n731), .ZN(n727) );
  INV_X4 U525 ( .A(n729), .ZN(n728) );
  INV_X4 U526 ( .A(n730), .ZN(n729) );
  INV_X4 U527 ( .A(n732), .ZN(n730) );
  INV_X4 U528 ( .A(n733), .ZN(n731) );
  NAND2_X4 U529 ( .A1(n1030), .A2(n733), .ZN(n467) );
  INV_X32 U530 ( .A(n732), .ZN(n1030) );
  NOR2_X4 U531 ( .A1(n1254), .A2(n1273), .ZN(n732) );
  NAND2_X4 U532 ( .A1(n1254), .A2(n1273), .ZN(n733) );
  XNOR2_X2 U533 ( .A(n749), .B(n468), .ZN(product[42]) );
  OAI21_X4 U534 ( .B1(n444), .B2(n735), .A(n736), .ZN(n734) );
  INV_X4 U535 ( .A(n737), .ZN(n735) );
  INV_X4 U536 ( .A(n738), .ZN(n736) );
  INV_X4 U537 ( .A(n739), .ZN(n737) );
  INV_X4 U538 ( .A(n740), .ZN(n738) );
  INV_X4 U539 ( .A(n741), .ZN(n739) );
  INV_X4 U540 ( .A(n742), .ZN(n740) );
  NOR2_X4 U541 ( .A1(n763), .A2(n743), .ZN(n741) );
  OAI21_X4 U542 ( .B1(n743), .B2(n764), .A(n744), .ZN(n742) );
  NAND2_X4 U543 ( .A1(n754), .A2(n745), .ZN(n743) );
  AOI21_X4 U544 ( .B1(n745), .B2(n755), .A(n746), .ZN(n744) );
  INV_X4 U545 ( .A(n747), .ZN(n745) );
  INV_X4 U546 ( .A(n748), .ZN(n746) );
  NAND2_X4 U547 ( .A1(n1031), .A2(n748), .ZN(n468) );
  INV_X32 U548 ( .A(n747), .ZN(n1031) );
  NOR2_X4 U549 ( .A1(n1274), .A2(n1293), .ZN(n747) );
  NAND2_X4 U550 ( .A1(n1274), .A2(n1293), .ZN(n748) );
  XNOR2_X2 U551 ( .A(n758), .B(n469), .ZN(product[41]) );
  OAI21_X4 U552 ( .B1(n444), .B2(n750), .A(n751), .ZN(n749) );
  NAND2_X4 U553 ( .A1(n761), .A2(n752), .ZN(n750) );
  AOI21_X4 U554 ( .B1(n762), .B2(n752), .A(n755), .ZN(n751) );
  INV_X4 U555 ( .A(n753), .ZN(n752) );
  INV_X4 U556 ( .A(n754), .ZN(n753) );
  INV_X4 U557 ( .A(n756), .ZN(n754) );
  INV_X4 U558 ( .A(n757), .ZN(n755) );
  NAND2_X4 U559 ( .A1(n1032), .A2(n757), .ZN(n469) );
  INV_X32 U560 ( .A(n756), .ZN(n1032) );
  NOR2_X4 U561 ( .A1(n1294), .A2(n1315), .ZN(n756) );
  NAND2_X4 U562 ( .A1(n1294), .A2(n1315), .ZN(n757) );
  XOR2_X2 U563 ( .A(n444), .B(n470), .Z(product[40]) );
  OAI21_X4 U564 ( .B1(n444), .B2(n759), .A(n760), .ZN(n758) );
  INV_X4 U565 ( .A(n761), .ZN(n759) );
  INV_X4 U566 ( .A(n762), .ZN(n760) );
  INV_X4 U567 ( .A(n763), .ZN(n761) );
  INV_X4 U568 ( .A(n764), .ZN(n762) );
  NAND2_X4 U569 ( .A1(n1033), .A2(n764), .ZN(n470) );
  INV_X32 U570 ( .A(n763), .ZN(n1033) );
  NOR2_X4 U571 ( .A1(n1316), .A2(n1337), .ZN(n763) );
  NAND2_X4 U572 ( .A1(n1316), .A2(n1337), .ZN(n764) );
  XNOR2_X2 U573 ( .A(n774), .B(n471), .ZN(product[39]) );
  AOI21_X4 U574 ( .B1(n766), .B2(n834), .A(n767), .ZN(n765) );
  NOR2_X4 U575 ( .A1(n806), .A2(n768), .ZN(n766) );
  OAI21_X4 U576 ( .B1(n807), .B2(n768), .A(n769), .ZN(n767) );
  NAND2_X4 U577 ( .A1(n790), .A2(n770), .ZN(n768) );
  AOI21_X4 U578 ( .B1(n770), .B2(n791), .A(n771), .ZN(n769) );
  NOR2_X4 U579 ( .A1(n781), .A2(n772), .ZN(n770) );
  OAI21_X4 U580 ( .B1(n782), .B2(n772), .A(n773), .ZN(n771) );
  NAND2_X4 U581 ( .A1(n1034), .A2(n773), .ZN(n471) );
  INV_X32 U582 ( .A(n772), .ZN(n1034) );
  NOR2_X4 U583 ( .A1(n1338), .A2(n1361), .ZN(n772) );
  NAND2_X4 U584 ( .A1(n1338), .A2(n1361), .ZN(n773) );
  XNOR2_X2 U585 ( .A(n783), .B(n472), .ZN(product[38]) );
  OAI21_X4 U586 ( .B1(n775), .B2(n833), .A(n776), .ZN(n774) );
  NAND2_X4 U587 ( .A1(n777), .A2(n804), .ZN(n775) );
  AOI21_X4 U588 ( .B1(n805), .B2(n777), .A(n778), .ZN(n776) );
  NOR2_X4 U589 ( .A1(n788), .A2(n779), .ZN(n777) );
  OAI21_X4 U590 ( .B1(n789), .B2(n779), .A(n782), .ZN(n778) );
  INV_X4 U591 ( .A(n780), .ZN(n779) );
  INV_X4 U592 ( .A(n781), .ZN(n780) );
  NAND2_X4 U593 ( .A1(n1035), .A2(n782), .ZN(n472) );
  INV_X32 U594 ( .A(n781), .ZN(n1035) );
  NOR2_X4 U595 ( .A1(n1362), .A2(n1385), .ZN(n781) );
  NAND2_X4 U596 ( .A1(n1362), .A2(n1385), .ZN(n782) );
  XNOR2_X2 U597 ( .A(n794), .B(n473), .ZN(product[37]) );
  OAI21_X4 U598 ( .B1(n833), .B2(n784), .A(n785), .ZN(n783) );
  NAND2_X4 U599 ( .A1(n804), .A2(n786), .ZN(n784) );
  AOI21_X4 U600 ( .B1(n805), .B2(n786), .A(n787), .ZN(n785) );
  INV_X4 U601 ( .A(n788), .ZN(n786) );
  INV_X4 U602 ( .A(n789), .ZN(n787) );
  INV_X4 U603 ( .A(n790), .ZN(n788) );
  INV_X4 U604 ( .A(n791), .ZN(n789) );
  NOR2_X4 U605 ( .A1(n799), .A2(n792), .ZN(n790) );
  OAI21_X4 U606 ( .B1(n792), .B2(n800), .A(n793), .ZN(n791) );
  NAND2_X4 U607 ( .A1(n1036), .A2(n793), .ZN(n473) );
  INV_X32 U608 ( .A(n792), .ZN(n1036) );
  NOR2_X4 U609 ( .A1(n1386), .A2(n1411), .ZN(n792) );
  NAND2_X4 U610 ( .A1(n1386), .A2(n1411), .ZN(n793) );
  XNOR2_X2 U611 ( .A(n801), .B(n474), .ZN(product[36]) );
  OAI21_X4 U612 ( .B1(n833), .B2(n795), .A(n796), .ZN(n794) );
  NAND2_X4 U613 ( .A1(n804), .A2(n797), .ZN(n795) );
  AOI21_X4 U614 ( .B1(n805), .B2(n797), .A(n798), .ZN(n796) );
  INV_X4 U615 ( .A(n799), .ZN(n797) );
  INV_X4 U616 ( .A(n800), .ZN(n798) );
  NAND2_X4 U617 ( .A1(n1037), .A2(n800), .ZN(n474) );
  INV_X32 U618 ( .A(n799), .ZN(n1037) );
  NOR2_X4 U619 ( .A1(n1412), .A2(n1437), .ZN(n799) );
  NAND2_X4 U620 ( .A1(n1412), .A2(n1437), .ZN(n800) );
  XNOR2_X2 U621 ( .A(n812), .B(n475), .ZN(product[35]) );
  OAI21_X4 U622 ( .B1(n833), .B2(n802), .A(n803), .ZN(n801) );
  INV_X4 U623 ( .A(n804), .ZN(n802) );
  INV_X4 U624 ( .A(n805), .ZN(n803) );
  INV_X4 U625 ( .A(n806), .ZN(n804) );
  INV_X4 U626 ( .A(n807), .ZN(n805) );
  NAND2_X4 U627 ( .A1(n826), .A2(n808), .ZN(n806) );
  AOI21_X4 U628 ( .B1(n808), .B2(n827), .A(n809), .ZN(n807) );
  NOR2_X4 U629 ( .A1(n810), .A2(n817), .ZN(n808) );
  OAI21_X4 U630 ( .B1(n810), .B2(n818), .A(n811), .ZN(n809) );
  NAND2_X4 U631 ( .A1(n1038), .A2(n811), .ZN(n475) );
  INV_X32 U632 ( .A(n810), .ZN(n1038) );
  NOR2_X4 U633 ( .A1(n1438), .A2(n1465), .ZN(n810) );
  NAND2_X4 U634 ( .A1(n1438), .A2(n1465), .ZN(n811) );
  XNOR2_X2 U635 ( .A(n819), .B(n476), .ZN(product[34]) );
  OAI21_X4 U636 ( .B1(n833), .B2(n813), .A(n814), .ZN(n812) );
  NAND2_X4 U637 ( .A1(n822), .A2(n815), .ZN(n813) );
  AOI21_X4 U638 ( .B1(n823), .B2(n815), .A(n816), .ZN(n814) );
  INV_X4 U639 ( .A(n817), .ZN(n815) );
  INV_X4 U640 ( .A(n818), .ZN(n816) );
  NAND2_X4 U641 ( .A1(n1039), .A2(n818), .ZN(n476) );
  INV_X32 U642 ( .A(n817), .ZN(n1039) );
  NOR2_X4 U643 ( .A1(n1466), .A2(n1493), .ZN(n817) );
  NAND2_X4 U644 ( .A1(n1466), .A2(n1493), .ZN(n818) );
  XNOR2_X2 U645 ( .A(n830), .B(n477), .ZN(product[33]) );
  OAI21_X4 U646 ( .B1(n833), .B2(n820), .A(n821), .ZN(n819) );
  INV_X4 U647 ( .A(n822), .ZN(n820) );
  INV_X4 U648 ( .A(n823), .ZN(n821) );
  INV_X4 U649 ( .A(n824), .ZN(n822) );
  INV_X4 U650 ( .A(n825), .ZN(n823) );
  INV_X4 U651 ( .A(n826), .ZN(n824) );
  INV_X4 U652 ( .A(n827), .ZN(n825) );
  NOR2_X4 U653 ( .A1(n831), .A2(n828), .ZN(n826) );
  OAI21_X4 U654 ( .B1(n828), .B2(n832), .A(n829), .ZN(n827) );
  NAND2_X4 U655 ( .A1(n1040), .A2(n829), .ZN(n477) );
  INV_X32 U656 ( .A(n828), .ZN(n1040) );
  NOR2_X4 U657 ( .A1(n1494), .A2(n1523), .ZN(n828) );
  NAND2_X4 U658 ( .A1(n1494), .A2(n1523), .ZN(n829) );
  XOR2_X2 U659 ( .A(n833), .B(n478), .Z(product[32]) );
  OAI21_X4 U660 ( .B1(n833), .B2(n831), .A(n832), .ZN(n830) );
  NAND2_X4 U661 ( .A1(n1041), .A2(n832), .ZN(n478) );
  INV_X32 U662 ( .A(n831), .ZN(n1041) );
  NOR2_X4 U663 ( .A1(n1524), .A2(n1553), .ZN(n831) );
  NAND2_X4 U664 ( .A1(n1524), .A2(n1553), .ZN(n832) );
  XNOR2_X2 U665 ( .A(n841), .B(n479), .ZN(product[31]) );
  INV_X4 U666 ( .A(n834), .ZN(n833) );
  OAI21_X4 U667 ( .B1(n835), .B2(n855), .A(n836), .ZN(n834) );
  NAND2_X4 U668 ( .A1(n837), .A2(n845), .ZN(n835) );
  AOI21_X4 U669 ( .B1(n837), .B2(n846), .A(n838), .ZN(n836) );
  NOR2_X4 U670 ( .A1(n842), .A2(n839), .ZN(n837) );
  OAI21_X4 U671 ( .B1(n839), .B2(n843), .A(n840), .ZN(n838) );
  NAND2_X4 U672 ( .A1(n1042), .A2(n840), .ZN(n479) );
  INV_X32 U673 ( .A(n839), .ZN(n1042) );
  NOR2_X4 U674 ( .A1(n1554), .A2(n1583), .ZN(n839) );
  NAND2_X4 U675 ( .A1(n1554), .A2(n1583), .ZN(n840) );
  XOR2_X2 U676 ( .A(n844), .B(n480), .Z(product[30]) );
  OAI21_X4 U677 ( .B1(n844), .B2(n842), .A(n843), .ZN(n841) );
  NAND2_X4 U678 ( .A1(n1043), .A2(n843), .ZN(n480) );
  INV_X32 U679 ( .A(n842), .ZN(n1043) );
  NOR2_X4 U680 ( .A1(n1584), .A2(n1611), .ZN(n842) );
  NAND2_X4 U681 ( .A1(n1584), .A2(n1611), .ZN(n843) );
  XOR2_X2 U682 ( .A(n849), .B(n481), .Z(product[29]) );
  AOI21_X4 U683 ( .B1(n854), .B2(n845), .A(n846), .ZN(n844) );
  NOR2_X4 U684 ( .A1(n847), .A2(n852), .ZN(n845) );
  OAI21_X4 U685 ( .B1(n847), .B2(n853), .A(n848), .ZN(n846) );
  NAND2_X4 U686 ( .A1(n1044), .A2(n848), .ZN(n481) );
  INV_X32 U687 ( .A(n847), .ZN(n1044) );
  NOR2_X4 U688 ( .A1(n1612), .A2(n1639), .ZN(n847) );
  NAND2_X4 U689 ( .A1(n1612), .A2(n1639), .ZN(n848) );
  XNOR2_X2 U690 ( .A(n854), .B(n482), .ZN(product[28]) );
  AOI21_X4 U691 ( .B1(n854), .B2(n850), .A(n851), .ZN(n849) );
  INV_X4 U692 ( .A(n852), .ZN(n850) );
  INV_X4 U693 ( .A(n853), .ZN(n851) );
  NAND2_X4 U694 ( .A1(n1045), .A2(n853), .ZN(n482) );
  INV_X32 U695 ( .A(n852), .ZN(n1045) );
  NOR2_X4 U696 ( .A1(n1640), .A2(n1665), .ZN(n852) );
  NAND2_X4 U697 ( .A1(n1640), .A2(n1665), .ZN(n853) );
  XOR2_X2 U698 ( .A(n864), .B(n483), .Z(product[27]) );
  INV_X4 U699 ( .A(n855), .ZN(n854) );
  AOI21_X4 U700 ( .B1(n884), .B2(n856), .A(n857), .ZN(n855) );
  NOR2_X4 U701 ( .A1(n858), .A2(n870), .ZN(n856) );
  OAI21_X4 U702 ( .B1(n871), .B2(n858), .A(n859), .ZN(n857) );
  NAND2_X4 U703 ( .A1(n860), .A2(n865), .ZN(n858) );
  AOI21_X4 U704 ( .B1(n860), .B2(n866), .A(n861), .ZN(n859) );
  INV_X4 U705 ( .A(n862), .ZN(n860) );
  INV_X4 U706 ( .A(n863), .ZN(n861) );
  NAND2_X4 U707 ( .A1(n1046), .A2(n863), .ZN(n483) );
  INV_X32 U708 ( .A(n862), .ZN(n1046) );
  NOR2_X4 U709 ( .A1(n1666), .A2(n1691), .ZN(n862) );
  NAND2_X4 U710 ( .A1(n1666), .A2(n1691), .ZN(n863) );
  XNOR2_X2 U711 ( .A(n869), .B(n484), .ZN(product[26]) );
  AOI21_X4 U712 ( .B1(n869), .B2(n865), .A(n866), .ZN(n864) );
  INV_X4 U713 ( .A(n867), .ZN(n865) );
  INV_X4 U714 ( .A(n868), .ZN(n866) );
  NAND2_X4 U715 ( .A1(n1047), .A2(n868), .ZN(n484) );
  INV_X32 U716 ( .A(n867), .ZN(n1047) );
  NOR2_X4 U717 ( .A1(n1692), .A2(n1715), .ZN(n867) );
  NAND2_X4 U718 ( .A1(n1692), .A2(n1715), .ZN(n868) );
  XNOR2_X2 U719 ( .A(n876), .B(n485), .ZN(product[25]) );
  OAI21_X4 U720 ( .B1(n883), .B2(n870), .A(n871), .ZN(n869) );
  NAND2_X4 U721 ( .A1(n872), .A2(n879), .ZN(n870) );
  AOI21_X4 U722 ( .B1(n872), .B2(n880), .A(n873), .ZN(n871) );
  INV_X4 U723 ( .A(n874), .ZN(n872) );
  INV_X4 U724 ( .A(n875), .ZN(n873) );
  NAND2_X4 U725 ( .A1(n1048), .A2(n875), .ZN(n485) );
  INV_X32 U726 ( .A(n874), .ZN(n1048) );
  NOR2_X4 U727 ( .A1(n1716), .A2(n1739), .ZN(n874) );
  NAND2_X4 U728 ( .A1(n1716), .A2(n1739), .ZN(n875) );
  XOR2_X2 U729 ( .A(n883), .B(n486), .Z(product[24]) );
  OAI21_X4 U730 ( .B1(n883), .B2(n877), .A(n878), .ZN(n876) );
  INV_X4 U731 ( .A(n879), .ZN(n877) );
  INV_X4 U732 ( .A(n880), .ZN(n878) );
  INV_X4 U733 ( .A(n881), .ZN(n879) );
  INV_X4 U734 ( .A(n882), .ZN(n880) );
  NAND2_X4 U735 ( .A1(n1049), .A2(n882), .ZN(n486) );
  INV_X32 U736 ( .A(n881), .ZN(n1049) );
  NOR2_X4 U737 ( .A1(n1740), .A2(n1761), .ZN(n881) );
  NAND2_X4 U738 ( .A1(n1740), .A2(n1761), .ZN(n882) );
  XNOR2_X2 U739 ( .A(n891), .B(n487), .ZN(product[23]) );
  INV_X4 U740 ( .A(n884), .ZN(n883) );
  OAI21_X4 U741 ( .B1(n885), .B2(n905), .A(n886), .ZN(n884) );
  NAND2_X4 U742 ( .A1(n887), .A2(n895), .ZN(n885) );
  AOI21_X4 U743 ( .B1(n887), .B2(n896), .A(n888), .ZN(n886) );
  NOR2_X4 U744 ( .A1(n889), .A2(n892), .ZN(n887) );
  OAI21_X4 U745 ( .B1(n889), .B2(n893), .A(n890), .ZN(n888) );
  NAND2_X4 U746 ( .A1(n1050), .A2(n890), .ZN(n487) );
  INV_X32 U747 ( .A(n889), .ZN(n1050) );
  NOR2_X4 U748 ( .A1(n1762), .A2(n1783), .ZN(n889) );
  NAND2_X4 U749 ( .A1(n1762), .A2(n1783), .ZN(n890) );
  XOR2_X2 U750 ( .A(n894), .B(n488), .Z(product[22]) );
  OAI21_X4 U751 ( .B1(n894), .B2(n892), .A(n893), .ZN(n891) );
  NAND2_X4 U752 ( .A1(n1051), .A2(n893), .ZN(n488) );
  INV_X32 U753 ( .A(n892), .ZN(n1051) );
  NOR2_X4 U754 ( .A1(n1784), .A2(n1803), .ZN(n892) );
  NAND2_X4 U755 ( .A1(n1784), .A2(n1803), .ZN(n893) );
  XOR2_X2 U756 ( .A(n899), .B(n489), .Z(product[21]) );
  AOI21_X4 U757 ( .B1(n904), .B2(n895), .A(n896), .ZN(n894) );
  NOR2_X4 U758 ( .A1(n897), .A2(n902), .ZN(n895) );
  OAI21_X4 U759 ( .B1(n897), .B2(n903), .A(n898), .ZN(n896) );
  NAND2_X4 U760 ( .A1(n1052), .A2(n898), .ZN(n489) );
  INV_X32 U761 ( .A(n897), .ZN(n1052) );
  NOR2_X4 U762 ( .A1(n1804), .A2(n1823), .ZN(n897) );
  NAND2_X4 U763 ( .A1(n1804), .A2(n1823), .ZN(n898) );
  XNOR2_X2 U764 ( .A(n904), .B(n490), .ZN(product[20]) );
  AOI21_X4 U765 ( .B1(n904), .B2(n900), .A(n901), .ZN(n899) );
  INV_X4 U766 ( .A(n902), .ZN(n900) );
  INV_X4 U767 ( .A(n903), .ZN(n901) );
  NAND2_X4 U768 ( .A1(n1053), .A2(n903), .ZN(n490) );
  INV_X32 U769 ( .A(n902), .ZN(n1053) );
  NOR2_X4 U770 ( .A1(n1824), .A2(n1841), .ZN(n902) );
  NAND2_X4 U771 ( .A1(n1824), .A2(n1841), .ZN(n903) );
  XOR2_X2 U772 ( .A(n914), .B(n491), .Z(product[19]) );
  INV_X4 U773 ( .A(n905), .ZN(n904) );
  AOI21_X4 U774 ( .B1(n906), .B2(n934), .A(n907), .ZN(n905) );
  NOR2_X4 U775 ( .A1(n908), .A2(n920), .ZN(n906) );
  OAI21_X4 U776 ( .B1(n908), .B2(n921), .A(n909), .ZN(n907) );
  NAND2_X4 U777 ( .A1(n910), .A2(n915), .ZN(n908) );
  AOI21_X4 U778 ( .B1(n910), .B2(n916), .A(n911), .ZN(n909) );
  INV_X4 U779 ( .A(n912), .ZN(n910) );
  INV_X4 U780 ( .A(n913), .ZN(n911) );
  NAND2_X4 U781 ( .A1(n1054), .A2(n913), .ZN(n491) );
  INV_X32 U782 ( .A(n912), .ZN(n1054) );
  NOR2_X4 U783 ( .A1(n1842), .A2(n1859), .ZN(n912) );
  NAND2_X4 U784 ( .A1(n1842), .A2(n1859), .ZN(n913) );
  XNOR2_X2 U785 ( .A(n919), .B(n492), .ZN(product[18]) );
  AOI21_X4 U786 ( .B1(n919), .B2(n915), .A(n916), .ZN(n914) );
  INV_X4 U787 ( .A(n917), .ZN(n915) );
  INV_X4 U788 ( .A(n918), .ZN(n916) );
  NAND2_X4 U789 ( .A1(n1055), .A2(n918), .ZN(n492) );
  INV_X32 U790 ( .A(n917), .ZN(n1055) );
  NOR2_X4 U791 ( .A1(n1860), .A2(n1875), .ZN(n917) );
  NAND2_X4 U792 ( .A1(n1860), .A2(n1875), .ZN(n918) );
  XNOR2_X2 U793 ( .A(n926), .B(n493), .ZN(product[17]) );
  OAI21_X4 U794 ( .B1(n933), .B2(n920), .A(n921), .ZN(n919) );
  NAND2_X4 U795 ( .A1(n922), .A2(n929), .ZN(n920) );
  AOI21_X4 U796 ( .B1(n922), .B2(n930), .A(n923), .ZN(n921) );
  INV_X4 U797 ( .A(n924), .ZN(n922) );
  INV_X4 U798 ( .A(n925), .ZN(n923) );
  NAND2_X4 U799 ( .A1(n1056), .A2(n925), .ZN(n493) );
  INV_X32 U800 ( .A(n924), .ZN(n1056) );
  NOR2_X4 U801 ( .A1(n1876), .A2(n1891), .ZN(n924) );
  NAND2_X4 U802 ( .A1(n1876), .A2(n1891), .ZN(n925) );
  XOR2_X2 U803 ( .A(n933), .B(n494), .Z(product[16]) );
  OAI21_X4 U804 ( .B1(n933), .B2(n927), .A(n928), .ZN(n926) );
  INV_X4 U805 ( .A(n929), .ZN(n927) );
  INV_X4 U806 ( .A(n930), .ZN(n928) );
  INV_X4 U807 ( .A(n931), .ZN(n929) );
  INV_X4 U808 ( .A(n932), .ZN(n930) );
  NAND2_X4 U809 ( .A1(n1057), .A2(n932), .ZN(n494) );
  INV_X32 U810 ( .A(n931), .ZN(n1057) );
  NOR2_X4 U811 ( .A1(n1892), .A2(n1905), .ZN(n931) );
  NAND2_X4 U812 ( .A1(n1892), .A2(n1905), .ZN(n932) );
  XOR2_X2 U813 ( .A(n941), .B(n495), .Z(product[15]) );
  INV_X4 U814 ( .A(n934), .ZN(n933) );
  OAI21_X4 U815 ( .B1(n947), .B2(n935), .A(n936), .ZN(n934) );
  NAND2_X4 U816 ( .A1(n937), .A2(n942), .ZN(n935) );
  AOI21_X4 U817 ( .B1(n937), .B2(n943), .A(n938), .ZN(n936) );
  INV_X4 U818 ( .A(n939), .ZN(n937) );
  INV_X4 U819 ( .A(n940), .ZN(n938) );
  NAND2_X4 U820 ( .A1(n1058), .A2(n940), .ZN(n495) );
  INV_X32 U821 ( .A(n939), .ZN(n1058) );
  NOR2_X4 U822 ( .A1(n1906), .A2(n1919), .ZN(n939) );
  NAND2_X4 U823 ( .A1(n1906), .A2(n1919), .ZN(n940) );
  XNOR2_X2 U824 ( .A(n946), .B(n496), .ZN(product[14]) );
  AOI21_X4 U825 ( .B1(n946), .B2(n942), .A(n943), .ZN(n941) );
  INV_X4 U826 ( .A(n944), .ZN(n942) );
  INV_X4 U827 ( .A(n945), .ZN(n943) );
  NAND2_X4 U828 ( .A1(n1059), .A2(n945), .ZN(n496) );
  INV_X32 U829 ( .A(n944), .ZN(n1059) );
  NOR2_X4 U830 ( .A1(n1920), .A2(n1931), .ZN(n944) );
  NAND2_X4 U831 ( .A1(n1920), .A2(n1931), .ZN(n945) );
  XNOR2_X2 U832 ( .A(n952), .B(n497), .ZN(product[13]) );
  INV_X4 U833 ( .A(n947), .ZN(n946) );
  AOI21_X4 U834 ( .B1(n948), .B2(n956), .A(n949), .ZN(n947) );
  NOR2_X4 U835 ( .A1(n950), .A2(n953), .ZN(n948) );
  OAI21_X4 U836 ( .B1(n950), .B2(n954), .A(n951), .ZN(n949) );
  NAND2_X4 U837 ( .A1(n1060), .A2(n951), .ZN(n497) );
  INV_X32 U838 ( .A(n950), .ZN(n1060) );
  NOR2_X4 U839 ( .A1(n1932), .A2(n1943), .ZN(n950) );
  NAND2_X4 U840 ( .A1(n1932), .A2(n1943), .ZN(n951) );
  XOR2_X2 U841 ( .A(n955), .B(n498), .Z(product[12]) );
  OAI21_X4 U842 ( .B1(n955), .B2(n953), .A(n954), .ZN(n952) );
  NAND2_X4 U843 ( .A1(n1061), .A2(n954), .ZN(n498) );
  INV_X32 U844 ( .A(n953), .ZN(n1061) );
  NOR2_X4 U845 ( .A1(n1944), .A2(n1953), .ZN(n953) );
  NAND2_X4 U846 ( .A1(n1944), .A2(n1953), .ZN(n954) );
  XOR2_X2 U847 ( .A(n963), .B(n499), .Z(product[11]) );
  INV_X4 U848 ( .A(n956), .ZN(n955) );
  OAI21_X4 U849 ( .B1(n957), .B2(n969), .A(n958), .ZN(n956) );
  NAND2_X4 U850 ( .A1(n964), .A2(n959), .ZN(n957) );
  AOI21_X4 U851 ( .B1(n959), .B2(n965), .A(n960), .ZN(n958) );
  INV_X4 U852 ( .A(n961), .ZN(n959) );
  INV_X4 U853 ( .A(n962), .ZN(n960) );
  NAND2_X4 U854 ( .A1(n1062), .A2(n962), .ZN(n499) );
  INV_X32 U855 ( .A(n961), .ZN(n1062) );
  NOR2_X4 U856 ( .A1(n1954), .A2(n1963), .ZN(n961) );
  NAND2_X4 U857 ( .A1(n1954), .A2(n1963), .ZN(n962) );
  XNOR2_X2 U858 ( .A(n500), .B(n968), .ZN(product[10]) );
  AOI21_X4 U859 ( .B1(n968), .B2(n964), .A(n965), .ZN(n963) );
  INV_X4 U860 ( .A(n966), .ZN(n964) );
  INV_X4 U861 ( .A(n967), .ZN(n965) );
  NAND2_X4 U862 ( .A1(n1063), .A2(n967), .ZN(n500) );
  INV_X32 U863 ( .A(n966), .ZN(n1063) );
  NOR2_X4 U864 ( .A1(n1964), .A2(n1971), .ZN(n966) );
  NAND2_X4 U865 ( .A1(n1964), .A2(n1971), .ZN(n967) );
  XNOR2_X2 U866 ( .A(n501), .B(n974), .ZN(product[9]) );
  INV_X4 U867 ( .A(n969), .ZN(n968) );
  AOI21_X4 U868 ( .B1(n974), .B2(n970), .A(n971), .ZN(n969) );
  INV_X4 U869 ( .A(n972), .ZN(n970) );
  INV_X4 U870 ( .A(n973), .ZN(n971) );
  NAND2_X4 U871 ( .A1(n1064), .A2(n973), .ZN(n501) );
  INV_X32 U872 ( .A(n972), .ZN(n1064) );
  NOR2_X4 U873 ( .A1(n1972), .A2(n1979), .ZN(n972) );
  NAND2_X4 U874 ( .A1(n1972), .A2(n1979), .ZN(n973) );
  XOR2_X2 U875 ( .A(n981), .B(n502), .Z(product[8]) );
  OAI21_X4 U876 ( .B1(n975), .B2(n987), .A(n976), .ZN(n974) );
  NAND2_X4 U877 ( .A1(n977), .A2(n982), .ZN(n975) );
  AOI21_X4 U878 ( .B1(n977), .B2(n983), .A(n978), .ZN(n976) );
  INV_X4 U879 ( .A(n979), .ZN(n977) );
  INV_X4 U880 ( .A(n980), .ZN(n978) );
  NAND2_X4 U881 ( .A1(n1065), .A2(n980), .ZN(n502) );
  INV_X32 U882 ( .A(n979), .ZN(n1065) );
  NOR2_X4 U883 ( .A1(n1980), .A2(n1985), .ZN(n979) );
  NAND2_X4 U884 ( .A1(n1980), .A2(n1985), .ZN(n980) );
  XNOR2_X2 U885 ( .A(n986), .B(n503), .ZN(product[7]) );
  AOI21_X4 U886 ( .B1(n986), .B2(n982), .A(n983), .ZN(n981) );
  INV_X4 U887 ( .A(n984), .ZN(n982) );
  INV_X4 U888 ( .A(n985), .ZN(n983) );
  NAND2_X4 U889 ( .A1(n1066), .A2(n985), .ZN(n503) );
  INV_X32 U890 ( .A(n984), .ZN(n1066) );
  NOR2_X4 U891 ( .A1(n1986), .A2(n1991), .ZN(n984) );
  NAND2_X4 U892 ( .A1(n1986), .A2(n1991), .ZN(n985) );
  XNOR2_X2 U893 ( .A(n504), .B(n992), .ZN(product[6]) );
  INV_X4 U894 ( .A(n987), .ZN(n986) );
  AOI21_X4 U895 ( .B1(n988), .B2(n992), .A(n989), .ZN(n987) );
  INV_X4 U896 ( .A(n990), .ZN(n988) );
  INV_X4 U897 ( .A(n991), .ZN(n989) );
  NAND2_X4 U898 ( .A1(n1067), .A2(n991), .ZN(n504) );
  INV_X32 U899 ( .A(n990), .ZN(n1067) );
  NOR2_X4 U900 ( .A1(n1992), .A2(n1995), .ZN(n990) );
  NAND2_X4 U901 ( .A1(n1992), .A2(n1995), .ZN(n991) );
  XNOR2_X2 U902 ( .A(n505), .B(n998), .ZN(product[5]) );
  INV_X4 U903 ( .A(n993), .ZN(n992) );
  AOI21_X4 U904 ( .B1(n994), .B2(n998), .A(n995), .ZN(n993) );
  INV_X4 U905 ( .A(n996), .ZN(n994) );
  INV_X4 U906 ( .A(n997), .ZN(n995) );
  NAND2_X4 U907 ( .A1(n1068), .A2(n997), .ZN(n505) );
  INV_X32 U908 ( .A(n996), .ZN(n1068) );
  NOR2_X4 U909 ( .A1(n1996), .A2(n1999), .ZN(n996) );
  NAND2_X4 U910 ( .A1(n1996), .A2(n1999), .ZN(n997) );
  XOR2_X2 U911 ( .A(n506), .B(n1001), .Z(product[4]) );
  OAI21_X4 U912 ( .B1(n999), .B2(n1001), .A(n1000), .ZN(n998) );
  NAND2_X4 U913 ( .A1(n1069), .A2(n1000), .ZN(n506) );
  INV_X32 U914 ( .A(n999), .ZN(n1069) );
  NOR2_X4 U915 ( .A1(n2000), .A2(n2001), .ZN(n999) );
  NAND2_X4 U916 ( .A1(n2000), .A2(n2001), .ZN(n1000) );
  XNOR2_X2 U917 ( .A(n507), .B(n1006), .ZN(product[3]) );
  AOI21_X4 U918 ( .B1(n1002), .B2(n1006), .A(n1003), .ZN(n1001) );
  INV_X4 U919 ( .A(n1004), .ZN(n1002) );
  INV_X4 U920 ( .A(n1005), .ZN(n1003) );
  NAND2_X4 U921 ( .A1(n1070), .A2(n1005), .ZN(n507) );
  INV_X32 U922 ( .A(n1004), .ZN(n1070) );
  NOR2_X4 U923 ( .A1(n2002), .A2(n2017), .ZN(n1004) );
  NAND2_X4 U924 ( .A1(n2002), .A2(n2017), .ZN(n1005) );
  XOR2_X2 U925 ( .A(n508), .B(n1010), .Z(product[2]) );
  OAI21_X4 U926 ( .B1(n1007), .B2(n1010), .A(n1008), .ZN(n1006) );
  NAND2_X4 U927 ( .A1(n1071), .A2(n1008), .ZN(n508) );
  INV_X32 U928 ( .A(n1007), .ZN(n1071) );
  NOR2_X4 U929 ( .A1(n2498), .A2(n2529), .ZN(n1007) );
  NAND2_X4 U930 ( .A1(n2498), .A2(n2529), .ZN(n1008) );
  INV_X32 U931 ( .A(n509), .ZN(product[1]) );
  NAND2_X4 U932 ( .A1(n1072), .A2(n1010), .ZN(n509) );
  INV_X32 U933 ( .A(n1009), .ZN(n1072) );
  NOR2_X4 U934 ( .A1(n2530), .A2(n2018), .ZN(n1009) );
  NAND2_X4 U935 ( .A1(n2530), .A2(n2018), .ZN(n1010) );
  INV_X32 U936 ( .A(n1073), .ZN(n1074) );
  FA_X1 U937 ( .A(n2020), .B(n1079), .CI(n2051), .CO(n1075), .S(n1076) );
  FA_X1 U938 ( .A(n1080), .B(n2021), .CI(n1083), .CO(n1077), .S(n1078) );
  INV_X32 U939 ( .A(n1079), .ZN(n1080) );
  FA_X1 U940 ( .A(n1087), .B(n2083), .CI(n1084), .CO(n1081), .S(n1082) );
  FA_X1 U941 ( .A(n2052), .B(n1089), .CI(n2022), .CO(n1083), .S(n1084) );
  FA_X1 U942 ( .A(n1088), .B(n1095), .CI(n1093), .CO(n1085), .S(n1086) );
  FA_X1 U943 ( .A(n2023), .B(n2053), .CI(n1090), .CO(n1087), .S(n1088) );
  INV_X32 U944 ( .A(n1089), .ZN(n1090) );
  FA_X1 U945 ( .A(n1099), .B(n1096), .CI(n1094), .CO(n1091), .S(n1092) );
  FA_X1 U946 ( .A(n2115), .B(n2084), .CI(n1101), .CO(n1093), .S(n1094) );
  FA_X1 U947 ( .A(n2054), .B(n2024), .CI(n1103), .CO(n1095), .S(n1096) );
  FA_X1 U948 ( .A(n1100), .B(n1102), .CI(n1107), .CO(n1097), .S(n1098) );
  FA_X1 U949 ( .A(n1111), .B(n2085), .CI(n1109), .CO(n1099), .S(n1100) );
  FA_X1 U950 ( .A(n2055), .B(n2025), .CI(n1104), .CO(n1101), .S(n1102) );
  INV_X32 U951 ( .A(n1103), .ZN(n1104) );
  FA_X1 U952 ( .A(n1115), .B(n1117), .CI(n1108), .CO(n1105), .S(n1106) );
  FA_X1 U953 ( .A(n1112), .B(n1119), .CI(n1110), .CO(n1107), .S(n1108) );
  FA_X1 U954 ( .A(n2086), .B(n2056), .CI(n2147), .CO(n1109), .S(n1110) );
  FA_X1 U955 ( .A(n2116), .B(n2026), .CI(n1121), .CO(n1111), .S(n1112) );
  FA_X1 U956 ( .A(n1125), .B(n1118), .CI(n1116), .CO(n1113), .S(n1114) );
  FA_X1 U957 ( .A(n1120), .B(n1129), .CI(n1127), .CO(n1115), .S(n1116) );
  FA_X1 U958 ( .A(n2027), .B(n2087), .CI(n1131), .CO(n1117), .S(n1118) );
  FA_X1 U959 ( .A(n2117), .B(n2057), .CI(n1122), .CO(n1119), .S(n1120) );
  INV_X32 U960 ( .A(n1121), .ZN(n1122) );
  FA_X1 U961 ( .A(n1135), .B(n1128), .CI(n1126), .CO(n1123), .S(n1124) );
  FA_X1 U962 ( .A(n1132), .B(n1130), .CI(n1137), .CO(n1125), .S(n1126) );
  FA_X1 U963 ( .A(n1141), .B(n2179), .CI(n1139), .CO(n1127), .S(n1128) );
  FA_X1 U964 ( .A(n2058), .B(n2148), .CI(n2118), .CO(n1129), .S(n1130) );
  FA_X1 U965 ( .A(n1143), .B(n2028), .CI(n2088), .CO(n1131), .S(n1132) );
  FA_X1 U966 ( .A(n1147), .B(n1138), .CI(n1136), .CO(n1133), .S(n1134) );
  FA_X1 U967 ( .A(n1151), .B(n1142), .CI(n1149), .CO(n1135), .S(n1136) );
  FA_X1 U968 ( .A(n1153), .B(n1155), .CI(n1140), .CO(n1137), .S(n1138) );
  FA_X1 U969 ( .A(n2059), .B(n2029), .CI(n2119), .CO(n1139), .S(n1140) );
  FA_X1 U970 ( .A(n2149), .B(n2089), .CI(n1144), .CO(n1141), .S(n1142) );
  INV_X32 U971 ( .A(n1143), .ZN(n1144) );
  FA_X1 U972 ( .A(n1159), .B(n1150), .CI(n1148), .CO(n1145), .S(n1146) );
  FA_X1 U973 ( .A(n1152), .B(n1163), .CI(n1161), .CO(n1147), .S(n1148) );
  FA_X1 U974 ( .A(n1154), .B(n1165), .CI(n1156), .CO(n1149), .S(n1150) );
  FA_X1 U975 ( .A(n2211), .B(n2120), .CI(n1167), .CO(n1151), .S(n1152) );
  FA_X1 U976 ( .A(n2090), .B(n2150), .CI(n2180), .CO(n1153), .S(n1154) );
  FA_X1 U977 ( .A(n1169), .B(n2030), .CI(n2060), .CO(n1155), .S(n1156) );
  FA_X1 U978 ( .A(n1173), .B(n1162), .CI(n1160), .CO(n1157), .S(n1158) );
  FA_X1 U979 ( .A(n1164), .B(n1177), .CI(n1175), .CO(n1159), .S(n1160) );
  FA_X1 U980 ( .A(n1166), .B(n1179), .CI(n1168), .CO(n1161), .S(n1162) );
  FA_X1 U981 ( .A(n1183), .B(n2061), .CI(n1181), .CO(n1163), .S(n1164) );
  FA_X1 U982 ( .A(n2031), .B(n2151), .CI(n2121), .CO(n1165), .S(n1166) );
  FA_X1 U983 ( .A(n2181), .B(n2091), .CI(n1170), .CO(n1167), .S(n1168) );
  INV_X32 U984 ( .A(n1169), .ZN(n1170) );
  FA_X1 U985 ( .A(n1187), .B(n1176), .CI(n1174), .CO(n1171), .S(n1172) );
  FA_X1 U986 ( .A(n1178), .B(n1191), .CI(n1189), .CO(n1173), .S(n1174) );
  FA_X1 U987 ( .A(n1180), .B(n1184), .CI(n1193), .CO(n1175), .S(n1176) );
  FA_X1 U988 ( .A(n1195), .B(n1197), .CI(n1182), .CO(n1177), .S(n1178) );
  FA_X1 U989 ( .A(n2212), .B(n2062), .CI(n2243), .CO(n1179), .S(n1180) );
  FA_X1 U990 ( .A(n2122), .B(n2182), .CI(n2152), .CO(n1181), .S(n1182) );
  FA_X1 U991 ( .A(n1199), .B(n2032), .CI(n2092), .CO(n1183), .S(n1184) );
  FA_X1 U992 ( .A(n1203), .B(n1190), .CI(n1188), .CO(n1185), .S(n1186) );
  FA_X1 U993 ( .A(n1192), .B(n1207), .CI(n1205), .CO(n1187), .S(n1188) );
  FA_X1 U994 ( .A(n1209), .B(n1198), .CI(n1194), .CO(n1189), .S(n1190) );
  FA_X1 U995 ( .A(n1211), .B(n1213), .CI(n1196), .CO(n1191), .S(n1192) );
  FA_X1 U996 ( .A(n2123), .B(n2153), .CI(n1215), .CO(n1193), .S(n1194) );
  FA_X1 U997 ( .A(n2033), .B(n2183), .CI(n2063), .CO(n1195), .S(n1196) );
  FA_X1 U998 ( .A(n2213), .B(n2093), .CI(n1200), .CO(n1197), .S(n1198) );
  INV_X32 U999 ( .A(n1199), .ZN(n1200) );
  FA_X1 U1000 ( .A(n1219), .B(n1206), .CI(n1204), .CO(n1201), .S(n1202) );
  FA_X1 U1001 ( .A(n1208), .B(n1223), .CI(n1221), .CO(n1203), .S(n1204) );
  FA_X1 U1002 ( .A(n1225), .B(n1216), .CI(n1210), .CO(n1205), .S(n1206) );
  FA_X1 U1003 ( .A(n1212), .B(n1227), .CI(n1214), .CO(n1207), .S(n1208) );
  FA_X1 U1004 ( .A(n1231), .B(n2275), .CI(n1229), .CO(n1209), .S(n1210) );
  FA_X1 U1005 ( .A(n2184), .B(n2094), .CI(n2214), .CO(n1211), .S(n1212) );
  FA_X1 U1006 ( .A(n2064), .B(n2154), .CI(n2124), .CO(n1213), .S(n1214) );
  FA_X1 U1007 ( .A(n2244), .B(n2034), .CI(n1233), .CO(n1215), .S(n1216) );
  FA_X1 U1008 ( .A(n1237), .B(n1222), .CI(n1220), .CO(n1217), .S(n1218) );
  FA_X1 U1009 ( .A(n1224), .B(n1241), .CI(n1239), .CO(n1219), .S(n1220) );
  FA_X1 U1010 ( .A(n1243), .B(n1245), .CI(n1226), .CO(n1221), .S(n1222) );
  FA_X1 U1011 ( .A(n1232), .B(n1228), .CI(n1230), .CO(n1223), .S(n1224) );
  FA_X1 U1012 ( .A(n1247), .B(n1251), .CI(n1249), .CO(n1225), .S(n1226) );
  FA_X1 U1013 ( .A(n2095), .B(n2185), .CI(n2155), .CO(n1227), .S(n1228) );
  FA_X1 U1014 ( .A(n2065), .B(n2245), .CI(n2215), .CO(n1229), .S(n1230) );
  FA_X1 U1015 ( .A(n2035), .B(n2125), .CI(n1234), .CO(n1231), .S(n1232) );
  INV_X32 U1016 ( .A(n1233), .ZN(n1234) );
  FA_X1 U1017 ( .A(n1255), .B(n1240), .CI(n1238), .CO(n1235), .S(n1236) );
  FA_X1 U1018 ( .A(n1242), .B(n1259), .CI(n1257), .CO(n1237), .S(n1238) );
  FA_X1 U1019 ( .A(n1246), .B(n1261), .CI(n1244), .CO(n1239), .S(n1240) );
  FA_X1 U1020 ( .A(n1252), .B(n1250), .CI(n1263), .CO(n1241), .S(n1242) );
  FA_X1 U1021 ( .A(n1265), .B(n1267), .CI(n1248), .CO(n1243), .S(n1244) );
  FA_X1 U1022 ( .A(n2307), .B(n2246), .CI(n1269), .CO(n1245), .S(n1246) );
  FA_X1 U1023 ( .A(n2216), .B(n2126), .CI(n2156), .CO(n1247), .S(n1248) );
  FA_X1 U1024 ( .A(n2096), .B(n2186), .CI(n1271), .CO(n1249), .S(n1250) );
  FA_X1 U1025 ( .A(n2276), .B(n2036), .CI(n2066), .CO(n1251), .S(n1252) );
  FA_X1 U1026 ( .A(n1275), .B(n1258), .CI(n1256), .CO(n1253), .S(n1254) );
  FA_X1 U1027 ( .A(n1260), .B(n1279), .CI(n1277), .CO(n1255), .S(n1256) );
  FA_X1 U1028 ( .A(n1281), .B(n1264), .CI(n1262), .CO(n1257), .S(n1258) );
  FA_X1 U1029 ( .A(n1270), .B(n1268), .CI(n1283), .CO(n1259), .S(n1260) );
  FA_X1 U1030 ( .A(n1285), .B(n1287), .CI(n1266), .CO(n1261), .S(n1262) );
  FA_X1 U1031 ( .A(n1291), .B(n2187), .CI(n1289), .CO(n1263), .S(n1264) );
  FA_X1 U1032 ( .A(n2097), .B(n2217), .CI(n2157), .CO(n1265), .S(n1266) );
  FA_X1 U1033 ( .A(n2037), .B(n2247), .CI(n2067), .CO(n1267), .S(n1268) );
  FA_X1 U1034 ( .A(n2277), .B(n2127), .CI(n1272), .CO(n1269), .S(n1270) );
  INV_X32 U1035 ( .A(n1271), .ZN(n1272) );
  FA_X1 U1036 ( .A(n1295), .B(n1278), .CI(n1276), .CO(n1273), .S(n1274) );
  FA_X1 U1037 ( .A(n1280), .B(n1299), .CI(n1297), .CO(n1275), .S(n1276) );
  FA_X1 U1038 ( .A(n1284), .B(n1301), .CI(n1282), .CO(n1277), .S(n1278) );
  FA_X1 U1039 ( .A(n1305), .B(n1286), .CI(n1303), .CO(n1279), .S(n1280) );
  FA_X1 U1040 ( .A(n1292), .B(n1288), .CI(n1290), .CO(n1281), .S(n1282) );
  FA_X1 U1041 ( .A(n1307), .B(n1311), .CI(n1309), .CO(n1283), .S(n1284) );
  FA_X1 U1042 ( .A(n2248), .B(n2278), .CI(n2339), .CO(n1285), .S(n1286) );
  FA_X1 U1043 ( .A(n2218), .B(n2098), .CI(n2158), .CO(n1287), .S(n1288) );
  FA_X1 U1044 ( .A(n1313), .B(n2188), .CI(n2128), .CO(n1289), .S(n1290) );
  FA_X1 U1045 ( .A(n2308), .B(n2038), .CI(n2068), .CO(n1291), .S(n1292) );
  FA_X1 U1046 ( .A(n1317), .B(n1298), .CI(n1296), .CO(n1293), .S(n1294) );
  FA_X1 U1047 ( .A(n1300), .B(n1321), .CI(n1319), .CO(n1295), .S(n1296) );
  FA_X1 U1048 ( .A(n1304), .B(n1323), .CI(n1302), .CO(n1297), .S(n1298) );
  FA_X1 U1049 ( .A(n1325), .B(n1327), .CI(n1306), .CO(n1299), .S(n1300) );
  FA_X1 U1050 ( .A(n1312), .B(n1308), .CI(n1310), .CO(n1301), .S(n1302) );
  FA_X1 U1051 ( .A(n1329), .B(n1333), .CI(n1331), .CO(n1303), .S(n1304) );
  FA_X1 U1052 ( .A(n2249), .B(n2279), .CI(n1335), .CO(n1305), .S(n1306) );
  FA_X1 U1053 ( .A(n2129), .B(n2219), .CI(n2189), .CO(n1307), .S(n1308) );
  FA_X1 U1054 ( .A(n2069), .B(n2309), .CI(n2099), .CO(n1309), .S(n1310) );
  FA_X1 U1055 ( .A(n2039), .B(n2159), .CI(n1314), .CO(n1311), .S(n1312) );
  INV_X32 U1056 ( .A(n1313), .ZN(n1314) );
  FA_X1 U1057 ( .A(n1339), .B(n1320), .CI(n1318), .CO(n1315), .S(n1316) );
  FA_X1 U1058 ( .A(n1322), .B(n1343), .CI(n1341), .CO(n1317), .S(n1318) );
  FA_X1 U1059 ( .A(n1345), .B(n1326), .CI(n1324), .CO(n1319), .S(n1320) );
  FA_X1 U1060 ( .A(n1328), .B(n1349), .CI(n1347), .CO(n1321), .S(n1322) );
  FA_X1 U1061 ( .A(n1336), .B(n1332), .CI(n1334), .CO(n1323), .S(n1324) );
  FA_X1 U1062 ( .A(n1351), .B(n1353), .CI(n1330), .CO(n1325), .S(n1326) );
  FA_X1 U1063 ( .A(n1357), .B(n2371), .CI(n1355), .CO(n1327), .S(n1328) );
  FA_X1 U1064 ( .A(n2190), .B(n2340), .CI(n2310), .CO(n1329), .S(n1330) );
  FA_X1 U1065 ( .A(n2160), .B(n2280), .CI(n2250), .CO(n1331), .S(n1332) );
  FA_X1 U1066 ( .A(n2130), .B(n2220), .CI(n2070), .CO(n1333), .S(n1334) );
  FA_X1 U1067 ( .A(n1359), .B(n2040), .CI(n2100), .CO(n1335), .S(n1336) );
  FA_X1 U1068 ( .A(n1363), .B(n1342), .CI(n1340), .CO(n1337), .S(n1338) );
  FA_X1 U1069 ( .A(n1344), .B(n1367), .CI(n1365), .CO(n1339), .S(n1340) );
  FA_X1 U1070 ( .A(n1369), .B(n1348), .CI(n1346), .CO(n1341), .S(n1342) );
  FA_X1 U1071 ( .A(n1371), .B(n1373), .CI(n1350), .CO(n1343), .S(n1344) );
  FA_X1 U1072 ( .A(n1358), .B(n1356), .CI(n1375), .CO(n1345), .S(n1346) );
  FA_X1 U1073 ( .A(n1352), .B(n1381), .CI(n1354), .CO(n1347), .S(n1348) );
  FA_X1 U1074 ( .A(n1377), .B(n1383), .CI(n1379), .CO(n1349), .S(n1350) );
  FA_X1 U1075 ( .A(n2221), .B(n2281), .CI(n2251), .CO(n1351), .S(n1352) );
  FA_X1 U1076 ( .A(n2311), .B(n2131), .CI(n2161), .CO(n1353), .S(n1354) );
  FA_X1 U1077 ( .A(n2071), .B(n2341), .CI(n2101), .CO(n1355), .S(n1356) );
  FA_X1 U1078 ( .A(n2041), .B(n2191), .CI(n1360), .CO(n1357), .S(n1358) );
  INV_X32 U1079 ( .A(n1359), .ZN(n1360) );
  FA_X1 U1080 ( .A(n1387), .B(n1366), .CI(n1364), .CO(n1361), .S(n1362) );
  FA_X1 U1081 ( .A(n1368), .B(n1391), .CI(n1389), .CO(n1363), .S(n1364) );
  FA_X1 U1082 ( .A(n1393), .B(n1372), .CI(n1370), .CO(n1365), .S(n1366) );
  FA_X1 U1083 ( .A(n1395), .B(n1376), .CI(n1374), .CO(n1367), .S(n1368) );
  FA_X1 U1084 ( .A(n1399), .B(n1380), .CI(n1397), .CO(n1369), .S(n1370) );
  FA_X1 U1085 ( .A(n1384), .B(n1378), .CI(n1382), .CO(n1371), .S(n1372) );
  FA_X1 U1086 ( .A(n1403), .B(n1401), .CI(n1405), .CO(n1373), .S(n1374) );
  FA_X1 U1087 ( .A(n2403), .B(n2342), .CI(n1407), .CO(n1375), .S(n1376) );
  FA_X1 U1088 ( .A(n2072), .B(n2312), .CI(n2282), .CO(n1377), .S(n1378) );
  FA_X1 U1089 ( .A(n2162), .B(n2252), .CI(n2192), .CO(n1379), .S(n1380) );
  FA_X1 U1090 ( .A(n2102), .B(n2222), .CI(n2132), .CO(n1381), .S(n1382) );
  FA_X1 U1091 ( .A(n2372), .B(n2042), .CI(n1409), .CO(n1383), .S(n1384) );
  FA_X1 U1092 ( .A(n1413), .B(n1390), .CI(n1388), .CO(n1385), .S(n1386) );
  FA_X1 U1093 ( .A(n1392), .B(n1417), .CI(n1415), .CO(n1387), .S(n1388) );
  FA_X1 U1094 ( .A(n1419), .B(n1396), .CI(n1394), .CO(n1389), .S(n1390) );
  FA_X1 U1095 ( .A(n1398), .B(n1423), .CI(n1421), .CO(n1391), .S(n1392) );
  FA_X1 U1096 ( .A(n1425), .B(n1404), .CI(n1400), .CO(n1393), .S(n1394) );
  FA_X1 U1097 ( .A(n1408), .B(n1402), .CI(n1406), .CO(n1395), .S(n1396) );
  FA_X1 U1098 ( .A(n1429), .B(n1431), .CI(n1427), .CO(n1397), .S(n1398) );
  FA_X1 U1099 ( .A(n1435), .B(n2253), .CI(n1433), .CO(n1399), .S(n1400) );
  FA_X1 U1100 ( .A(n2163), .B(n2283), .CI(n2223), .CO(n1401), .S(n1402) );
  FA_X1 U1101 ( .A(n2103), .B(n2313), .CI(n2133), .CO(n1403), .S(n1404) );
  FA_X1 U1102 ( .A(n2043), .B(n2343), .CI(n2073), .CO(n1405), .S(n1406) );
  FA_X1 U1103 ( .A(n2373), .B(n2193), .CI(n1410), .CO(n1407), .S(n1408) );
  INV_X32 U1104 ( .A(n1409), .ZN(n1410) );
  FA_X1 U1105 ( .A(n1439), .B(n1416), .CI(n1414), .CO(n1411), .S(n1412) );
  FA_X1 U1106 ( .A(n1418), .B(n1443), .CI(n1441), .CO(n1413), .S(n1414) );
  FA_X1 U1107 ( .A(n1445), .B(n1422), .CI(n1420), .CO(n1415), .S(n1416) );
  FA_X1 U1108 ( .A(n1424), .B(n1426), .CI(n1447), .CO(n1417), .S(n1418) );
  FA_X1 U1109 ( .A(n1451), .B(n1453), .CI(n1449), .CO(n1419), .S(n1420) );
  FA_X1 U1110 ( .A(n1436), .B(n1434), .CI(n1428), .CO(n1421), .S(n1422) );
  FA_X1 U1111 ( .A(n1430), .B(n1455), .CI(n1432), .CO(n1423), .S(n1424) );
  FA_X1 U1112 ( .A(n1461), .B(n1457), .CI(n1459), .CO(n1425), .S(n1426) );
  FA_X1 U1113 ( .A(n2344), .B(n2374), .CI(n2435), .CO(n1427), .S(n1428) );
  FA_X1 U1114 ( .A(n2314), .B(n2194), .CI(n2224), .CO(n1429), .S(n1430) );
  FA_X1 U1115 ( .A(n1463), .B(n2284), .CI(n2164), .CO(n1431), .S(n1432) );
  FA_X1 U1116 ( .A(n2104), .B(n2254), .CI(n2134), .CO(n1433), .S(n1434) );
  FA_X1 U1117 ( .A(n2404), .B(n2044), .CI(n2074), .CO(n1435), .S(n1436) );
  FA_X1 U1118 ( .A(n1467), .B(n1442), .CI(n1440), .CO(n1437), .S(n1438) );
  FA_X1 U1119 ( .A(n1444), .B(n1471), .CI(n1469), .CO(n1439), .S(n1440) );
  FA_X1 U1120 ( .A(n1473), .B(n1448), .CI(n1446), .CO(n1441), .S(n1442) );
  FA_X1 U1121 ( .A(n1450), .B(n1452), .CI(n1475), .CO(n1443), .S(n1444) );
  FA_X1 U1122 ( .A(n1454), .B(n1479), .CI(n1477), .CO(n1445), .S(n1446) );
  FA_X1 U1123 ( .A(n1460), .B(n1462), .CI(n1481), .CO(n1447), .S(n1448) );
  FA_X1 U1124 ( .A(n1456), .B(n1487), .CI(n1458), .CO(n1449), .S(n1450) );
  FA_X1 U1125 ( .A(n1489), .B(n1485), .CI(n1483), .CO(n1451), .S(n1452) );
  FA_X1 U1126 ( .A(n2285), .B(n2315), .CI(n1491), .CO(n1453), .S(n1454) );
  FA_X1 U1127 ( .A(n2165), .B(n2345), .CI(n2195), .CO(n1455), .S(n1456) );
  FA_X1 U1128 ( .A(n2135), .B(n2405), .CI(n2375), .CO(n1457), .S(n1458) );
  FA_X1 U1129 ( .A(n2075), .B(n2255), .CI(n2105), .CO(n1459), .S(n1460) );
  FA_X1 U1130 ( .A(n2045), .B(n2225), .CI(n1464), .CO(n1461), .S(n1462) );
  INV_X32 U1131 ( .A(n1463), .ZN(n1464) );
  FA_X1 U1132 ( .A(n1495), .B(n1470), .CI(n1468), .CO(n1465), .S(n1466) );
  FA_X1 U1133 ( .A(n1472), .B(n1499), .CI(n1497), .CO(n1467), .S(n1468) );
  FA_X1 U1134 ( .A(n1501), .B(n1476), .CI(n1474), .CO(n1469), .S(n1470) );
  FA_X1 U1135 ( .A(n1503), .B(n1480), .CI(n1478), .CO(n1471), .S(n1472) );
  FA_X1 U1136 ( .A(n1482), .B(n1507), .CI(n1505), .CO(n1473), .S(n1474) );
  FA_X1 U1137 ( .A(n1486), .B(n1488), .CI(n1509), .CO(n1475), .S(n1476) );
  FA_X1 U1138 ( .A(n1492), .B(n1484), .CI(n1490), .CO(n1477), .S(n1478) );
  FA_X1 U1139 ( .A(n1515), .B(n1511), .CI(n1513), .CO(n1479), .S(n1480) );
  FA_X1 U1140 ( .A(n1519), .B(n2467), .CI(n1517), .CO(n1481), .S(n1482) );
  FA_X1 U1141 ( .A(n2436), .B(n2406), .CI(n2256), .CO(n1483), .S(n1484) );
  FA_X1 U1142 ( .A(n2346), .B(n2226), .CI(n2376), .CO(n1485), .S(n1486) );
  FA_X1 U1143 ( .A(n2196), .B(n2316), .CI(n2136), .CO(n1487), .S(n1488) );
  FA_X1 U1144 ( .A(n2106), .B(n2286), .CI(n2166), .CO(n1489), .S(n1490) );
  FA_X1 U1145 ( .A(n1521), .B(n2046), .CI(n2076), .CO(n1491), .S(n1492) );
  FA_X1 U1146 ( .A(n1525), .B(n1498), .CI(n1496), .CO(n1493), .S(n1494) );
  FA_X1 U1147 ( .A(n1500), .B(n1502), .CI(n1527), .CO(n1495), .S(n1496) );
  FA_X1 U1148 ( .A(n1531), .B(n1504), .CI(n1529), .CO(n1497), .S(n1498) );
  FA_X1 U1149 ( .A(n1533), .B(n1508), .CI(n1506), .CO(n1499), .S(n1500) );
  FA_X1 U1150 ( .A(n1510), .B(n1537), .CI(n1535), .CO(n1501), .S(n1502) );
  FA_X1 U1151 ( .A(n1516), .B(n1514), .CI(n1539), .CO(n1503), .S(n1504) );
  FA_X1 U1152 ( .A(n1520), .B(n1512), .CI(n1518), .CO(n1505), .S(n1506) );
  FA_X1 U1153 ( .A(n1543), .B(n1545), .CI(n1541), .CO(n1507), .S(n1508) );
  FA_X1 U1154 ( .A(n1549), .B(n1551), .CI(n1547), .CO(n1509), .S(n1510) );
  FA_X1 U1155 ( .A(n2287), .B(n2347), .CI(n2317), .CO(n1511), .S(n1512) );
  FA_X1 U1156 ( .A(n2167), .B(n2377), .CI(n2197), .CO(n1513), .S(n1514) );
  FA_X1 U1157 ( .A(n2107), .B(n2407), .CI(n2137), .CO(n1515), .S(n1516) );
  FA_X1 U1158 ( .A(n2437), .B(n2257), .CI(n2077), .CO(n1517), .S(n1518) );
  FA_X1 U1159 ( .A(n2047), .B(n2227), .CI(n1522), .CO(n1519), .S(n1520) );
  INV_X32 U1160 ( .A(n1521), .ZN(n1522) );
  FA_X1 U1161 ( .A(n1555), .B(n1528), .CI(n1526), .CO(n1523), .S(n1524) );
  FA_X1 U1162 ( .A(n1530), .B(n1532), .CI(n1557), .CO(n1525), .S(n1526) );
  FA_X1 U1163 ( .A(n1561), .B(n1534), .CI(n1559), .CO(n1527), .S(n1528) );
  FA_X1 U1164 ( .A(n1563), .B(n1538), .CI(n1536), .CO(n1529), .S(n1530) );
  FA_X1 U1165 ( .A(n1540), .B(n1567), .CI(n1565), .CO(n1531), .S(n1532) );
  FA_X1 U1166 ( .A(n1542), .B(n1546), .CI(n1569), .CO(n1533), .S(n1534) );
  FA_X1 U1167 ( .A(n1550), .B(n1548), .CI(n1544), .CO(n1535), .S(n1536) );
  FA_X1 U1168 ( .A(n1579), .B(n1571), .CI(n1577), .CO(n1537), .S(n1538) );
  FA_X1 U1169 ( .A(n1573), .B(n1552), .CI(n1575), .CO(n1539), .S(n1540) );
  FA_X1 U1170 ( .A(n2499), .B(n2408), .CI(n1581), .CO(n1541), .S(n1542) );
  FA_X1 U1171 ( .A(n2378), .B(n2438), .CI(n2468), .CO(n1543), .S(n1544) );
  FA_X1 U1172 ( .A(n2198), .B(n2348), .CI(n2228), .CO(n1545), .S(n1546) );
  FA_X1 U1173 ( .A(n2138), .B(n2288), .CI(n2168), .CO(n1547), .S(n1548) );
  FA_X1 U1174 ( .A(n2048), .B(n2258), .CI(n2108), .CO(n1549), .S(n1550) );
  XNOR2_X2 U1175 ( .A(n2318), .B(n2078), .ZN(n1552) );
  OR2_X4 U1176 ( .A1(n2318), .A2(n2078), .ZN(n1551) );
  FA_X1 U1177 ( .A(n1585), .B(n1558), .CI(n1556), .CO(n1553), .S(n1554) );
  FA_X1 U1178 ( .A(n1560), .B(n1562), .CI(n1587), .CO(n1555), .S(n1556) );
  FA_X1 U1179 ( .A(n1591), .B(n1564), .CI(n1589), .CO(n1557), .S(n1558) );
  FA_X1 U1180 ( .A(n1593), .B(n1568), .CI(n1566), .CO(n1559), .S(n1560) );
  FA_X1 U1181 ( .A(n1570), .B(n1597), .CI(n1595), .CO(n1561), .S(n1562) );
  FA_X1 U1182 ( .A(n1574), .B(n1576), .CI(n1599), .CO(n1563), .S(n1564) );
  FA_X1 U1183 ( .A(n1580), .B(n1572), .CI(n1578), .CO(n1565), .S(n1566) );
  FA_X1 U1184 ( .A(n1605), .B(n1601), .CI(n1603), .CO(n1567), .S(n1568) );
  FA_X1 U1185 ( .A(n1609), .B(n1582), .CI(n1607), .CO(n1569), .S(n1570) );
  FA_X1 U1186 ( .A(n2319), .B(n2199), .CI(n2259), .CO(n1571), .S(n1572) );
  FA_X1 U1187 ( .A(n2109), .B(n2349), .CI(n2139), .CO(n1573), .S(n1574) );
  FA_X1 U1188 ( .A(n2079), .B(n2169), .CI(n2379), .CO(n1575), .S(n1576) );
  FA_X1 U1189 ( .A(n2439), .B(n2229), .CI(n2409), .CO(n1577), .S(n1578) );
  FA_X1 U1190 ( .A(n2500), .B(n2289), .CI(n2469), .CO(n1579), .S(n1580) );
  HA_X1 U1191 ( .A(n2049), .B(n2003), .CO(n1581), .S(n1582) );
  FA_X1 U1192 ( .A(n1613), .B(n1588), .CI(n1586), .CO(n1583), .S(n1584) );
  FA_X1 U1193 ( .A(n1590), .B(n1592), .CI(n1615), .CO(n1585), .S(n1586) );
  FA_X1 U1194 ( .A(n1619), .B(n1594), .CI(n1617), .CO(n1587), .S(n1588) );
  FA_X1 U1195 ( .A(n1598), .B(n1621), .CI(n1596), .CO(n1589), .S(n1590) );
  FA_X1 U1196 ( .A(n1623), .B(n1625), .CI(n1600), .CO(n1591), .S(n1592) );
  FA_X1 U1197 ( .A(n1606), .B(n1604), .CI(n1627), .CO(n1593), .S(n1594) );
  FA_X1 U1198 ( .A(n1610), .B(n1602), .CI(n1608), .CO(n1595), .S(n1596) );
  FA_X1 U1199 ( .A(n1633), .B(n1629), .CI(n1631), .CO(n1597), .S(n1598) );
  FA_X1 U1200 ( .A(n1637), .B(n2350), .CI(n1635), .CO(n1599), .S(n1600) );
  FA_X1 U1201 ( .A(n2290), .B(n2380), .CI(n2320), .CO(n1601), .S(n1602) );
  FA_X1 U1202 ( .A(n2230), .B(n2200), .CI(n2260), .CO(n1603), .S(n1604) );
  FA_X1 U1203 ( .A(n2140), .B(n2410), .CI(n2170), .CO(n1605), .S(n1606) );
  FA_X1 U1204 ( .A(n2110), .B(n2470), .CI(n2440), .CO(n1607), .S(n1608) );
  FA_X1 U1205 ( .A(n2080), .B(n2501), .CI(n2050), .CO(n1609), .S(n1610) );
  FA_X1 U1206 ( .A(n1641), .B(n1616), .CI(n1614), .CO(n1611), .S(n1612) );
  FA_X1 U1207 ( .A(n1618), .B(n1620), .CI(n1643), .CO(n1613), .S(n1614) );
  FA_X1 U1208 ( .A(n1647), .B(n1622), .CI(n1645), .CO(n1615), .S(n1616) );
  FA_X1 U1209 ( .A(n1626), .B(n1649), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1210 ( .A(n1628), .B(n1653), .CI(n1651), .CO(n1619), .S(n1620) );
  FA_X1 U1211 ( .A(n1632), .B(n1634), .CI(n1636), .CO(n1621), .S(n1622) );
  FA_X1 U1212 ( .A(n1655), .B(n1659), .CI(n1630), .CO(n1623), .S(n1624) );
  FA_X1 U1213 ( .A(n1663), .B(n1657), .CI(n1661), .CO(n1625), .S(n1626) );
  FA_X1 U1214 ( .A(n2381), .B(n2351), .CI(n1638), .CO(n1627), .S(n1628) );
  FA_X1 U1215 ( .A(n2201), .B(n2411), .CI(n2231), .CO(n1629), .S(n1630) );
  FA_X1 U1216 ( .A(n2441), .B(n2321), .CI(n2171), .CO(n1631), .S(n1632) );
  FA_X1 U1217 ( .A(n2471), .B(n2261), .CI(n2141), .CO(n1633), .S(n1634) );
  FA_X1 U1218 ( .A(n2502), .B(n2291), .CI(n2111), .CO(n1635), .S(n1636) );
  HA_X1 U1219 ( .A(n2081), .B(n2004), .CO(n1637), .S(n1638) );
  FA_X1 U1220 ( .A(n1667), .B(n1644), .CI(n1642), .CO(n1639), .S(n1640) );
  FA_X1 U1221 ( .A(n1646), .B(n1671), .CI(n1669), .CO(n1641), .S(n1642) );
  FA_X1 U1222 ( .A(n1673), .B(n1650), .CI(n1648), .CO(n1643), .S(n1644) );
  FA_X1 U1223 ( .A(n1675), .B(n1654), .CI(n1652), .CO(n1645), .S(n1646) );
  FA_X1 U1224 ( .A(n1679), .B(n1660), .CI(n1677), .CO(n1647), .S(n1648) );
  FA_X1 U1225 ( .A(n1664), .B(n1658), .CI(n1662), .CO(n1649), .S(n1650) );
  FA_X1 U1226 ( .A(n1683), .B(n1681), .CI(n1656), .CO(n1651), .S(n1652) );
  FA_X1 U1227 ( .A(n1687), .B(n1689), .CI(n1685), .CO(n1653), .S(n1654) );
  FA_X1 U1228 ( .A(n2292), .B(n2352), .CI(n2322), .CO(n1655), .S(n1656) );
  FA_X1 U1229 ( .A(n2232), .B(n2382), .CI(n2262), .CO(n1657), .S(n1658) );
  FA_X1 U1230 ( .A(n2172), .B(n2412), .CI(n2202), .CO(n1659), .S(n1660) );
  FA_X1 U1231 ( .A(n2142), .B(n2472), .CI(n2442), .CO(n1661), .S(n1662) );
  FA_X1 U1232 ( .A(n2112), .B(n2503), .CI(n2082), .CO(n1663), .S(n1664) );
  FA_X1 U1233 ( .A(n1693), .B(n1670), .CI(n1668), .CO(n1665), .S(n1666) );
  FA_X1 U1234 ( .A(n1672), .B(n1674), .CI(n1695), .CO(n1667), .S(n1668) );
  FA_X1 U1235 ( .A(n1676), .B(n1699), .CI(n1697), .CO(n1669), .S(n1670) );
  FA_X1 U1236 ( .A(n1701), .B(n1680), .CI(n1678), .CO(n1671), .S(n1672) );
  FA_X1 U1237 ( .A(n1686), .B(n1688), .CI(n1703), .CO(n1673), .S(n1674) );
  FA_X1 U1238 ( .A(n1682), .B(n1705), .CI(n1684), .CO(n1675), .S(n1676) );
  FA_X1 U1239 ( .A(n1709), .B(n1707), .CI(n1711), .CO(n1677), .S(n1678) );
  FA_X1 U1240 ( .A(n1690), .B(n2413), .CI(n1713), .CO(n1679), .S(n1680) );
  FA_X1 U1241 ( .A(n2353), .B(n2443), .CI(n2383), .CO(n1681), .S(n1682) );
  FA_X1 U1242 ( .A(n2473), .B(n2263), .CI(n2233), .CO(n1683), .S(n1684) );
  FA_X1 U1243 ( .A(n2173), .B(n2293), .CI(n2203), .CO(n1685), .S(n1686) );
  FA_X1 U1244 ( .A(n2143), .B(n2323), .CI(n2504), .CO(n1687), .S(n1688) );
  HA_X1 U1245 ( .A(n2113), .B(n2005), .CO(n1689), .S(n1690) );
  FA_X1 U1246 ( .A(n1717), .B(n1696), .CI(n1694), .CO(n1691), .S(n1692) );
  FA_X1 U1247 ( .A(n1719), .B(n1721), .CI(n1698), .CO(n1693), .S(n1694) );
  FA_X1 U1248 ( .A(n1702), .B(n1704), .CI(n1700), .CO(n1695), .S(n1696) );
  FA_X1 U1249 ( .A(n1725), .B(n1727), .CI(n1723), .CO(n1697), .S(n1698) );
  FA_X1 U1250 ( .A(n1712), .B(n1714), .CI(n1706), .CO(n1699), .S(n1700) );
  FA_X1 U1251 ( .A(n1708), .B(n1735), .CI(n1710), .CO(n1701), .S(n1702) );
  FA_X1 U1252 ( .A(n1729), .B(n1731), .CI(n1733), .CO(n1703), .S(n1704) );
  FA_X1 U1253 ( .A(n2354), .B(n2384), .CI(n1737), .CO(n1705), .S(n1706) );
  FA_X1 U1254 ( .A(n2294), .B(n2414), .CI(n2324), .CO(n1707), .S(n1708) );
  FA_X1 U1255 ( .A(n2234), .B(n2444), .CI(n2264), .CO(n1709), .S(n1710) );
  FA_X1 U1256 ( .A(n2174), .B(n2474), .CI(n2204), .CO(n1711), .S(n1712) );
  FA_X1 U1257 ( .A(n2144), .B(n2505), .CI(n2114), .CO(n1713), .S(n1714) );
  FA_X1 U1258 ( .A(n1741), .B(n1720), .CI(n1718), .CO(n1715), .S(n1716) );
  FA_X1 U1259 ( .A(n1722), .B(n1745), .CI(n1743), .CO(n1717), .S(n1718) );
  FA_X1 U1260 ( .A(n1726), .B(n1747), .CI(n1724), .CO(n1719), .S(n1720) );
  FA_X1 U1261 ( .A(n1749), .B(n1751), .CI(n1728), .CO(n1721), .S(n1722) );
  FA_X1 U1262 ( .A(n1736), .B(n1732), .CI(n1734), .CO(n1723), .S(n1724) );
  FA_X1 U1263 ( .A(n1753), .B(n1755), .CI(n1730), .CO(n1725), .S(n1726) );
  FA_X1 U1264 ( .A(n1759), .B(n1738), .CI(n1757), .CO(n1727), .S(n1728) );
  FA_X1 U1265 ( .A(n2265), .B(n2385), .CI(n2355), .CO(n1729), .S(n1730) );
  FA_X1 U1266 ( .A(n2205), .B(n2415), .CI(n2235), .CO(n1731), .S(n1732) );
  FA_X1 U1267 ( .A(n2475), .B(n2295), .CI(n2445), .CO(n1733), .S(n1734) );
  FA_X1 U1268 ( .A(n2506), .B(n2325), .CI(n2175), .CO(n1735), .S(n1736) );
  HA_X1 U1269 ( .A(n2145), .B(n2006), .CO(n1737), .S(n1738) );
  FA_X1 U1270 ( .A(n1763), .B(n1744), .CI(n1742), .CO(n1739), .S(n1740) );
  FA_X1 U1271 ( .A(n1746), .B(n1767), .CI(n1765), .CO(n1741), .S(n1742) );
  FA_X1 U1272 ( .A(n1750), .B(n1769), .CI(n1748), .CO(n1743), .S(n1744) );
  FA_X1 U1273 ( .A(n1771), .B(n1773), .CI(n1752), .CO(n1745), .S(n1746) );
  FA_X1 U1274 ( .A(n1760), .B(n1756), .CI(n1758), .CO(n1747), .S(n1748) );
  FA_X1 U1275 ( .A(n1775), .B(n1777), .CI(n1754), .CO(n1749), .S(n1750) );
  FA_X1 U1276 ( .A(n1781), .B(n2356), .CI(n1779), .CO(n1751), .S(n1752) );
  FA_X1 U1277 ( .A(n2296), .B(n2386), .CI(n2326), .CO(n1753), .S(n1754) );
  FA_X1 U1278 ( .A(n2266), .B(n2446), .CI(n2416), .CO(n1755), .S(n1756) );
  FA_X1 U1279 ( .A(n2206), .B(n2476), .CI(n2236), .CO(n1757), .S(n1758) );
  FA_X1 U1280 ( .A(n2176), .B(n2507), .CI(n2146), .CO(n1759), .S(n1760) );
  FA_X1 U1281 ( .A(n1785), .B(n1766), .CI(n1764), .CO(n1761), .S(n1762) );
  FA_X1 U1282 ( .A(n1787), .B(n1770), .CI(n1768), .CO(n1763), .S(n1764) );
  FA_X1 U1283 ( .A(n1772), .B(n1791), .CI(n1789), .CO(n1765), .S(n1766) );
  FA_X1 U1284 ( .A(n1793), .B(n1780), .CI(n1774), .CO(n1767), .S(n1768) );
  FA_X1 U1285 ( .A(n1776), .B(n1799), .CI(n1778), .CO(n1769), .S(n1770) );
  FA_X1 U1286 ( .A(n1795), .B(n1801), .CI(n1797), .CO(n1771), .S(n1772) );
  FA_X1 U1287 ( .A(n2387), .B(n2417), .CI(n1782), .CO(n1773), .S(n1774) );
  FA_X1 U1288 ( .A(n2267), .B(n2447), .CI(n2297), .CO(n1775), .S(n1776) );
  FA_X1 U1289 ( .A(n2477), .B(n2327), .CI(n2237), .CO(n1777), .S(n1778) );
  FA_X1 U1290 ( .A(n2508), .B(n2357), .CI(n2207), .CO(n1779), .S(n1780) );
  HA_X1 U1291 ( .A(n2177), .B(n2007), .CO(n1781), .S(n1782) );
  FA_X1 U1292 ( .A(n1805), .B(n1788), .CI(n1786), .CO(n1783), .S(n1784) );
  FA_X1 U1293 ( .A(n1790), .B(n1792), .CI(n1807), .CO(n1785), .S(n1786) );
  FA_X1 U1294 ( .A(n1794), .B(n1811), .CI(n1809), .CO(n1787), .S(n1788) );
  FA_X1 U1295 ( .A(n1802), .B(n1800), .CI(n1813), .CO(n1789), .S(n1790) );
  FA_X1 U1296 ( .A(n1796), .B(n1815), .CI(n1798), .CO(n1791), .S(n1792) );
  FA_X1 U1297 ( .A(n1819), .B(n1821), .CI(n1817), .CO(n1793), .S(n1794) );
  FA_X1 U1298 ( .A(n2358), .B(n2418), .CI(n2388), .CO(n1795), .S(n1796) );
  FA_X1 U1299 ( .A(n2298), .B(n2448), .CI(n2328), .CO(n1797), .S(n1798) );
  FA_X1 U1300 ( .A(n2238), .B(n2478), .CI(n2268), .CO(n1799), .S(n1800) );
  FA_X1 U1301 ( .A(n2208), .B(n2509), .CI(n2178), .CO(n1801), .S(n1802) );
  FA_X1 U1302 ( .A(n1825), .B(n1808), .CI(n1806), .CO(n1803), .S(n1804) );
  FA_X1 U1303 ( .A(n1810), .B(n1812), .CI(n1827), .CO(n1805), .S(n1806) );
  FA_X1 U1304 ( .A(n1814), .B(n1831), .CI(n1829), .CO(n1807), .S(n1808) );
  FA_X1 U1305 ( .A(n1820), .B(n1816), .CI(n1818), .CO(n1809), .S(n1810) );
  FA_X1 U1306 ( .A(n1835), .B(n1837), .CI(n1833), .CO(n1811), .S(n1812) );
  FA_X1 U1307 ( .A(n1822), .B(n2389), .CI(n1839), .CO(n1813), .S(n1814) );
  FA_X1 U1308 ( .A(n2269), .B(n2419), .CI(n2299), .CO(n1815), .S(n1816) );
  FA_X1 U1309 ( .A(n2239), .B(n2329), .CI(n2449), .CO(n1817), .S(n1818) );
  FA_X1 U1310 ( .A(n2510), .B(n2359), .CI(n2479), .CO(n1819), .S(n1820) );
  HA_X1 U1311 ( .A(n2209), .B(n2008), .CO(n1821), .S(n1822) );
  FA_X1 U1312 ( .A(n1843), .B(n1828), .CI(n1826), .CO(n1823), .S(n1824) );
  FA_X1 U1313 ( .A(n1830), .B(n1832), .CI(n1845), .CO(n1825), .S(n1826) );
  FA_X1 U1314 ( .A(n1849), .B(n1834), .CI(n1847), .CO(n1827), .S(n1828) );
  FA_X1 U1315 ( .A(n1840), .B(n1836), .CI(n1838), .CO(n1829), .S(n1830) );
  FA_X1 U1316 ( .A(n1851), .B(n1855), .CI(n1853), .CO(n1831), .S(n1832) );
  FA_X1 U1317 ( .A(n2390), .B(n2420), .CI(n1857), .CO(n1833), .S(n1834) );
  FA_X1 U1318 ( .A(n2330), .B(n2450), .CI(n2360), .CO(n1835), .S(n1836) );
  FA_X1 U1319 ( .A(n2270), .B(n2480), .CI(n2300), .CO(n1837), .S(n1838) );
  FA_X1 U1320 ( .A(n2240), .B(n2511), .CI(n2210), .CO(n1839), .S(n1840) );
  FA_X1 U1321 ( .A(n1861), .B(n1846), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1322 ( .A(n1848), .B(n1865), .CI(n1863), .CO(n1843), .S(n1844) );
  FA_X1 U1323 ( .A(n1867), .B(n1856), .CI(n1850), .CO(n1845), .S(n1846) );
  FA_X1 U1324 ( .A(n1852), .B(n1869), .CI(n1854), .CO(n1847), .S(n1848) );
  FA_X1 U1325 ( .A(n1873), .B(n1858), .CI(n1871), .CO(n1849), .S(n1850) );
  FA_X1 U1326 ( .A(n2361), .B(n2481), .CI(n2451), .CO(n1851), .S(n1852) );
  FA_X1 U1327 ( .A(n2512), .B(n2421), .CI(n2331), .CO(n1853), .S(n1854) );
  FA_X1 U1328 ( .A(n2271), .B(n2391), .CI(n2301), .CO(n1855), .S(n1856) );
  HA_X1 U1329 ( .A(n2241), .B(n2009), .CO(n1857), .S(n1858) );
  FA_X1 U1330 ( .A(n1877), .B(n1864), .CI(n1862), .CO(n1859), .S(n1860) );
  FA_X1 U1331 ( .A(n1866), .B(n1868), .CI(n1879), .CO(n1861), .S(n1862) );
  FA_X1 U1332 ( .A(n1883), .B(n1874), .CI(n1881), .CO(n1863), .S(n1864) );
  FA_X1 U1333 ( .A(n1870), .B(n1885), .CI(n1872), .CO(n1865), .S(n1866) );
  FA_X1 U1334 ( .A(n1889), .B(n2422), .CI(n1887), .CO(n1867), .S(n1868) );
  FA_X1 U1335 ( .A(n2362), .B(n2452), .CI(n2392), .CO(n1869), .S(n1870) );
  FA_X1 U1336 ( .A(n2302), .B(n2482), .CI(n2332), .CO(n1871), .S(n1872) );
  FA_X1 U1337 ( .A(n2272), .B(n2513), .CI(n2242), .CO(n1873), .S(n1874) );
  FA_X1 U1338 ( .A(n1880), .B(n1893), .CI(n1878), .CO(n1875), .S(n1876) );
  FA_X1 U1339 ( .A(n1895), .B(n1884), .CI(n1882), .CO(n1877), .S(n1878) );
  FA_X1 U1340 ( .A(n1888), .B(n1886), .CI(n1897), .CO(n1879), .S(n1880) );
  FA_X1 U1341 ( .A(n1899), .B(n1903), .CI(n1901), .CO(n1881), .S(n1882) );
  FA_X1 U1342 ( .A(n2453), .B(n2483), .CI(n1890), .CO(n1883), .S(n1884) );
  FA_X1 U1343 ( .A(n2333), .B(n2423), .CI(n2363), .CO(n1885), .S(n1886) );
  FA_X1 U1344 ( .A(n2303), .B(n2393), .CI(n2514), .CO(n1887), .S(n1888) );
  HA_X1 U1345 ( .A(n2273), .B(n2010), .CO(n1889), .S(n1890) );
  FA_X1 U1346 ( .A(n1907), .B(n1896), .CI(n1894), .CO(n1891), .S(n1892) );
  FA_X1 U1347 ( .A(n1909), .B(n1911), .CI(n1898), .CO(n1893), .S(n1894) );
  FA_X1 U1348 ( .A(n1902), .B(n1904), .CI(n1900), .CO(n1895), .S(n1896) );
  FA_X1 U1349 ( .A(n1915), .B(n1917), .CI(n1913), .CO(n1897), .S(n1898) );
  FA_X1 U1350 ( .A(n2394), .B(n2454), .CI(n2424), .CO(n1899), .S(n1900) );
  FA_X1 U1351 ( .A(n2334), .B(n2484), .CI(n2364), .CO(n1901), .S(n1902) );
  FA_X1 U1352 ( .A(n2304), .B(n2515), .CI(n2274), .CO(n1903), .S(n1904) );
  FA_X1 U1353 ( .A(n1921), .B(n1910), .CI(n1908), .CO(n1905), .S(n1906) );
  FA_X1 U1354 ( .A(n1923), .B(n1916), .CI(n1912), .CO(n1907), .S(n1908) );
  FA_X1 U1355 ( .A(n1925), .B(n1927), .CI(n1914), .CO(n1909), .S(n1910) );
  FA_X1 U1356 ( .A(n1918), .B(n2395), .CI(n1929), .CO(n1911), .S(n1912) );
  FA_X1 U1357 ( .A(n2455), .B(n2335), .CI(n2365), .CO(n1913), .S(n1914) );
  FA_X1 U1358 ( .A(n2516), .B(n2425), .CI(n2485), .CO(n1915), .S(n1916) );
  HA_X1 U1359 ( .A(n2305), .B(n2011), .CO(n1917), .S(n1918) );
  FA_X1 U1360 ( .A(n1933), .B(n1924), .CI(n1922), .CO(n1919), .S(n1920) );
  FA_X1 U1361 ( .A(n1926), .B(n1930), .CI(n1935), .CO(n1921), .S(n1922) );
  FA_X1 U1362 ( .A(n1937), .B(n1939), .CI(n1928), .CO(n1923), .S(n1924) );
  FA_X1 U1363 ( .A(n2426), .B(n2456), .CI(n1941), .CO(n1925), .S(n1926) );
  FA_X1 U1364 ( .A(n2366), .B(n2486), .CI(n2396), .CO(n1927), .S(n1928) );
  FA_X1 U1365 ( .A(n2336), .B(n2517), .CI(n2306), .CO(n1929), .S(n1930) );
  FA_X1 U1366 ( .A(n1945), .B(n1936), .CI(n1934), .CO(n1931), .S(n1932) );
  FA_X1 U1367 ( .A(n1940), .B(n1938), .CI(n1947), .CO(n1933), .S(n1934) );
  FA_X1 U1368 ( .A(n1951), .B(n1942), .CI(n1949), .CO(n1935), .S(n1936) );
  FA_X1 U1369 ( .A(n2367), .B(n2457), .CI(n2397), .CO(n1937), .S(n1938) );
  FA_X1 U1370 ( .A(n2518), .B(n2427), .CI(n2487), .CO(n1939), .S(n1940) );
  HA_X1 U1371 ( .A(n2337), .B(n2012), .CO(n1941), .S(n1942) );
  FA_X1 U1372 ( .A(n1948), .B(n1955), .CI(n1946), .CO(n1943), .S(n1944) );
  FA_X1 U1373 ( .A(n1952), .B(n1950), .CI(n1957), .CO(n1945), .S(n1946) );
  FA_X1 U1374 ( .A(n1961), .B(n2458), .CI(n1959), .CO(n1947), .S(n1948) );
  FA_X1 U1375 ( .A(n2398), .B(n2488), .CI(n2428), .CO(n1949), .S(n1950) );
  FA_X1 U1376 ( .A(n2368), .B(n2519), .CI(n2338), .CO(n1951), .S(n1952) );
  FA_X1 U1377 ( .A(n1965), .B(n1958), .CI(n1956), .CO(n1953), .S(n1954) );
  FA_X1 U1378 ( .A(n1967), .B(n1969), .CI(n1960), .CO(n1955), .S(n1956) );
  FA_X1 U1379 ( .A(n2399), .B(n2429), .CI(n1962), .CO(n1957), .S(n1958) );
  FA_X1 U1380 ( .A(n2520), .B(n2459), .CI(n2489), .CO(n1959), .S(n1960) );
  HA_X1 U1381 ( .A(n2369), .B(n2013), .CO(n1961), .S(n1962) );
  FA_X1 U1382 ( .A(n1973), .B(n1970), .CI(n1966), .CO(n1963), .S(n1964) );
  FA_X1 U1383 ( .A(n1975), .B(n1977), .CI(n1968), .CO(n1965), .S(n1966) );
  FA_X1 U1384 ( .A(n2430), .B(n2490), .CI(n2460), .CO(n1967), .S(n1968) );
  FA_X1 U1385 ( .A(n2400), .B(n2521), .CI(n2370), .CO(n1969), .S(n1970) );
  FA_X1 U1386 ( .A(n1976), .B(n1981), .CI(n1974), .CO(n1971), .S(n1972) );
  FA_X1 U1387 ( .A(n1978), .B(n2522), .CI(n1983), .CO(n1973), .S(n1974) );
  FA_X1 U1388 ( .A(n2431), .B(n2461), .CI(n2491), .CO(n1975), .S(n1976) );
  HA_X1 U1389 ( .A(n2401), .B(n2014), .CO(n1977), .S(n1978) );
  FA_X1 U1390 ( .A(n1984), .B(n1987), .CI(n1982), .CO(n1979), .S(n1980) );
  FA_X1 U1391 ( .A(n2462), .B(n2492), .CI(n1989), .CO(n1981), .S(n1982) );
  FA_X1 U1392 ( .A(n2432), .B(n2523), .CI(n2402), .CO(n1983), .S(n1984) );
  FA_X1 U1393 ( .A(n1993), .B(n1990), .CI(n1988), .CO(n1985), .S(n1986) );
  FA_X1 U1394 ( .A(n2463), .B(n2524), .CI(n2493), .CO(n1987), .S(n1988) );
  HA_X1 U1395 ( .A(n2433), .B(n2015), .CO(n1989), .S(n1990) );
  FA_X1 U1396 ( .A(n1997), .B(n2494), .CI(n1994), .CO(n1991), .S(n1992) );
  FA_X1 U1397 ( .A(n2464), .B(n2525), .CI(n2434), .CO(n1993), .S(n1994) );
  FA_X1 U1398 ( .A(n2495), .B(n2526), .CI(n1998), .CO(n1995), .S(n1996) );
  HA_X1 U1399 ( .A(n2465), .B(n2016), .CO(n1997), .S(n1998) );
  FA_X1 U1400 ( .A(n2496), .B(n2527), .CI(n2466), .CO(n1999), .S(n2000) );
  HA_X1 U1401 ( .A(n2528), .B(n2497), .CO(n2001), .S(n2002) );
  OAI22_X2 U1402 ( .A1(n440), .A2(n3139), .B1(n2563), .B2(n392), .ZN(n2003) );
  OAI22_X2 U1404 ( .A1(n440), .A2(n2533), .B1(n2532), .B2(n392), .ZN(n2020) );
  OAI22_X2 U1405 ( .A1(n440), .A2(n2534), .B1(n2533), .B2(n392), .ZN(n2021) );
  OAI22_X2 U1406 ( .A1(n440), .A2(n2535), .B1(n2534), .B2(n392), .ZN(n2022) );
  OAI22_X2 U1407 ( .A1(n440), .A2(n2536), .B1(n2535), .B2(n392), .ZN(n2023) );
  OAI22_X2 U1408 ( .A1(n440), .A2(n2537), .B1(n2536), .B2(n392), .ZN(n2024) );
  OAI22_X2 U1409 ( .A1(n440), .A2(n2538), .B1(n2537), .B2(n392), .ZN(n2025) );
  OAI22_X2 U1410 ( .A1(n440), .A2(n2539), .B1(n2538), .B2(n392), .ZN(n2026) );
  OAI22_X2 U1411 ( .A1(n440), .A2(n2540), .B1(n2539), .B2(n392), .ZN(n2027) );
  OAI22_X2 U1412 ( .A1(n439), .A2(n2541), .B1(n2540), .B2(n391), .ZN(n2028) );
  OAI22_X2 U1413 ( .A1(n439), .A2(n2542), .B1(n2541), .B2(n391), .ZN(n2029) );
  OAI22_X2 U1414 ( .A1(n439), .A2(n2543), .B1(n2542), .B2(n391), .ZN(n2030) );
  OAI22_X2 U1415 ( .A1(n439), .A2(n2544), .B1(n2543), .B2(n391), .ZN(n2031) );
  OAI22_X2 U1416 ( .A1(n439), .A2(n2545), .B1(n2544), .B2(n391), .ZN(n2032) );
  OAI22_X2 U1417 ( .A1(n439), .A2(n2546), .B1(n2545), .B2(n391), .ZN(n2033) );
  OAI22_X2 U1418 ( .A1(n439), .A2(n2547), .B1(n2546), .B2(n391), .ZN(n2034) );
  OAI22_X2 U1419 ( .A1(n439), .A2(n2548), .B1(n2547), .B2(n391), .ZN(n2035) );
  OAI22_X2 U1420 ( .A1(n439), .A2(n2549), .B1(n2548), .B2(n391), .ZN(n2036) );
  OAI22_X2 U1421 ( .A1(n439), .A2(n2550), .B1(n2549), .B2(n391), .ZN(n2037) );
  OAI22_X2 U1422 ( .A1(n439), .A2(n2551), .B1(n2550), .B2(n391), .ZN(n2038) );
  OAI22_X2 U1423 ( .A1(n438), .A2(n2552), .B1(n2551), .B2(n391), .ZN(n2039) );
  OAI22_X2 U1424 ( .A1(n438), .A2(n2553), .B1(n2552), .B2(n390), .ZN(n2040) );
  OAI22_X2 U1425 ( .A1(n438), .A2(n2554), .B1(n2553), .B2(n390), .ZN(n2041) );
  OAI22_X2 U1426 ( .A1(n438), .A2(n2555), .B1(n2554), .B2(n390), .ZN(n2042) );
  OAI22_X2 U1427 ( .A1(n438), .A2(n2556), .B1(n2555), .B2(n390), .ZN(n2043) );
  OAI22_X2 U1428 ( .A1(n438), .A2(n2557), .B1(n2556), .B2(n390), .ZN(n2044) );
  OAI22_X2 U1429 ( .A1(n438), .A2(n2558), .B1(n2557), .B2(n390), .ZN(n2045) );
  OAI22_X2 U1430 ( .A1(n438), .A2(n2559), .B1(n2558), .B2(n390), .ZN(n2046) );
  OAI22_X2 U1431 ( .A1(n438), .A2(n2560), .B1(n2559), .B2(n390), .ZN(n2047) );
  OAI22_X2 U1432 ( .A1(n438), .A2(n2561), .B1(n2560), .B2(n390), .ZN(n2048) );
  OAI22_X2 U1433 ( .A1(n438), .A2(n2562), .B1(n2561), .B2(n390), .ZN(n2049) );
  XNOR2_X2 U1434 ( .A(n3059), .B(n342), .ZN(n2531) );
  XNOR2_X2 U1435 ( .A(n3060), .B(n342), .ZN(n2532) );
  XNOR2_X2 U1436 ( .A(n3061), .B(n342), .ZN(n2533) );
  XNOR2_X2 U1437 ( .A(n3062), .B(n342), .ZN(n2534) );
  XNOR2_X2 U1438 ( .A(n3063), .B(n342), .ZN(n2535) );
  XNOR2_X2 U1439 ( .A(n3064), .B(n342), .ZN(n2536) );
  XNOR2_X2 U1440 ( .A(n3065), .B(n342), .ZN(n2537) );
  XNOR2_X2 U1441 ( .A(n3066), .B(n342), .ZN(n2538) );
  XNOR2_X2 U1442 ( .A(n3067), .B(n342), .ZN(n2539) );
  XNOR2_X2 U1443 ( .A(n3068), .B(n342), .ZN(n2540) );
  XNOR2_X2 U1444 ( .A(n3069), .B(n342), .ZN(n2541) );
  XNOR2_X2 U1445 ( .A(n3070), .B(n342), .ZN(n2542) );
  XNOR2_X2 U1446 ( .A(n3071), .B(n342), .ZN(n2543) );
  XNOR2_X2 U1447 ( .A(n3072), .B(n342), .ZN(n2544) );
  XNOR2_X2 U1448 ( .A(n3073), .B(n342), .ZN(n2545) );
  XNOR2_X2 U1449 ( .A(n3074), .B(n342), .ZN(n2546) );
  XNOR2_X2 U1450 ( .A(n3075), .B(n342), .ZN(n2547) );
  XNOR2_X2 U1451 ( .A(n3076), .B(n342), .ZN(n2548) );
  XNOR2_X2 U1452 ( .A(n3077), .B(n342), .ZN(n2549) );
  XNOR2_X2 U1453 ( .A(n3078), .B(n342), .ZN(n2550) );
  XNOR2_X2 U1454 ( .A(n3079), .B(n342), .ZN(n2551) );
  XNOR2_X2 U1455 ( .A(n3080), .B(n342), .ZN(n2552) );
  XNOR2_X2 U1456 ( .A(n3081), .B(n342), .ZN(n2553) );
  XNOR2_X2 U1457 ( .A(n3082), .B(n342), .ZN(n2554) );
  XNOR2_X2 U1458 ( .A(n3083), .B(n342), .ZN(n2555) );
  XNOR2_X2 U1459 ( .A(n3084), .B(n342), .ZN(n2556) );
  XNOR2_X2 U1460 ( .A(n3085), .B(n342), .ZN(n2557) );
  XNOR2_X2 U1461 ( .A(n3086), .B(n342), .ZN(n2558) );
  XNOR2_X2 U1462 ( .A(n3087), .B(n342), .ZN(n2559) );
  XNOR2_X2 U1463 ( .A(n3088), .B(n342), .ZN(n2560) );
  XNOR2_X2 U1464 ( .A(n3089), .B(n342), .ZN(n2561) );
  XNOR2_X2 U1465 ( .A(n441), .B(n342), .ZN(n2562) );
  OAI22_X2 U1466 ( .A1(n437), .A2(n3140), .B1(n2596), .B2(n389), .ZN(n2004) );
  OAI22_X2 U1468 ( .A1(n437), .A2(n2566), .B1(n2565), .B2(n389), .ZN(n2052) );
  OAI22_X2 U1469 ( .A1(n437), .A2(n2567), .B1(n2566), .B2(n389), .ZN(n2053) );
  OAI22_X2 U1470 ( .A1(n437), .A2(n2568), .B1(n2567), .B2(n389), .ZN(n2054) );
  OAI22_X2 U1471 ( .A1(n437), .A2(n2569), .B1(n2568), .B2(n389), .ZN(n2055) );
  OAI22_X2 U1472 ( .A1(n437), .A2(n2570), .B1(n2569), .B2(n389), .ZN(n2056) );
  OAI22_X2 U1473 ( .A1(n437), .A2(n2571), .B1(n2570), .B2(n389), .ZN(n2057) );
  OAI22_X2 U1474 ( .A1(n437), .A2(n2572), .B1(n2571), .B2(n389), .ZN(n2058) );
  OAI22_X2 U1475 ( .A1(n437), .A2(n2573), .B1(n2572), .B2(n389), .ZN(n2059) );
  OAI22_X2 U1476 ( .A1(n436), .A2(n2574), .B1(n2573), .B2(n388), .ZN(n2060) );
  OAI22_X2 U1477 ( .A1(n436), .A2(n2575), .B1(n2574), .B2(n388), .ZN(n2061) );
  OAI22_X2 U1478 ( .A1(n436), .A2(n2576), .B1(n2575), .B2(n388), .ZN(n2062) );
  OAI22_X2 U1479 ( .A1(n436), .A2(n2577), .B1(n2576), .B2(n388), .ZN(n2063) );
  OAI22_X2 U1480 ( .A1(n436), .A2(n2578), .B1(n2577), .B2(n388), .ZN(n2064) );
  OAI22_X2 U1481 ( .A1(n436), .A2(n2579), .B1(n2578), .B2(n388), .ZN(n2065) );
  OAI22_X2 U1482 ( .A1(n436), .A2(n2580), .B1(n2579), .B2(n388), .ZN(n2066) );
  OAI22_X2 U1483 ( .A1(n436), .A2(n2581), .B1(n2580), .B2(n388), .ZN(n2067) );
  OAI22_X2 U1484 ( .A1(n436), .A2(n2582), .B1(n2581), .B2(n388), .ZN(n2068) );
  OAI22_X2 U1485 ( .A1(n436), .A2(n2583), .B1(n2582), .B2(n388), .ZN(n2069) );
  OAI22_X2 U1486 ( .A1(n436), .A2(n2584), .B1(n2583), .B2(n388), .ZN(n2070) );
  OAI22_X2 U1487 ( .A1(n435), .A2(n2585), .B1(n2584), .B2(n388), .ZN(n2071) );
  OAI22_X2 U1488 ( .A1(n435), .A2(n2586), .B1(n2585), .B2(n387), .ZN(n2072) );
  OAI22_X2 U1489 ( .A1(n435), .A2(n2587), .B1(n2586), .B2(n387), .ZN(n2073) );
  OAI22_X2 U1490 ( .A1(n435), .A2(n2588), .B1(n2587), .B2(n387), .ZN(n2074) );
  OAI22_X2 U1491 ( .A1(n435), .A2(n2589), .B1(n2588), .B2(n387), .ZN(n2075) );
  OAI22_X2 U1492 ( .A1(n435), .A2(n2590), .B1(n2589), .B2(n387), .ZN(n2076) );
  OAI22_X2 U1493 ( .A1(n435), .A2(n2591), .B1(n2590), .B2(n387), .ZN(n2077) );
  OAI22_X2 U1494 ( .A1(n435), .A2(n2592), .B1(n2591), .B2(n387), .ZN(n2078) );
  OAI22_X2 U1495 ( .A1(n435), .A2(n2593), .B1(n2592), .B2(n387), .ZN(n2079) );
  OAI22_X2 U1496 ( .A1(n435), .A2(n2594), .B1(n2593), .B2(n387), .ZN(n2080) );
  OAI22_X2 U1497 ( .A1(n435), .A2(n2595), .B1(n2594), .B2(n387), .ZN(n2081) );
  XNOR2_X2 U1498 ( .A(n3059), .B(n341), .ZN(n2564) );
  XNOR2_X2 U1499 ( .A(n3060), .B(n341), .ZN(n2565) );
  XNOR2_X2 U1500 ( .A(n3061), .B(n341), .ZN(n2566) );
  XNOR2_X2 U1501 ( .A(n3062), .B(n341), .ZN(n2567) );
  XNOR2_X2 U1502 ( .A(n3063), .B(n341), .ZN(n2568) );
  XNOR2_X2 U1503 ( .A(n3064), .B(n341), .ZN(n2569) );
  XNOR2_X2 U1504 ( .A(n3065), .B(n341), .ZN(n2570) );
  XNOR2_X2 U1505 ( .A(n3066), .B(n341), .ZN(n2571) );
  XNOR2_X2 U1506 ( .A(n3067), .B(n341), .ZN(n2572) );
  XNOR2_X2 U1507 ( .A(n3068), .B(n341), .ZN(n2573) );
  XNOR2_X2 U1508 ( .A(n3069), .B(n341), .ZN(n2574) );
  XNOR2_X2 U1509 ( .A(n3070), .B(n340), .ZN(n2575) );
  XNOR2_X2 U1510 ( .A(n3071), .B(n340), .ZN(n2576) );
  XNOR2_X2 U1511 ( .A(n3072), .B(n340), .ZN(n2577) );
  XNOR2_X2 U1512 ( .A(n3073), .B(n340), .ZN(n2578) );
  XNOR2_X2 U1513 ( .A(n3074), .B(n340), .ZN(n2579) );
  XNOR2_X2 U1514 ( .A(n3075), .B(n340), .ZN(n2580) );
  XNOR2_X2 U1515 ( .A(n3076), .B(n340), .ZN(n2581) );
  XNOR2_X2 U1516 ( .A(n3077), .B(n340), .ZN(n2582) );
  XNOR2_X2 U1517 ( .A(n3078), .B(n340), .ZN(n2583) );
  XNOR2_X2 U1518 ( .A(n3079), .B(n340), .ZN(n2584) );
  XNOR2_X2 U1519 ( .A(n3080), .B(n340), .ZN(n2585) );
  XNOR2_X2 U1520 ( .A(n3081), .B(n340), .ZN(n2586) );
  XNOR2_X2 U1521 ( .A(n3082), .B(n339), .ZN(n2587) );
  XNOR2_X2 U1522 ( .A(n3083), .B(n339), .ZN(n2588) );
  XNOR2_X2 U1523 ( .A(n3084), .B(n339), .ZN(n2589) );
  XNOR2_X2 U1524 ( .A(n3085), .B(n339), .ZN(n2590) );
  XNOR2_X2 U1525 ( .A(n3086), .B(n339), .ZN(n2591) );
  XNOR2_X2 U1526 ( .A(n3087), .B(n339), .ZN(n2592) );
  XNOR2_X2 U1527 ( .A(n3088), .B(n339), .ZN(n2593) );
  XNOR2_X2 U1528 ( .A(n3089), .B(n339), .ZN(n2594) );
  XNOR2_X2 U1529 ( .A(n441), .B(n339), .ZN(n2595) );
  OAI22_X2 U1530 ( .A1(n434), .A2(n3141), .B1(n2629), .B2(n386), .ZN(n2005) );
  OAI22_X2 U1532 ( .A1(n434), .A2(n2599), .B1(n2598), .B2(n386), .ZN(n2084) );
  OAI22_X2 U1533 ( .A1(n434), .A2(n2600), .B1(n2599), .B2(n386), .ZN(n2085) );
  OAI22_X2 U1534 ( .A1(n434), .A2(n2601), .B1(n2600), .B2(n386), .ZN(n2086) );
  OAI22_X2 U1535 ( .A1(n434), .A2(n2602), .B1(n2601), .B2(n386), .ZN(n2087) );
  OAI22_X2 U1536 ( .A1(n434), .A2(n2603), .B1(n2602), .B2(n386), .ZN(n2088) );
  OAI22_X2 U1537 ( .A1(n434), .A2(n2604), .B1(n2603), .B2(n386), .ZN(n2089) );
  OAI22_X2 U1538 ( .A1(n434), .A2(n2605), .B1(n2604), .B2(n386), .ZN(n2090) );
  OAI22_X2 U1539 ( .A1(n434), .A2(n2606), .B1(n2605), .B2(n386), .ZN(n2091) );
  OAI22_X2 U1540 ( .A1(n433), .A2(n2607), .B1(n2606), .B2(n385), .ZN(n2092) );
  OAI22_X2 U1541 ( .A1(n433), .A2(n2608), .B1(n2607), .B2(n385), .ZN(n2093) );
  OAI22_X2 U1542 ( .A1(n433), .A2(n2609), .B1(n2608), .B2(n385), .ZN(n2094) );
  OAI22_X2 U1543 ( .A1(n433), .A2(n2610), .B1(n2609), .B2(n385), .ZN(n2095) );
  OAI22_X2 U1544 ( .A1(n433), .A2(n2611), .B1(n2610), .B2(n385), .ZN(n2096) );
  OAI22_X2 U1545 ( .A1(n433), .A2(n2612), .B1(n2611), .B2(n385), .ZN(n2097) );
  OAI22_X2 U1546 ( .A1(n433), .A2(n2613), .B1(n2612), .B2(n385), .ZN(n2098) );
  OAI22_X2 U1547 ( .A1(n433), .A2(n2614), .B1(n2613), .B2(n385), .ZN(n2099) );
  OAI22_X2 U1548 ( .A1(n433), .A2(n2615), .B1(n2614), .B2(n385), .ZN(n2100) );
  OAI22_X2 U1549 ( .A1(n433), .A2(n2616), .B1(n2615), .B2(n385), .ZN(n2101) );
  OAI22_X2 U1550 ( .A1(n433), .A2(n2617), .B1(n2616), .B2(n385), .ZN(n2102) );
  OAI22_X2 U1551 ( .A1(n432), .A2(n2618), .B1(n2617), .B2(n385), .ZN(n2103) );
  OAI22_X2 U1552 ( .A1(n432), .A2(n2619), .B1(n2618), .B2(n384), .ZN(n2104) );
  OAI22_X2 U1553 ( .A1(n432), .A2(n2620), .B1(n2619), .B2(n384), .ZN(n2105) );
  OAI22_X2 U1554 ( .A1(n432), .A2(n2621), .B1(n2620), .B2(n384), .ZN(n2106) );
  OAI22_X2 U1555 ( .A1(n432), .A2(n2622), .B1(n2621), .B2(n384), .ZN(n2107) );
  OAI22_X2 U1556 ( .A1(n432), .A2(n2623), .B1(n2622), .B2(n384), .ZN(n2108) );
  OAI22_X2 U1557 ( .A1(n432), .A2(n2624), .B1(n2623), .B2(n384), .ZN(n2109) );
  OAI22_X2 U1558 ( .A1(n432), .A2(n2625), .B1(n2624), .B2(n384), .ZN(n2110) );
  OAI22_X2 U1559 ( .A1(n432), .A2(n2626), .B1(n2625), .B2(n384), .ZN(n2111) );
  OAI22_X2 U1560 ( .A1(n432), .A2(n2627), .B1(n2626), .B2(n384), .ZN(n2112) );
  OAI22_X2 U1561 ( .A1(n432), .A2(n2628), .B1(n2627), .B2(n384), .ZN(n2113) );
  XNOR2_X2 U1562 ( .A(n3059), .B(n338), .ZN(n2597) );
  XNOR2_X2 U1563 ( .A(n3060), .B(n338), .ZN(n2598) );
  XNOR2_X2 U1564 ( .A(n3061), .B(n338), .ZN(n2599) );
  XNOR2_X2 U1565 ( .A(n3062), .B(n338), .ZN(n2600) );
  XNOR2_X2 U1566 ( .A(n3063), .B(n338), .ZN(n2601) );
  XNOR2_X2 U1567 ( .A(n3064), .B(n338), .ZN(n2602) );
  XNOR2_X2 U1568 ( .A(n3065), .B(n338), .ZN(n2603) );
  XNOR2_X2 U1569 ( .A(n3066), .B(n338), .ZN(n2604) );
  XNOR2_X2 U1570 ( .A(n3067), .B(n338), .ZN(n2605) );
  XNOR2_X2 U1571 ( .A(n3068), .B(n338), .ZN(n2606) );
  XNOR2_X2 U1572 ( .A(n3069), .B(n338), .ZN(n2607) );
  XNOR2_X2 U1573 ( .A(n3070), .B(n337), .ZN(n2608) );
  XNOR2_X2 U1574 ( .A(n3071), .B(n337), .ZN(n2609) );
  XNOR2_X2 U1575 ( .A(n3072), .B(n337), .ZN(n2610) );
  XNOR2_X2 U1576 ( .A(n3073), .B(n337), .ZN(n2611) );
  XNOR2_X2 U1577 ( .A(n3074), .B(n337), .ZN(n2612) );
  XNOR2_X2 U1578 ( .A(n3075), .B(n337), .ZN(n2613) );
  XNOR2_X2 U1579 ( .A(n3076), .B(n337), .ZN(n2614) );
  XNOR2_X2 U1580 ( .A(n3077), .B(n337), .ZN(n2615) );
  XNOR2_X2 U1581 ( .A(n3078), .B(n337), .ZN(n2616) );
  XNOR2_X2 U1582 ( .A(n3079), .B(n337), .ZN(n2617) );
  XNOR2_X2 U1583 ( .A(n3080), .B(n337), .ZN(n2618) );
  XNOR2_X2 U1584 ( .A(n3081), .B(n337), .ZN(n2619) );
  XNOR2_X2 U1585 ( .A(n3082), .B(n336), .ZN(n2620) );
  XNOR2_X2 U1586 ( .A(n3083), .B(n336), .ZN(n2621) );
  XNOR2_X2 U1587 ( .A(n3084), .B(n336), .ZN(n2622) );
  XNOR2_X2 U1588 ( .A(n3085), .B(n336), .ZN(n2623) );
  XNOR2_X2 U1589 ( .A(n3086), .B(n336), .ZN(n2624) );
  XNOR2_X2 U1590 ( .A(n3087), .B(n336), .ZN(n2625) );
  XNOR2_X2 U1591 ( .A(n3088), .B(n336), .ZN(n2626) );
  XNOR2_X2 U1592 ( .A(n3089), .B(n336), .ZN(n2627) );
  XNOR2_X2 U1593 ( .A(n441), .B(n336), .ZN(n2628) );
  OAI22_X2 U1594 ( .A1(n431), .A2(n3142), .B1(n2662), .B2(n383), .ZN(n2006) );
  OAI22_X2 U1596 ( .A1(n431), .A2(n2632), .B1(n2631), .B2(n383), .ZN(n2116) );
  OAI22_X2 U1597 ( .A1(n431), .A2(n2633), .B1(n2632), .B2(n383), .ZN(n2117) );
  OAI22_X2 U1598 ( .A1(n431), .A2(n2634), .B1(n2633), .B2(n383), .ZN(n2118) );
  OAI22_X2 U1599 ( .A1(n431), .A2(n2635), .B1(n2634), .B2(n383), .ZN(n2119) );
  OAI22_X2 U1600 ( .A1(n431), .A2(n2636), .B1(n2635), .B2(n383), .ZN(n2120) );
  OAI22_X2 U1601 ( .A1(n431), .A2(n2637), .B1(n2636), .B2(n383), .ZN(n2121) );
  OAI22_X2 U1602 ( .A1(n431), .A2(n2638), .B1(n2637), .B2(n383), .ZN(n2122) );
  OAI22_X2 U1603 ( .A1(n431), .A2(n2639), .B1(n2638), .B2(n383), .ZN(n2123) );
  OAI22_X2 U1604 ( .A1(n430), .A2(n2640), .B1(n2639), .B2(n382), .ZN(n2124) );
  OAI22_X2 U1605 ( .A1(n430), .A2(n2641), .B1(n2640), .B2(n382), .ZN(n2125) );
  OAI22_X2 U1606 ( .A1(n430), .A2(n2642), .B1(n2641), .B2(n382), .ZN(n2126) );
  OAI22_X2 U1607 ( .A1(n430), .A2(n2643), .B1(n2642), .B2(n382), .ZN(n2127) );
  OAI22_X2 U1608 ( .A1(n430), .A2(n2644), .B1(n2643), .B2(n382), .ZN(n2128) );
  OAI22_X2 U1609 ( .A1(n430), .A2(n2645), .B1(n2644), .B2(n382), .ZN(n2129) );
  OAI22_X2 U1610 ( .A1(n430), .A2(n2646), .B1(n2645), .B2(n382), .ZN(n2130) );
  OAI22_X2 U1611 ( .A1(n430), .A2(n2647), .B1(n2646), .B2(n382), .ZN(n2131) );
  OAI22_X2 U1612 ( .A1(n430), .A2(n2648), .B1(n2647), .B2(n382), .ZN(n2132) );
  OAI22_X2 U1613 ( .A1(n430), .A2(n2649), .B1(n2648), .B2(n382), .ZN(n2133) );
  OAI22_X2 U1614 ( .A1(n430), .A2(n2650), .B1(n2649), .B2(n382), .ZN(n2134) );
  OAI22_X2 U1615 ( .A1(n429), .A2(n2651), .B1(n2650), .B2(n382), .ZN(n2135) );
  OAI22_X2 U1616 ( .A1(n429), .A2(n2652), .B1(n2651), .B2(n381), .ZN(n2136) );
  OAI22_X2 U1617 ( .A1(n429), .A2(n2653), .B1(n2652), .B2(n381), .ZN(n2137) );
  OAI22_X2 U1618 ( .A1(n429), .A2(n2654), .B1(n2653), .B2(n381), .ZN(n2138) );
  OAI22_X2 U1619 ( .A1(n429), .A2(n2655), .B1(n2654), .B2(n381), .ZN(n2139) );
  OAI22_X2 U1620 ( .A1(n429), .A2(n2656), .B1(n2655), .B2(n381), .ZN(n2140) );
  OAI22_X2 U1621 ( .A1(n429), .A2(n2657), .B1(n2656), .B2(n381), .ZN(n2141) );
  OAI22_X2 U1622 ( .A1(n429), .A2(n2658), .B1(n2657), .B2(n381), .ZN(n2142) );
  OAI22_X2 U1623 ( .A1(n429), .A2(n2659), .B1(n2658), .B2(n381), .ZN(n2143) );
  OAI22_X2 U1624 ( .A1(n429), .A2(n2660), .B1(n2659), .B2(n381), .ZN(n2144) );
  OAI22_X2 U1625 ( .A1(n429), .A2(n2661), .B1(n2660), .B2(n381), .ZN(n2145) );
  XNOR2_X2 U1626 ( .A(n3059), .B(n335), .ZN(n2630) );
  XNOR2_X2 U1627 ( .A(n3060), .B(n335), .ZN(n2631) );
  XNOR2_X2 U1628 ( .A(n3061), .B(n335), .ZN(n2632) );
  XNOR2_X2 U1629 ( .A(n3062), .B(n335), .ZN(n2633) );
  XNOR2_X2 U1630 ( .A(n3063), .B(n335), .ZN(n2634) );
  XNOR2_X2 U1631 ( .A(n3064), .B(n335), .ZN(n2635) );
  XNOR2_X2 U1632 ( .A(n3065), .B(n335), .ZN(n2636) );
  XNOR2_X2 U1633 ( .A(n3066), .B(n335), .ZN(n2637) );
  XNOR2_X2 U1634 ( .A(n3067), .B(n335), .ZN(n2638) );
  XNOR2_X2 U1635 ( .A(n3068), .B(n335), .ZN(n2639) );
  XNOR2_X2 U1636 ( .A(n3069), .B(n335), .ZN(n2640) );
  XNOR2_X2 U1637 ( .A(n3070), .B(n334), .ZN(n2641) );
  XNOR2_X2 U1638 ( .A(n3071), .B(n334), .ZN(n2642) );
  XNOR2_X2 U1639 ( .A(n3072), .B(n334), .ZN(n2643) );
  XNOR2_X2 U1640 ( .A(n3073), .B(n334), .ZN(n2644) );
  XNOR2_X2 U1641 ( .A(n3074), .B(n334), .ZN(n2645) );
  XNOR2_X2 U1642 ( .A(n3075), .B(n334), .ZN(n2646) );
  XNOR2_X2 U1643 ( .A(n3076), .B(n334), .ZN(n2647) );
  XNOR2_X2 U1644 ( .A(n3077), .B(n334), .ZN(n2648) );
  XNOR2_X2 U1645 ( .A(n3078), .B(n334), .ZN(n2649) );
  XNOR2_X2 U1646 ( .A(n3079), .B(n334), .ZN(n2650) );
  XNOR2_X2 U1647 ( .A(n3080), .B(n334), .ZN(n2651) );
  XNOR2_X2 U1648 ( .A(n3081), .B(n334), .ZN(n2652) );
  XNOR2_X2 U1649 ( .A(n3082), .B(n333), .ZN(n2653) );
  XNOR2_X2 U1650 ( .A(n3083), .B(n333), .ZN(n2654) );
  XNOR2_X2 U1651 ( .A(n3084), .B(n333), .ZN(n2655) );
  XNOR2_X2 U1652 ( .A(n3085), .B(n333), .ZN(n2656) );
  XNOR2_X2 U1653 ( .A(n3086), .B(n333), .ZN(n2657) );
  XNOR2_X2 U1654 ( .A(n3087), .B(n333), .ZN(n2658) );
  XNOR2_X2 U1655 ( .A(n3088), .B(n333), .ZN(n2659) );
  XNOR2_X2 U1656 ( .A(n3089), .B(n333), .ZN(n2660) );
  XNOR2_X2 U1657 ( .A(n441), .B(n333), .ZN(n2661) );
  OAI22_X2 U1658 ( .A1(n428), .A2(n3143), .B1(n2695), .B2(n380), .ZN(n2007) );
  OAI22_X2 U1660 ( .A1(n428), .A2(n2665), .B1(n2664), .B2(n380), .ZN(n2148) );
  OAI22_X2 U1661 ( .A1(n428), .A2(n2666), .B1(n2665), .B2(n380), .ZN(n2149) );
  OAI22_X2 U1662 ( .A1(n428), .A2(n2667), .B1(n2666), .B2(n380), .ZN(n2150) );
  OAI22_X2 U1663 ( .A1(n428), .A2(n2668), .B1(n2667), .B2(n380), .ZN(n2151) );
  OAI22_X2 U1664 ( .A1(n428), .A2(n2669), .B1(n2668), .B2(n380), .ZN(n2152) );
  OAI22_X2 U1665 ( .A1(n428), .A2(n2670), .B1(n2669), .B2(n380), .ZN(n2153) );
  OAI22_X2 U1666 ( .A1(n428), .A2(n2671), .B1(n2670), .B2(n380), .ZN(n2154) );
  OAI22_X2 U1667 ( .A1(n428), .A2(n2672), .B1(n2671), .B2(n380), .ZN(n2155) );
  OAI22_X2 U1668 ( .A1(n427), .A2(n2673), .B1(n2672), .B2(n379), .ZN(n2156) );
  OAI22_X2 U1669 ( .A1(n427), .A2(n2674), .B1(n2673), .B2(n379), .ZN(n2157) );
  OAI22_X2 U1670 ( .A1(n427), .A2(n2675), .B1(n2674), .B2(n379), .ZN(n2158) );
  OAI22_X2 U1671 ( .A1(n427), .A2(n2676), .B1(n2675), .B2(n379), .ZN(n2159) );
  OAI22_X2 U1672 ( .A1(n427), .A2(n2677), .B1(n2676), .B2(n379), .ZN(n2160) );
  OAI22_X2 U1673 ( .A1(n427), .A2(n2678), .B1(n2677), .B2(n379), .ZN(n2161) );
  OAI22_X2 U1674 ( .A1(n427), .A2(n2679), .B1(n2678), .B2(n379), .ZN(n2162) );
  OAI22_X2 U1675 ( .A1(n427), .A2(n2680), .B1(n2679), .B2(n379), .ZN(n2163) );
  OAI22_X2 U1676 ( .A1(n427), .A2(n2681), .B1(n2680), .B2(n379), .ZN(n2164) );
  OAI22_X2 U1677 ( .A1(n427), .A2(n2682), .B1(n2681), .B2(n379), .ZN(n2165) );
  OAI22_X2 U1678 ( .A1(n427), .A2(n2683), .B1(n2682), .B2(n379), .ZN(n2166) );
  OAI22_X2 U1679 ( .A1(n426), .A2(n2684), .B1(n2683), .B2(n379), .ZN(n2167) );
  OAI22_X2 U1680 ( .A1(n426), .A2(n2685), .B1(n2684), .B2(n378), .ZN(n2168) );
  OAI22_X2 U1681 ( .A1(n426), .A2(n2686), .B1(n2685), .B2(n378), .ZN(n2169) );
  OAI22_X2 U1682 ( .A1(n426), .A2(n2687), .B1(n2686), .B2(n378), .ZN(n2170) );
  OAI22_X2 U1683 ( .A1(n426), .A2(n2688), .B1(n2687), .B2(n378), .ZN(n2171) );
  OAI22_X2 U1684 ( .A1(n426), .A2(n2689), .B1(n2688), .B2(n378), .ZN(n2172) );
  OAI22_X2 U1685 ( .A1(n426), .A2(n2690), .B1(n2689), .B2(n378), .ZN(n2173) );
  OAI22_X2 U1686 ( .A1(n426), .A2(n2691), .B1(n2690), .B2(n378), .ZN(n2174) );
  OAI22_X2 U1687 ( .A1(n426), .A2(n2692), .B1(n2691), .B2(n378), .ZN(n2175) );
  OAI22_X2 U1688 ( .A1(n426), .A2(n2693), .B1(n2692), .B2(n378), .ZN(n2176) );
  OAI22_X2 U1689 ( .A1(n426), .A2(n2694), .B1(n2693), .B2(n378), .ZN(n2177) );
  XNOR2_X2 U1690 ( .A(n3059), .B(n332), .ZN(n2663) );
  XNOR2_X2 U1691 ( .A(n3060), .B(n332), .ZN(n2664) );
  XNOR2_X2 U1692 ( .A(n3061), .B(n332), .ZN(n2665) );
  XNOR2_X2 U1693 ( .A(n3062), .B(n332), .ZN(n2666) );
  XNOR2_X2 U1694 ( .A(n3063), .B(n332), .ZN(n2667) );
  XNOR2_X2 U1695 ( .A(n3064), .B(n332), .ZN(n2668) );
  XNOR2_X2 U1696 ( .A(n3065), .B(n332), .ZN(n2669) );
  XNOR2_X2 U1697 ( .A(n3066), .B(n332), .ZN(n2670) );
  XNOR2_X2 U1698 ( .A(n3067), .B(n332), .ZN(n2671) );
  XNOR2_X2 U1699 ( .A(n3068), .B(n332), .ZN(n2672) );
  XNOR2_X2 U1700 ( .A(n3069), .B(n332), .ZN(n2673) );
  XNOR2_X2 U1701 ( .A(n3070), .B(n331), .ZN(n2674) );
  XNOR2_X2 U1702 ( .A(n3071), .B(n331), .ZN(n2675) );
  XNOR2_X2 U1703 ( .A(n3072), .B(n331), .ZN(n2676) );
  XNOR2_X2 U1704 ( .A(n3073), .B(n331), .ZN(n2677) );
  XNOR2_X2 U1705 ( .A(n3074), .B(n331), .ZN(n2678) );
  XNOR2_X2 U1706 ( .A(n3075), .B(n331), .ZN(n2679) );
  XNOR2_X2 U1707 ( .A(n3076), .B(n331), .ZN(n2680) );
  XNOR2_X2 U1708 ( .A(n3077), .B(n331), .ZN(n2681) );
  XNOR2_X2 U1709 ( .A(n3078), .B(n331), .ZN(n2682) );
  XNOR2_X2 U1710 ( .A(n3079), .B(n331), .ZN(n2683) );
  XNOR2_X2 U1711 ( .A(n3080), .B(n331), .ZN(n2684) );
  XNOR2_X2 U1712 ( .A(n3081), .B(n331), .ZN(n2685) );
  XNOR2_X2 U1713 ( .A(n3082), .B(n330), .ZN(n2686) );
  XNOR2_X2 U1714 ( .A(n3083), .B(n330), .ZN(n2687) );
  XNOR2_X2 U1715 ( .A(n3084), .B(n330), .ZN(n2688) );
  XNOR2_X2 U1716 ( .A(n3085), .B(n330), .ZN(n2689) );
  XNOR2_X2 U1717 ( .A(n3086), .B(n330), .ZN(n2690) );
  XNOR2_X2 U1718 ( .A(n3087), .B(n330), .ZN(n2691) );
  XNOR2_X2 U1719 ( .A(n3088), .B(n330), .ZN(n2692) );
  XNOR2_X2 U1720 ( .A(n3089), .B(n330), .ZN(n2693) );
  XNOR2_X2 U1721 ( .A(n441), .B(n330), .ZN(n2694) );
  OAI22_X2 U1722 ( .A1(n425), .A2(n3144), .B1(n2728), .B2(n377), .ZN(n2008) );
  OAI22_X2 U1724 ( .A1(n425), .A2(n2698), .B1(n2697), .B2(n377), .ZN(n2180) );
  OAI22_X2 U1725 ( .A1(n425), .A2(n2699), .B1(n2698), .B2(n377), .ZN(n2181) );
  OAI22_X2 U1726 ( .A1(n425), .A2(n2700), .B1(n2699), .B2(n377), .ZN(n2182) );
  OAI22_X2 U1727 ( .A1(n425), .A2(n2701), .B1(n2700), .B2(n377), .ZN(n2183) );
  OAI22_X2 U1728 ( .A1(n425), .A2(n2702), .B1(n2701), .B2(n377), .ZN(n2184) );
  OAI22_X2 U1729 ( .A1(n425), .A2(n2703), .B1(n2702), .B2(n377), .ZN(n2185) );
  OAI22_X2 U1730 ( .A1(n425), .A2(n2704), .B1(n2703), .B2(n377), .ZN(n2186) );
  OAI22_X2 U1731 ( .A1(n425), .A2(n2705), .B1(n2704), .B2(n377), .ZN(n2187) );
  OAI22_X2 U1732 ( .A1(n424), .A2(n2706), .B1(n2705), .B2(n376), .ZN(n2188) );
  OAI22_X2 U1733 ( .A1(n424), .A2(n2707), .B1(n2706), .B2(n376), .ZN(n2189) );
  OAI22_X2 U1734 ( .A1(n424), .A2(n2708), .B1(n2707), .B2(n376), .ZN(n2190) );
  OAI22_X2 U1735 ( .A1(n424), .A2(n2709), .B1(n2708), .B2(n376), .ZN(n2191) );
  OAI22_X2 U1736 ( .A1(n424), .A2(n2710), .B1(n2709), .B2(n376), .ZN(n2192) );
  OAI22_X2 U1737 ( .A1(n424), .A2(n2711), .B1(n2710), .B2(n376), .ZN(n2193) );
  OAI22_X2 U1738 ( .A1(n424), .A2(n2712), .B1(n2711), .B2(n376), .ZN(n2194) );
  OAI22_X2 U1739 ( .A1(n424), .A2(n2713), .B1(n2712), .B2(n376), .ZN(n2195) );
  OAI22_X2 U1740 ( .A1(n424), .A2(n2714), .B1(n2713), .B2(n376), .ZN(n2196) );
  OAI22_X2 U1741 ( .A1(n424), .A2(n2715), .B1(n2714), .B2(n376), .ZN(n2197) );
  OAI22_X2 U1742 ( .A1(n424), .A2(n2716), .B1(n2715), .B2(n376), .ZN(n2198) );
  OAI22_X2 U1743 ( .A1(n423), .A2(n2717), .B1(n2716), .B2(n376), .ZN(n2199) );
  OAI22_X2 U1744 ( .A1(n423), .A2(n2718), .B1(n2717), .B2(n375), .ZN(n2200) );
  OAI22_X2 U1745 ( .A1(n423), .A2(n2719), .B1(n2718), .B2(n375), .ZN(n2201) );
  OAI22_X2 U1746 ( .A1(n423), .A2(n2720), .B1(n2719), .B2(n375), .ZN(n2202) );
  OAI22_X2 U1747 ( .A1(n423), .A2(n2721), .B1(n2720), .B2(n375), .ZN(n2203) );
  OAI22_X2 U1748 ( .A1(n423), .A2(n2722), .B1(n2721), .B2(n375), .ZN(n2204) );
  OAI22_X2 U1749 ( .A1(n423), .A2(n2723), .B1(n2722), .B2(n375), .ZN(n2205) );
  OAI22_X2 U1750 ( .A1(n423), .A2(n2724), .B1(n2723), .B2(n375), .ZN(n2206) );
  OAI22_X2 U1751 ( .A1(n423), .A2(n2725), .B1(n2724), .B2(n375), .ZN(n2207) );
  OAI22_X2 U1752 ( .A1(n423), .A2(n2726), .B1(n2725), .B2(n375), .ZN(n2208) );
  OAI22_X2 U1753 ( .A1(n423), .A2(n2727), .B1(n2726), .B2(n375), .ZN(n2209) );
  XNOR2_X2 U1754 ( .A(n3059), .B(n329), .ZN(n2696) );
  XNOR2_X2 U1755 ( .A(n3060), .B(n329), .ZN(n2697) );
  XNOR2_X2 U1756 ( .A(n3061), .B(n329), .ZN(n2698) );
  XNOR2_X2 U1757 ( .A(n3062), .B(n329), .ZN(n2699) );
  XNOR2_X2 U1758 ( .A(n3063), .B(n329), .ZN(n2700) );
  XNOR2_X2 U1759 ( .A(n3064), .B(n329), .ZN(n2701) );
  XNOR2_X2 U1760 ( .A(n3065), .B(n329), .ZN(n2702) );
  XNOR2_X2 U1761 ( .A(n3066), .B(n329), .ZN(n2703) );
  XNOR2_X2 U1762 ( .A(n3067), .B(n329), .ZN(n2704) );
  XNOR2_X2 U1763 ( .A(n3068), .B(n329), .ZN(n2705) );
  XNOR2_X2 U1764 ( .A(n3069), .B(n329), .ZN(n2706) );
  XNOR2_X2 U1765 ( .A(n3070), .B(n328), .ZN(n2707) );
  XNOR2_X2 U1766 ( .A(n3071), .B(n328), .ZN(n2708) );
  XNOR2_X2 U1767 ( .A(n3072), .B(n328), .ZN(n2709) );
  XNOR2_X2 U1768 ( .A(n3073), .B(n328), .ZN(n2710) );
  XNOR2_X2 U1769 ( .A(n3074), .B(n328), .ZN(n2711) );
  XNOR2_X2 U1770 ( .A(n3075), .B(n328), .ZN(n2712) );
  XNOR2_X2 U1771 ( .A(n3076), .B(n328), .ZN(n2713) );
  XNOR2_X2 U1772 ( .A(n3077), .B(n328), .ZN(n2714) );
  XNOR2_X2 U1773 ( .A(n3078), .B(n328), .ZN(n2715) );
  XNOR2_X2 U1774 ( .A(n3079), .B(n328), .ZN(n2716) );
  XNOR2_X2 U1775 ( .A(n3080), .B(n328), .ZN(n2717) );
  XNOR2_X2 U1776 ( .A(n3081), .B(n328), .ZN(n2718) );
  XNOR2_X2 U1777 ( .A(n3082), .B(n327), .ZN(n2719) );
  XNOR2_X2 U1778 ( .A(n3083), .B(n327), .ZN(n2720) );
  XNOR2_X2 U1779 ( .A(n3084), .B(n327), .ZN(n2721) );
  XNOR2_X2 U1780 ( .A(n3085), .B(n327), .ZN(n2722) );
  XNOR2_X2 U1781 ( .A(n3086), .B(n327), .ZN(n2723) );
  XNOR2_X2 U1782 ( .A(n3087), .B(n327), .ZN(n2724) );
  XNOR2_X2 U1783 ( .A(n3088), .B(n327), .ZN(n2725) );
  XNOR2_X2 U1784 ( .A(n3089), .B(n327), .ZN(n2726) );
  XNOR2_X2 U1785 ( .A(n441), .B(n327), .ZN(n2727) );
  OAI22_X2 U1786 ( .A1(n422), .A2(n3145), .B1(n2761), .B2(n374), .ZN(n2009) );
  OAI22_X2 U1788 ( .A1(n422), .A2(n2731), .B1(n2730), .B2(n374), .ZN(n2212) );
  OAI22_X2 U1789 ( .A1(n422), .A2(n2732), .B1(n2731), .B2(n374), .ZN(n2213) );
  OAI22_X2 U1790 ( .A1(n422), .A2(n2733), .B1(n2732), .B2(n374), .ZN(n2214) );
  OAI22_X2 U1791 ( .A1(n422), .A2(n2734), .B1(n2733), .B2(n374), .ZN(n2215) );
  OAI22_X2 U1792 ( .A1(n422), .A2(n2735), .B1(n2734), .B2(n374), .ZN(n2216) );
  OAI22_X2 U1793 ( .A1(n422), .A2(n2736), .B1(n2735), .B2(n374), .ZN(n2217) );
  OAI22_X2 U1794 ( .A1(n422), .A2(n2737), .B1(n2736), .B2(n374), .ZN(n2218) );
  OAI22_X2 U1795 ( .A1(n422), .A2(n2738), .B1(n2737), .B2(n374), .ZN(n2219) );
  OAI22_X2 U1796 ( .A1(n421), .A2(n2739), .B1(n2738), .B2(n373), .ZN(n2220) );
  OAI22_X2 U1797 ( .A1(n421), .A2(n2740), .B1(n2739), .B2(n373), .ZN(n2221) );
  OAI22_X2 U1798 ( .A1(n421), .A2(n2741), .B1(n2740), .B2(n373), .ZN(n2222) );
  OAI22_X2 U1799 ( .A1(n421), .A2(n2742), .B1(n2741), .B2(n373), .ZN(n2223) );
  OAI22_X2 U1800 ( .A1(n421), .A2(n2743), .B1(n2742), .B2(n373), .ZN(n2224) );
  OAI22_X2 U1801 ( .A1(n421), .A2(n2744), .B1(n2743), .B2(n373), .ZN(n2225) );
  OAI22_X2 U1802 ( .A1(n421), .A2(n2745), .B1(n2744), .B2(n373), .ZN(n2226) );
  OAI22_X2 U1803 ( .A1(n421), .A2(n2746), .B1(n2745), .B2(n373), .ZN(n2227) );
  OAI22_X2 U1804 ( .A1(n421), .A2(n2747), .B1(n2746), .B2(n373), .ZN(n2228) );
  OAI22_X2 U1805 ( .A1(n421), .A2(n2748), .B1(n2747), .B2(n373), .ZN(n2229) );
  OAI22_X2 U1806 ( .A1(n421), .A2(n2749), .B1(n2748), .B2(n373), .ZN(n2230) );
  OAI22_X2 U1807 ( .A1(n420), .A2(n2750), .B1(n2749), .B2(n373), .ZN(n2231) );
  OAI22_X2 U1808 ( .A1(n420), .A2(n2751), .B1(n2750), .B2(n372), .ZN(n2232) );
  OAI22_X2 U1809 ( .A1(n420), .A2(n2752), .B1(n2751), .B2(n372), .ZN(n2233) );
  OAI22_X2 U1810 ( .A1(n420), .A2(n2753), .B1(n2752), .B2(n372), .ZN(n2234) );
  OAI22_X2 U1811 ( .A1(n420), .A2(n2754), .B1(n2753), .B2(n372), .ZN(n2235) );
  OAI22_X2 U1812 ( .A1(n420), .A2(n2755), .B1(n2754), .B2(n372), .ZN(n2236) );
  OAI22_X2 U1813 ( .A1(n420), .A2(n2756), .B1(n2755), .B2(n372), .ZN(n2237) );
  OAI22_X2 U1814 ( .A1(n420), .A2(n2757), .B1(n2756), .B2(n372), .ZN(n2238) );
  OAI22_X2 U1815 ( .A1(n420), .A2(n2758), .B1(n2757), .B2(n372), .ZN(n2239) );
  OAI22_X2 U1816 ( .A1(n420), .A2(n2759), .B1(n2758), .B2(n372), .ZN(n2240) );
  OAI22_X2 U1817 ( .A1(n420), .A2(n2760), .B1(n2759), .B2(n372), .ZN(n2241) );
  XNOR2_X2 U1818 ( .A(n3059), .B(n326), .ZN(n2729) );
  XNOR2_X2 U1819 ( .A(n3060), .B(n326), .ZN(n2730) );
  XNOR2_X2 U1820 ( .A(n3061), .B(n326), .ZN(n2731) );
  XNOR2_X2 U1821 ( .A(n3062), .B(n326), .ZN(n2732) );
  XNOR2_X2 U1822 ( .A(n3063), .B(n326), .ZN(n2733) );
  XNOR2_X2 U1823 ( .A(n3064), .B(n326), .ZN(n2734) );
  XNOR2_X2 U1824 ( .A(n3065), .B(n326), .ZN(n2735) );
  XNOR2_X2 U1825 ( .A(n3066), .B(n326), .ZN(n2736) );
  XNOR2_X2 U1826 ( .A(n3067), .B(n326), .ZN(n2737) );
  XNOR2_X2 U1827 ( .A(n3068), .B(n326), .ZN(n2738) );
  XNOR2_X2 U1828 ( .A(n3069), .B(n326), .ZN(n2739) );
  XNOR2_X2 U1829 ( .A(n3070), .B(n325), .ZN(n2740) );
  XNOR2_X2 U1830 ( .A(n3071), .B(n325), .ZN(n2741) );
  XNOR2_X2 U1831 ( .A(n3072), .B(n325), .ZN(n2742) );
  XNOR2_X2 U1832 ( .A(n3073), .B(n325), .ZN(n2743) );
  XNOR2_X2 U1833 ( .A(n3074), .B(n325), .ZN(n2744) );
  XNOR2_X2 U1834 ( .A(n3075), .B(n325), .ZN(n2745) );
  XNOR2_X2 U1835 ( .A(n3076), .B(n325), .ZN(n2746) );
  XNOR2_X2 U1836 ( .A(n3077), .B(n325), .ZN(n2747) );
  XNOR2_X2 U1837 ( .A(n3078), .B(n325), .ZN(n2748) );
  XNOR2_X2 U1838 ( .A(n3079), .B(n325), .ZN(n2749) );
  XNOR2_X2 U1839 ( .A(n3080), .B(n325), .ZN(n2750) );
  XNOR2_X2 U1840 ( .A(n3081), .B(n325), .ZN(n2751) );
  XNOR2_X2 U1841 ( .A(n3082), .B(n324), .ZN(n2752) );
  XNOR2_X2 U1842 ( .A(n3083), .B(n324), .ZN(n2753) );
  XNOR2_X2 U1843 ( .A(n3084), .B(n324), .ZN(n2754) );
  XNOR2_X2 U1844 ( .A(n3085), .B(n324), .ZN(n2755) );
  XNOR2_X2 U1845 ( .A(n3086), .B(n324), .ZN(n2756) );
  XNOR2_X2 U1846 ( .A(n3087), .B(n324), .ZN(n2757) );
  XNOR2_X2 U1847 ( .A(n3088), .B(n324), .ZN(n2758) );
  XNOR2_X2 U1848 ( .A(n3089), .B(n324), .ZN(n2759) );
  XNOR2_X2 U1849 ( .A(n441), .B(n324), .ZN(n2760) );
  OAI22_X2 U1850 ( .A1(n419), .A2(n3146), .B1(n2794), .B2(n371), .ZN(n2010) );
  OAI22_X2 U1852 ( .A1(n419), .A2(n2764), .B1(n2763), .B2(n371), .ZN(n2244) );
  OAI22_X2 U1853 ( .A1(n419), .A2(n2765), .B1(n2764), .B2(n371), .ZN(n2245) );
  OAI22_X2 U1854 ( .A1(n419), .A2(n2766), .B1(n2765), .B2(n371), .ZN(n2246) );
  OAI22_X2 U1855 ( .A1(n419), .A2(n2767), .B1(n2766), .B2(n371), .ZN(n2247) );
  OAI22_X2 U1856 ( .A1(n419), .A2(n2768), .B1(n2767), .B2(n371), .ZN(n2248) );
  OAI22_X2 U1857 ( .A1(n419), .A2(n2769), .B1(n2768), .B2(n371), .ZN(n2249) );
  OAI22_X2 U1858 ( .A1(n419), .A2(n2770), .B1(n2769), .B2(n371), .ZN(n2250) );
  OAI22_X2 U1859 ( .A1(n419), .A2(n2771), .B1(n2770), .B2(n371), .ZN(n2251) );
  OAI22_X2 U1860 ( .A1(n418), .A2(n2772), .B1(n2771), .B2(n370), .ZN(n2252) );
  OAI22_X2 U1861 ( .A1(n418), .A2(n2773), .B1(n2772), .B2(n370), .ZN(n2253) );
  OAI22_X2 U1862 ( .A1(n418), .A2(n2774), .B1(n2773), .B2(n370), .ZN(n2254) );
  OAI22_X2 U1863 ( .A1(n418), .A2(n2775), .B1(n2774), .B2(n370), .ZN(n2255) );
  OAI22_X2 U1864 ( .A1(n418), .A2(n2776), .B1(n2775), .B2(n370), .ZN(n2256) );
  OAI22_X2 U1865 ( .A1(n418), .A2(n2777), .B1(n2776), .B2(n370), .ZN(n2257) );
  OAI22_X2 U1866 ( .A1(n418), .A2(n2778), .B1(n2777), .B2(n370), .ZN(n2258) );
  OAI22_X2 U1867 ( .A1(n418), .A2(n2779), .B1(n2778), .B2(n370), .ZN(n2259) );
  OAI22_X2 U1868 ( .A1(n418), .A2(n2780), .B1(n2779), .B2(n370), .ZN(n2260) );
  OAI22_X2 U1869 ( .A1(n418), .A2(n2781), .B1(n2780), .B2(n370), .ZN(n2261) );
  OAI22_X2 U1870 ( .A1(n418), .A2(n2782), .B1(n2781), .B2(n370), .ZN(n2262) );
  OAI22_X2 U1871 ( .A1(n417), .A2(n2783), .B1(n2782), .B2(n370), .ZN(n2263) );
  OAI22_X2 U1872 ( .A1(n417), .A2(n2784), .B1(n2783), .B2(n369), .ZN(n2264) );
  OAI22_X2 U1873 ( .A1(n417), .A2(n2785), .B1(n2784), .B2(n369), .ZN(n2265) );
  OAI22_X2 U1874 ( .A1(n417), .A2(n2786), .B1(n2785), .B2(n369), .ZN(n2266) );
  OAI22_X2 U1875 ( .A1(n417), .A2(n2787), .B1(n2786), .B2(n369), .ZN(n2267) );
  OAI22_X2 U1876 ( .A1(n417), .A2(n2788), .B1(n2787), .B2(n369), .ZN(n2268) );
  OAI22_X2 U1877 ( .A1(n417), .A2(n2789), .B1(n2788), .B2(n369), .ZN(n2269) );
  OAI22_X2 U1878 ( .A1(n417), .A2(n2790), .B1(n2789), .B2(n369), .ZN(n2270) );
  OAI22_X2 U1879 ( .A1(n417), .A2(n2791), .B1(n2790), .B2(n369), .ZN(n2271) );
  OAI22_X2 U1880 ( .A1(n417), .A2(n2792), .B1(n2791), .B2(n369), .ZN(n2272) );
  OAI22_X2 U1881 ( .A1(n417), .A2(n2793), .B1(n2792), .B2(n369), .ZN(n2273) );
  XNOR2_X2 U1882 ( .A(n3059), .B(n323), .ZN(n2762) );
  XNOR2_X2 U1883 ( .A(n3060), .B(n323), .ZN(n2763) );
  XNOR2_X2 U1884 ( .A(n3061), .B(n323), .ZN(n2764) );
  XNOR2_X2 U1885 ( .A(n3062), .B(n323), .ZN(n2765) );
  XNOR2_X2 U1886 ( .A(n3063), .B(n323), .ZN(n2766) );
  XNOR2_X2 U1887 ( .A(n3064), .B(n323), .ZN(n2767) );
  XNOR2_X2 U1888 ( .A(n3065), .B(n323), .ZN(n2768) );
  XNOR2_X2 U1889 ( .A(n3066), .B(n323), .ZN(n2769) );
  XNOR2_X2 U1890 ( .A(n3067), .B(n323), .ZN(n2770) );
  XNOR2_X2 U1891 ( .A(n3068), .B(n323), .ZN(n2771) );
  XNOR2_X2 U1892 ( .A(n3069), .B(n323), .ZN(n2772) );
  XNOR2_X2 U1893 ( .A(n3070), .B(n322), .ZN(n2773) );
  XNOR2_X2 U1894 ( .A(n3071), .B(n322), .ZN(n2774) );
  XNOR2_X2 U1895 ( .A(n3072), .B(n322), .ZN(n2775) );
  XNOR2_X2 U1896 ( .A(n3073), .B(n322), .ZN(n2776) );
  XNOR2_X2 U1897 ( .A(n3074), .B(n322), .ZN(n2777) );
  XNOR2_X2 U1898 ( .A(n3075), .B(n322), .ZN(n2778) );
  XNOR2_X2 U1899 ( .A(n3076), .B(n322), .ZN(n2779) );
  XNOR2_X2 U1900 ( .A(n3077), .B(n322), .ZN(n2780) );
  XNOR2_X2 U1901 ( .A(n3078), .B(n322), .ZN(n2781) );
  XNOR2_X2 U1902 ( .A(n3079), .B(n322), .ZN(n2782) );
  XNOR2_X2 U1903 ( .A(n3080), .B(n322), .ZN(n2783) );
  XNOR2_X2 U1904 ( .A(n3081), .B(n322), .ZN(n2784) );
  XNOR2_X2 U1905 ( .A(n3082), .B(n321), .ZN(n2785) );
  XNOR2_X2 U1906 ( .A(n3083), .B(n321), .ZN(n2786) );
  XNOR2_X2 U1907 ( .A(n3084), .B(n321), .ZN(n2787) );
  XNOR2_X2 U1908 ( .A(n3085), .B(n321), .ZN(n2788) );
  XNOR2_X2 U1909 ( .A(n3086), .B(n321), .ZN(n2789) );
  XNOR2_X2 U1910 ( .A(n3087), .B(n321), .ZN(n2790) );
  XNOR2_X2 U1911 ( .A(n3088), .B(n321), .ZN(n2791) );
  XNOR2_X2 U1912 ( .A(n3089), .B(n321), .ZN(n2792) );
  XNOR2_X2 U1913 ( .A(n441), .B(n321), .ZN(n2793) );
  OAI22_X2 U1914 ( .A1(n416), .A2(n3147), .B1(n2827), .B2(n368), .ZN(n2011) );
  OAI22_X2 U1916 ( .A1(n416), .A2(n2797), .B1(n2796), .B2(n368), .ZN(n2276) );
  OAI22_X2 U1917 ( .A1(n416), .A2(n2798), .B1(n2797), .B2(n368), .ZN(n2277) );
  OAI22_X2 U1918 ( .A1(n416), .A2(n2799), .B1(n2798), .B2(n368), .ZN(n2278) );
  OAI22_X2 U1919 ( .A1(n416), .A2(n2800), .B1(n2799), .B2(n368), .ZN(n2279) );
  OAI22_X2 U1920 ( .A1(n416), .A2(n2801), .B1(n2800), .B2(n368), .ZN(n2280) );
  OAI22_X2 U1921 ( .A1(n416), .A2(n2802), .B1(n2801), .B2(n368), .ZN(n2281) );
  OAI22_X2 U1922 ( .A1(n416), .A2(n2803), .B1(n2802), .B2(n368), .ZN(n2282) );
  OAI22_X2 U1923 ( .A1(n416), .A2(n2804), .B1(n2803), .B2(n368), .ZN(n2283) );
  OAI22_X2 U1924 ( .A1(n415), .A2(n2805), .B1(n2804), .B2(n367), .ZN(n2284) );
  OAI22_X2 U1925 ( .A1(n415), .A2(n2806), .B1(n2805), .B2(n367), .ZN(n2285) );
  OAI22_X2 U1926 ( .A1(n415), .A2(n2807), .B1(n2806), .B2(n367), .ZN(n2286) );
  OAI22_X2 U1927 ( .A1(n415), .A2(n2808), .B1(n2807), .B2(n367), .ZN(n2287) );
  OAI22_X2 U1928 ( .A1(n415), .A2(n2809), .B1(n2808), .B2(n367), .ZN(n2288) );
  OAI22_X2 U1929 ( .A1(n415), .A2(n2810), .B1(n2809), .B2(n367), .ZN(n2289) );
  OAI22_X2 U1930 ( .A1(n415), .A2(n2811), .B1(n2810), .B2(n367), .ZN(n2290) );
  OAI22_X2 U1931 ( .A1(n415), .A2(n2812), .B1(n2811), .B2(n367), .ZN(n2291) );
  OAI22_X2 U1932 ( .A1(n415), .A2(n2813), .B1(n2812), .B2(n367), .ZN(n2292) );
  OAI22_X2 U1933 ( .A1(n415), .A2(n2814), .B1(n2813), .B2(n367), .ZN(n2293) );
  OAI22_X2 U1934 ( .A1(n415), .A2(n2815), .B1(n2814), .B2(n367), .ZN(n2294) );
  OAI22_X2 U1935 ( .A1(n414), .A2(n2816), .B1(n2815), .B2(n367), .ZN(n2295) );
  OAI22_X2 U1936 ( .A1(n414), .A2(n2817), .B1(n2816), .B2(n366), .ZN(n2296) );
  OAI22_X2 U1937 ( .A1(n414), .A2(n2818), .B1(n2817), .B2(n366), .ZN(n2297) );
  OAI22_X2 U1938 ( .A1(n414), .A2(n2819), .B1(n2818), .B2(n366), .ZN(n2298) );
  OAI22_X2 U1939 ( .A1(n414), .A2(n2820), .B1(n2819), .B2(n366), .ZN(n2299) );
  OAI22_X2 U1940 ( .A1(n414), .A2(n2821), .B1(n2820), .B2(n366), .ZN(n2300) );
  OAI22_X2 U1941 ( .A1(n414), .A2(n2822), .B1(n2821), .B2(n366), .ZN(n2301) );
  OAI22_X2 U1942 ( .A1(n414), .A2(n2823), .B1(n2822), .B2(n366), .ZN(n2302) );
  OAI22_X2 U1943 ( .A1(n414), .A2(n2824), .B1(n2823), .B2(n366), .ZN(n2303) );
  OAI22_X2 U1944 ( .A1(n414), .A2(n2825), .B1(n2824), .B2(n366), .ZN(n2304) );
  OAI22_X2 U1945 ( .A1(n414), .A2(n2826), .B1(n2825), .B2(n366), .ZN(n2305) );
  XNOR2_X2 U1946 ( .A(n3059), .B(n320), .ZN(n2795) );
  XNOR2_X2 U1947 ( .A(n3060), .B(n320), .ZN(n2796) );
  XNOR2_X2 U1948 ( .A(n3061), .B(n320), .ZN(n2797) );
  XNOR2_X2 U1949 ( .A(n3062), .B(n320), .ZN(n2798) );
  XNOR2_X2 U1950 ( .A(n3063), .B(n320), .ZN(n2799) );
  XNOR2_X2 U1951 ( .A(n3064), .B(n320), .ZN(n2800) );
  XNOR2_X2 U1952 ( .A(n3065), .B(n320), .ZN(n2801) );
  XNOR2_X2 U1953 ( .A(n3066), .B(n320), .ZN(n2802) );
  XNOR2_X2 U1954 ( .A(n3067), .B(n320), .ZN(n2803) );
  XNOR2_X2 U1955 ( .A(n3068), .B(n320), .ZN(n2804) );
  XNOR2_X2 U1956 ( .A(n3069), .B(n320), .ZN(n2805) );
  XNOR2_X2 U1957 ( .A(n3070), .B(n319), .ZN(n2806) );
  XNOR2_X2 U1958 ( .A(n3071), .B(n319), .ZN(n2807) );
  XNOR2_X2 U1959 ( .A(n3072), .B(n319), .ZN(n2808) );
  XNOR2_X2 U1960 ( .A(n3073), .B(n319), .ZN(n2809) );
  XNOR2_X2 U1961 ( .A(n3074), .B(n319), .ZN(n2810) );
  XNOR2_X2 U1962 ( .A(n3075), .B(n319), .ZN(n2811) );
  XNOR2_X2 U1963 ( .A(n3076), .B(n319), .ZN(n2812) );
  XNOR2_X2 U1964 ( .A(n3077), .B(n319), .ZN(n2813) );
  XNOR2_X2 U1965 ( .A(n3078), .B(n319), .ZN(n2814) );
  XNOR2_X2 U1966 ( .A(n3079), .B(n319), .ZN(n2815) );
  XNOR2_X2 U1967 ( .A(n3080), .B(n319), .ZN(n2816) );
  XNOR2_X2 U1968 ( .A(n3081), .B(n319), .ZN(n2817) );
  XNOR2_X2 U1969 ( .A(n3082), .B(n318), .ZN(n2818) );
  XNOR2_X2 U1970 ( .A(n3083), .B(n318), .ZN(n2819) );
  XNOR2_X2 U1971 ( .A(n3084), .B(n318), .ZN(n2820) );
  XNOR2_X2 U1972 ( .A(n3085), .B(n318), .ZN(n2821) );
  XNOR2_X2 U1973 ( .A(n3086), .B(n318), .ZN(n2822) );
  XNOR2_X2 U1974 ( .A(n3087), .B(n318), .ZN(n2823) );
  XNOR2_X2 U1975 ( .A(n3088), .B(n318), .ZN(n2824) );
  XNOR2_X2 U1976 ( .A(n3089), .B(n318), .ZN(n2825) );
  XNOR2_X2 U1977 ( .A(n441), .B(n318), .ZN(n2826) );
  OAI22_X2 U1978 ( .A1(n413), .A2(n3148), .B1(n2860), .B2(n365), .ZN(n2012) );
  OAI22_X2 U1980 ( .A1(n413), .A2(n2830), .B1(n2829), .B2(n365), .ZN(n2308) );
  OAI22_X2 U1981 ( .A1(n413), .A2(n2831), .B1(n2830), .B2(n365), .ZN(n2309) );
  OAI22_X2 U1982 ( .A1(n413), .A2(n2832), .B1(n2831), .B2(n365), .ZN(n2310) );
  OAI22_X2 U1983 ( .A1(n413), .A2(n2833), .B1(n2832), .B2(n365), .ZN(n2311) );
  OAI22_X2 U1984 ( .A1(n413), .A2(n2834), .B1(n2833), .B2(n365), .ZN(n2312) );
  OAI22_X2 U1985 ( .A1(n413), .A2(n2835), .B1(n2834), .B2(n365), .ZN(n2313) );
  OAI22_X2 U1986 ( .A1(n413), .A2(n2836), .B1(n2835), .B2(n365), .ZN(n2314) );
  OAI22_X2 U1987 ( .A1(n413), .A2(n2837), .B1(n2836), .B2(n365), .ZN(n2315) );
  OAI22_X2 U1988 ( .A1(n412), .A2(n2838), .B1(n2837), .B2(n364), .ZN(n2316) );
  OAI22_X2 U1989 ( .A1(n412), .A2(n2839), .B1(n2838), .B2(n364), .ZN(n2317) );
  OAI22_X2 U1990 ( .A1(n412), .A2(n2840), .B1(n2839), .B2(n364), .ZN(n2318) );
  OAI22_X2 U1991 ( .A1(n412), .A2(n2841), .B1(n2840), .B2(n364), .ZN(n2319) );
  OAI22_X2 U1992 ( .A1(n412), .A2(n2842), .B1(n2841), .B2(n364), .ZN(n2320) );
  OAI22_X2 U1993 ( .A1(n412), .A2(n2843), .B1(n2842), .B2(n364), .ZN(n2321) );
  OAI22_X2 U1994 ( .A1(n412), .A2(n2844), .B1(n2843), .B2(n364), .ZN(n2322) );
  OAI22_X2 U1995 ( .A1(n412), .A2(n2845), .B1(n2844), .B2(n364), .ZN(n2323) );
  OAI22_X2 U1996 ( .A1(n412), .A2(n2846), .B1(n2845), .B2(n364), .ZN(n2324) );
  OAI22_X2 U1997 ( .A1(n412), .A2(n2847), .B1(n2846), .B2(n364), .ZN(n2325) );
  OAI22_X2 U1998 ( .A1(n412), .A2(n2848), .B1(n2847), .B2(n364), .ZN(n2326) );
  OAI22_X2 U1999 ( .A1(n411), .A2(n2849), .B1(n2848), .B2(n364), .ZN(n2327) );
  OAI22_X2 U2000 ( .A1(n411), .A2(n2850), .B1(n2849), .B2(n363), .ZN(n2328) );
  OAI22_X2 U2001 ( .A1(n411), .A2(n2851), .B1(n2850), .B2(n363), .ZN(n2329) );
  OAI22_X2 U2002 ( .A1(n411), .A2(n2852), .B1(n2851), .B2(n363), .ZN(n2330) );
  OAI22_X2 U2003 ( .A1(n411), .A2(n2853), .B1(n2852), .B2(n363), .ZN(n2331) );
  OAI22_X2 U2004 ( .A1(n411), .A2(n2854), .B1(n2853), .B2(n363), .ZN(n2332) );
  OAI22_X2 U2005 ( .A1(n411), .A2(n2855), .B1(n2854), .B2(n363), .ZN(n2333) );
  OAI22_X2 U2006 ( .A1(n411), .A2(n2856), .B1(n2855), .B2(n363), .ZN(n2334) );
  OAI22_X2 U2007 ( .A1(n411), .A2(n2857), .B1(n2856), .B2(n363), .ZN(n2335) );
  OAI22_X2 U2008 ( .A1(n411), .A2(n2858), .B1(n2857), .B2(n363), .ZN(n2336) );
  OAI22_X2 U2009 ( .A1(n411), .A2(n2859), .B1(n2858), .B2(n363), .ZN(n2337) );
  XNOR2_X2 U2010 ( .A(n3059), .B(n317), .ZN(n2828) );
  XNOR2_X2 U2011 ( .A(n3060), .B(n317), .ZN(n2829) );
  XNOR2_X2 U2012 ( .A(n3061), .B(n317), .ZN(n2830) );
  XNOR2_X2 U2013 ( .A(n3062), .B(n317), .ZN(n2831) );
  XNOR2_X2 U2014 ( .A(n3063), .B(n317), .ZN(n2832) );
  XNOR2_X2 U2015 ( .A(n3064), .B(n317), .ZN(n2833) );
  XNOR2_X2 U2016 ( .A(n3065), .B(n317), .ZN(n2834) );
  XNOR2_X2 U2017 ( .A(n3066), .B(n317), .ZN(n2835) );
  XNOR2_X2 U2018 ( .A(n3067), .B(n317), .ZN(n2836) );
  XNOR2_X2 U2019 ( .A(n3068), .B(n317), .ZN(n2837) );
  XNOR2_X2 U2020 ( .A(n3069), .B(n317), .ZN(n2838) );
  XNOR2_X2 U2021 ( .A(n3070), .B(n316), .ZN(n2839) );
  XNOR2_X2 U2022 ( .A(n3071), .B(n316), .ZN(n2840) );
  XNOR2_X2 U2023 ( .A(n3072), .B(n316), .ZN(n2841) );
  XNOR2_X2 U2024 ( .A(n3073), .B(n316), .ZN(n2842) );
  XNOR2_X2 U2025 ( .A(n3074), .B(n316), .ZN(n2843) );
  XNOR2_X2 U2026 ( .A(n3075), .B(n316), .ZN(n2844) );
  XNOR2_X2 U2027 ( .A(n3076), .B(n316), .ZN(n2845) );
  XNOR2_X2 U2028 ( .A(n3077), .B(n316), .ZN(n2846) );
  XNOR2_X2 U2029 ( .A(n3078), .B(n316), .ZN(n2847) );
  XNOR2_X2 U2030 ( .A(n3079), .B(n316), .ZN(n2848) );
  XNOR2_X2 U2031 ( .A(n3080), .B(n316), .ZN(n2849) );
  XNOR2_X2 U2032 ( .A(n3081), .B(n316), .ZN(n2850) );
  XNOR2_X2 U2033 ( .A(n3082), .B(n315), .ZN(n2851) );
  XNOR2_X2 U2034 ( .A(n3083), .B(n315), .ZN(n2852) );
  XNOR2_X2 U2035 ( .A(n3084), .B(n315), .ZN(n2853) );
  XNOR2_X2 U2036 ( .A(n3085), .B(n315), .ZN(n2854) );
  XNOR2_X2 U2037 ( .A(n3086), .B(n315), .ZN(n2855) );
  XNOR2_X2 U2038 ( .A(n3087), .B(n315), .ZN(n2856) );
  XNOR2_X2 U2039 ( .A(n3088), .B(n315), .ZN(n2857) );
  XNOR2_X2 U2040 ( .A(n3089), .B(n315), .ZN(n2858) );
  XNOR2_X2 U2041 ( .A(n441), .B(n315), .ZN(n2859) );
  OAI22_X2 U2042 ( .A1(n410), .A2(n3149), .B1(n2893), .B2(n362), .ZN(n2013) );
  OAI22_X2 U2044 ( .A1(n410), .A2(n2863), .B1(n2862), .B2(n362), .ZN(n2340) );
  OAI22_X2 U2045 ( .A1(n410), .A2(n2864), .B1(n2863), .B2(n362), .ZN(n2341) );
  OAI22_X2 U2046 ( .A1(n410), .A2(n2865), .B1(n2864), .B2(n362), .ZN(n2342) );
  OAI22_X2 U2047 ( .A1(n410), .A2(n2866), .B1(n2865), .B2(n362), .ZN(n2343) );
  OAI22_X2 U2048 ( .A1(n410), .A2(n2867), .B1(n2866), .B2(n362), .ZN(n2344) );
  OAI22_X2 U2049 ( .A1(n410), .A2(n2868), .B1(n2867), .B2(n362), .ZN(n2345) );
  OAI22_X2 U2050 ( .A1(n410), .A2(n2869), .B1(n2868), .B2(n362), .ZN(n2346) );
  OAI22_X2 U2051 ( .A1(n410), .A2(n2870), .B1(n2869), .B2(n362), .ZN(n2347) );
  OAI22_X2 U2052 ( .A1(n409), .A2(n2871), .B1(n2870), .B2(n361), .ZN(n2348) );
  OAI22_X2 U2053 ( .A1(n409), .A2(n2872), .B1(n2871), .B2(n361), .ZN(n2349) );
  OAI22_X2 U2054 ( .A1(n409), .A2(n2873), .B1(n2872), .B2(n361), .ZN(n2350) );
  OAI22_X2 U2055 ( .A1(n409), .A2(n2874), .B1(n2873), .B2(n361), .ZN(n2351) );
  OAI22_X2 U2056 ( .A1(n409), .A2(n2875), .B1(n2874), .B2(n361), .ZN(n2352) );
  OAI22_X2 U2057 ( .A1(n409), .A2(n2876), .B1(n2875), .B2(n361), .ZN(n2353) );
  OAI22_X2 U2058 ( .A1(n409), .A2(n2877), .B1(n2876), .B2(n361), .ZN(n2354) );
  OAI22_X2 U2059 ( .A1(n409), .A2(n2878), .B1(n2877), .B2(n361), .ZN(n2355) );
  OAI22_X2 U2060 ( .A1(n409), .A2(n2879), .B1(n2878), .B2(n361), .ZN(n2356) );
  OAI22_X2 U2061 ( .A1(n409), .A2(n2880), .B1(n2879), .B2(n361), .ZN(n2357) );
  OAI22_X2 U2062 ( .A1(n409), .A2(n2881), .B1(n2880), .B2(n361), .ZN(n2358) );
  OAI22_X2 U2063 ( .A1(n408), .A2(n2882), .B1(n2881), .B2(n361), .ZN(n2359) );
  OAI22_X2 U2064 ( .A1(n408), .A2(n2883), .B1(n2882), .B2(n360), .ZN(n2360) );
  OAI22_X2 U2065 ( .A1(n408), .A2(n2884), .B1(n2883), .B2(n360), .ZN(n2361) );
  OAI22_X2 U2066 ( .A1(n408), .A2(n2885), .B1(n2884), .B2(n360), .ZN(n2362) );
  OAI22_X2 U2067 ( .A1(n408), .A2(n2886), .B1(n2885), .B2(n360), .ZN(n2363) );
  OAI22_X2 U2068 ( .A1(n408), .A2(n2887), .B1(n2886), .B2(n360), .ZN(n2364) );
  OAI22_X2 U2069 ( .A1(n408), .A2(n2888), .B1(n2887), .B2(n360), .ZN(n2365) );
  OAI22_X2 U2070 ( .A1(n408), .A2(n2889), .B1(n2888), .B2(n360), .ZN(n2366) );
  OAI22_X2 U2071 ( .A1(n408), .A2(n2890), .B1(n2889), .B2(n360), .ZN(n2367) );
  OAI22_X2 U2072 ( .A1(n408), .A2(n2891), .B1(n2890), .B2(n360), .ZN(n2368) );
  OAI22_X2 U2073 ( .A1(n408), .A2(n2892), .B1(n2891), .B2(n360), .ZN(n2369) );
  XNOR2_X2 U2074 ( .A(n3059), .B(n314), .ZN(n2861) );
  XNOR2_X2 U2075 ( .A(n3060), .B(n314), .ZN(n2862) );
  XNOR2_X2 U2076 ( .A(n3061), .B(n314), .ZN(n2863) );
  XNOR2_X2 U2077 ( .A(n3062), .B(n314), .ZN(n2864) );
  XNOR2_X2 U2078 ( .A(n3063), .B(n314), .ZN(n2865) );
  XNOR2_X2 U2079 ( .A(n3064), .B(n314), .ZN(n2866) );
  XNOR2_X2 U2080 ( .A(n3065), .B(n314), .ZN(n2867) );
  XNOR2_X2 U2081 ( .A(n3066), .B(n314), .ZN(n2868) );
  XNOR2_X2 U2082 ( .A(n3067), .B(n314), .ZN(n2869) );
  XNOR2_X2 U2083 ( .A(n3068), .B(n314), .ZN(n2870) );
  XNOR2_X2 U2084 ( .A(n3069), .B(n314), .ZN(n2871) );
  XNOR2_X2 U2085 ( .A(n3070), .B(n313), .ZN(n2872) );
  XNOR2_X2 U2086 ( .A(n3071), .B(n313), .ZN(n2873) );
  XNOR2_X2 U2087 ( .A(n3072), .B(n313), .ZN(n2874) );
  XNOR2_X2 U2088 ( .A(n3073), .B(n313), .ZN(n2875) );
  XNOR2_X2 U2089 ( .A(n3074), .B(n313), .ZN(n2876) );
  XNOR2_X2 U2090 ( .A(n3075), .B(n313), .ZN(n2877) );
  XNOR2_X2 U2091 ( .A(n3076), .B(n313), .ZN(n2878) );
  XNOR2_X2 U2092 ( .A(n3077), .B(n313), .ZN(n2879) );
  XNOR2_X2 U2093 ( .A(n3078), .B(n313), .ZN(n2880) );
  XNOR2_X2 U2094 ( .A(n3079), .B(n313), .ZN(n2881) );
  XNOR2_X2 U2095 ( .A(n3080), .B(n313), .ZN(n2882) );
  XNOR2_X2 U2096 ( .A(n3081), .B(n313), .ZN(n2883) );
  XNOR2_X2 U2097 ( .A(n3082), .B(n312), .ZN(n2884) );
  XNOR2_X2 U2098 ( .A(n3083), .B(n312), .ZN(n2885) );
  XNOR2_X2 U2099 ( .A(n3084), .B(n312), .ZN(n2886) );
  XNOR2_X2 U2100 ( .A(n3085), .B(n312), .ZN(n2887) );
  XNOR2_X2 U2101 ( .A(n3086), .B(n312), .ZN(n2888) );
  XNOR2_X2 U2102 ( .A(n3087), .B(n312), .ZN(n2889) );
  XNOR2_X2 U2103 ( .A(n3088), .B(n312), .ZN(n2890) );
  XNOR2_X2 U2104 ( .A(n3089), .B(n312), .ZN(n2891) );
  XNOR2_X2 U2105 ( .A(n441), .B(n312), .ZN(n2892) );
  OAI22_X2 U2106 ( .A1(n407), .A2(n3150), .B1(n2926), .B2(n359), .ZN(n2014) );
  OAI22_X2 U2108 ( .A1(n407), .A2(n2896), .B1(n2895), .B2(n359), .ZN(n2372) );
  OAI22_X2 U2109 ( .A1(n407), .A2(n2897), .B1(n2896), .B2(n359), .ZN(n2373) );
  OAI22_X2 U2110 ( .A1(n407), .A2(n2898), .B1(n2897), .B2(n359), .ZN(n2374) );
  OAI22_X2 U2111 ( .A1(n407), .A2(n2899), .B1(n2898), .B2(n359), .ZN(n2375) );
  OAI22_X2 U2112 ( .A1(n407), .A2(n2900), .B1(n2899), .B2(n359), .ZN(n2376) );
  OAI22_X2 U2113 ( .A1(n407), .A2(n2901), .B1(n2900), .B2(n359), .ZN(n2377) );
  OAI22_X2 U2114 ( .A1(n407), .A2(n2902), .B1(n2901), .B2(n359), .ZN(n2378) );
  OAI22_X2 U2115 ( .A1(n407), .A2(n2903), .B1(n2902), .B2(n359), .ZN(n2379) );
  OAI22_X2 U2116 ( .A1(n406), .A2(n2904), .B1(n2903), .B2(n358), .ZN(n2380) );
  OAI22_X2 U2117 ( .A1(n406), .A2(n2905), .B1(n2904), .B2(n358), .ZN(n2381) );
  OAI22_X2 U2118 ( .A1(n406), .A2(n2906), .B1(n2905), .B2(n358), .ZN(n2382) );
  OAI22_X2 U2119 ( .A1(n406), .A2(n2907), .B1(n2906), .B2(n358), .ZN(n2383) );
  OAI22_X2 U2120 ( .A1(n406), .A2(n2908), .B1(n2907), .B2(n358), .ZN(n2384) );
  OAI22_X2 U2121 ( .A1(n406), .A2(n2909), .B1(n2908), .B2(n358), .ZN(n2385) );
  OAI22_X2 U2122 ( .A1(n406), .A2(n2910), .B1(n2909), .B2(n358), .ZN(n2386) );
  OAI22_X2 U2123 ( .A1(n406), .A2(n2911), .B1(n2910), .B2(n358), .ZN(n2387) );
  OAI22_X2 U2124 ( .A1(n406), .A2(n2912), .B1(n2911), .B2(n358), .ZN(n2388) );
  OAI22_X2 U2125 ( .A1(n406), .A2(n2913), .B1(n2912), .B2(n358), .ZN(n2389) );
  OAI22_X2 U2126 ( .A1(n406), .A2(n2914), .B1(n2913), .B2(n358), .ZN(n2390) );
  OAI22_X2 U2127 ( .A1(n405), .A2(n2915), .B1(n2914), .B2(n358), .ZN(n2391) );
  OAI22_X2 U2128 ( .A1(n405), .A2(n2916), .B1(n2915), .B2(n357), .ZN(n2392) );
  OAI22_X2 U2129 ( .A1(n405), .A2(n2917), .B1(n2916), .B2(n357), .ZN(n2393) );
  OAI22_X2 U2130 ( .A1(n405), .A2(n2918), .B1(n2917), .B2(n357), .ZN(n2394) );
  OAI22_X2 U2131 ( .A1(n405), .A2(n2919), .B1(n2918), .B2(n357), .ZN(n2395) );
  OAI22_X2 U2132 ( .A1(n405), .A2(n2920), .B1(n2919), .B2(n357), .ZN(n2396) );
  OAI22_X2 U2133 ( .A1(n405), .A2(n2921), .B1(n2920), .B2(n357), .ZN(n2397) );
  OAI22_X2 U2134 ( .A1(n405), .A2(n2922), .B1(n2921), .B2(n357), .ZN(n2398) );
  OAI22_X2 U2135 ( .A1(n405), .A2(n2923), .B1(n2922), .B2(n357), .ZN(n2399) );
  OAI22_X2 U2136 ( .A1(n405), .A2(n2924), .B1(n2923), .B2(n357), .ZN(n2400) );
  OAI22_X2 U2137 ( .A1(n405), .A2(n2925), .B1(n2924), .B2(n357), .ZN(n2401) );
  XNOR2_X2 U2138 ( .A(n3059), .B(n311), .ZN(n2894) );
  XNOR2_X2 U2139 ( .A(n3060), .B(n311), .ZN(n2895) );
  XNOR2_X2 U2140 ( .A(n3061), .B(n311), .ZN(n2896) );
  XNOR2_X2 U2141 ( .A(n3062), .B(n311), .ZN(n2897) );
  XNOR2_X2 U2142 ( .A(n3063), .B(n311), .ZN(n2898) );
  XNOR2_X2 U2143 ( .A(n3064), .B(n311), .ZN(n2899) );
  XNOR2_X2 U2144 ( .A(n3065), .B(n311), .ZN(n2900) );
  XNOR2_X2 U2145 ( .A(n3066), .B(n311), .ZN(n2901) );
  XNOR2_X2 U2146 ( .A(n3067), .B(n311), .ZN(n2902) );
  XNOR2_X2 U2147 ( .A(n3068), .B(n311), .ZN(n2903) );
  XNOR2_X2 U2148 ( .A(n3069), .B(n311), .ZN(n2904) );
  XNOR2_X2 U2149 ( .A(n3070), .B(n310), .ZN(n2905) );
  XNOR2_X2 U2150 ( .A(n3071), .B(n310), .ZN(n2906) );
  XNOR2_X2 U2151 ( .A(n3072), .B(n310), .ZN(n2907) );
  XNOR2_X2 U2152 ( .A(n3073), .B(n310), .ZN(n2908) );
  XNOR2_X2 U2153 ( .A(n3074), .B(n310), .ZN(n2909) );
  XNOR2_X2 U2154 ( .A(n3075), .B(n310), .ZN(n2910) );
  XNOR2_X2 U2155 ( .A(n3076), .B(n310), .ZN(n2911) );
  XNOR2_X2 U2156 ( .A(n3077), .B(n310), .ZN(n2912) );
  XNOR2_X2 U2157 ( .A(n3078), .B(n310), .ZN(n2913) );
  XNOR2_X2 U2158 ( .A(n3079), .B(n310), .ZN(n2914) );
  XNOR2_X2 U2159 ( .A(n3080), .B(n310), .ZN(n2915) );
  XNOR2_X2 U2160 ( .A(n3081), .B(n310), .ZN(n2916) );
  XNOR2_X2 U2161 ( .A(n3082), .B(n309), .ZN(n2917) );
  XNOR2_X2 U2162 ( .A(n3083), .B(n309), .ZN(n2918) );
  XNOR2_X2 U2163 ( .A(n3084), .B(n309), .ZN(n2919) );
  XNOR2_X2 U2164 ( .A(n3085), .B(n309), .ZN(n2920) );
  XNOR2_X2 U2165 ( .A(n3086), .B(n309), .ZN(n2921) );
  XNOR2_X2 U2166 ( .A(n3087), .B(n309), .ZN(n2922) );
  XNOR2_X2 U2167 ( .A(n3088), .B(n309), .ZN(n2923) );
  XNOR2_X2 U2168 ( .A(n3089), .B(n309), .ZN(n2924) );
  XNOR2_X2 U2169 ( .A(n441), .B(n309), .ZN(n2925) );
  OAI22_X2 U2170 ( .A1(n404), .A2(n3151), .B1(n2959), .B2(n356), .ZN(n2015) );
  OAI22_X2 U2172 ( .A1(n404), .A2(n2929), .B1(n2928), .B2(n356), .ZN(n2404) );
  OAI22_X2 U2173 ( .A1(n404), .A2(n2930), .B1(n2929), .B2(n356), .ZN(n2405) );
  OAI22_X2 U2174 ( .A1(n404), .A2(n2931), .B1(n2930), .B2(n356), .ZN(n2406) );
  OAI22_X2 U2175 ( .A1(n404), .A2(n2932), .B1(n2931), .B2(n356), .ZN(n2407) );
  OAI22_X2 U2176 ( .A1(n404), .A2(n2933), .B1(n2932), .B2(n356), .ZN(n2408) );
  OAI22_X2 U2177 ( .A1(n404), .A2(n2934), .B1(n2933), .B2(n356), .ZN(n2409) );
  OAI22_X2 U2178 ( .A1(n404), .A2(n2935), .B1(n2934), .B2(n356), .ZN(n2410) );
  OAI22_X2 U2179 ( .A1(n404), .A2(n2936), .B1(n2935), .B2(n356), .ZN(n2411) );
  OAI22_X2 U2180 ( .A1(n403), .A2(n2937), .B1(n2936), .B2(n355), .ZN(n2412) );
  OAI22_X2 U2181 ( .A1(n403), .A2(n2938), .B1(n2937), .B2(n355), .ZN(n2413) );
  OAI22_X2 U2182 ( .A1(n403), .A2(n2939), .B1(n2938), .B2(n355), .ZN(n2414) );
  OAI22_X2 U2183 ( .A1(n403), .A2(n2940), .B1(n2939), .B2(n355), .ZN(n2415) );
  OAI22_X2 U2184 ( .A1(n403), .A2(n2941), .B1(n2940), .B2(n355), .ZN(n2416) );
  OAI22_X2 U2185 ( .A1(n403), .A2(n2942), .B1(n2941), .B2(n355), .ZN(n2417) );
  OAI22_X2 U2186 ( .A1(n403), .A2(n2943), .B1(n2942), .B2(n355), .ZN(n2418) );
  OAI22_X2 U2187 ( .A1(n403), .A2(n2944), .B1(n2943), .B2(n355), .ZN(n2419) );
  OAI22_X2 U2188 ( .A1(n403), .A2(n2945), .B1(n2944), .B2(n355), .ZN(n2420) );
  OAI22_X2 U2189 ( .A1(n403), .A2(n2946), .B1(n2945), .B2(n355), .ZN(n2421) );
  OAI22_X2 U2190 ( .A1(n403), .A2(n2947), .B1(n2946), .B2(n355), .ZN(n2422) );
  OAI22_X2 U2191 ( .A1(n402), .A2(n2948), .B1(n2947), .B2(n355), .ZN(n2423) );
  OAI22_X2 U2192 ( .A1(n402), .A2(n2949), .B1(n2948), .B2(n354), .ZN(n2424) );
  OAI22_X2 U2193 ( .A1(n402), .A2(n2950), .B1(n2949), .B2(n354), .ZN(n2425) );
  OAI22_X2 U2194 ( .A1(n402), .A2(n2951), .B1(n2950), .B2(n354), .ZN(n2426) );
  OAI22_X2 U2195 ( .A1(n402), .A2(n2952), .B1(n2951), .B2(n354), .ZN(n2427) );
  OAI22_X2 U2196 ( .A1(n402), .A2(n2953), .B1(n2952), .B2(n354), .ZN(n2428) );
  OAI22_X2 U2197 ( .A1(n402), .A2(n2954), .B1(n2953), .B2(n354), .ZN(n2429) );
  OAI22_X2 U2198 ( .A1(n402), .A2(n2955), .B1(n2954), .B2(n354), .ZN(n2430) );
  OAI22_X2 U2199 ( .A1(n402), .A2(n2956), .B1(n2955), .B2(n354), .ZN(n2431) );
  OAI22_X2 U2200 ( .A1(n402), .A2(n2957), .B1(n2956), .B2(n354), .ZN(n2432) );
  OAI22_X2 U2201 ( .A1(n402), .A2(n2958), .B1(n2957), .B2(n354), .ZN(n2433) );
  XNOR2_X2 U2202 ( .A(n3059), .B(n308), .ZN(n2927) );
  XNOR2_X2 U2203 ( .A(n3060), .B(n308), .ZN(n2928) );
  XNOR2_X2 U2204 ( .A(n3061), .B(n308), .ZN(n2929) );
  XNOR2_X2 U2205 ( .A(n3062), .B(n308), .ZN(n2930) );
  XNOR2_X2 U2206 ( .A(n3063), .B(n308), .ZN(n2931) );
  XNOR2_X2 U2207 ( .A(n3064), .B(n308), .ZN(n2932) );
  XNOR2_X2 U2208 ( .A(n3065), .B(n308), .ZN(n2933) );
  XNOR2_X2 U2209 ( .A(n3066), .B(n308), .ZN(n2934) );
  XNOR2_X2 U2210 ( .A(n3067), .B(n308), .ZN(n2935) );
  XNOR2_X2 U2211 ( .A(n3068), .B(n308), .ZN(n2936) );
  XNOR2_X2 U2212 ( .A(n3069), .B(n308), .ZN(n2937) );
  XNOR2_X2 U2213 ( .A(n3070), .B(n307), .ZN(n2938) );
  XNOR2_X2 U2214 ( .A(n3071), .B(n307), .ZN(n2939) );
  XNOR2_X2 U2215 ( .A(n3072), .B(n307), .ZN(n2940) );
  XNOR2_X2 U2216 ( .A(n3073), .B(n307), .ZN(n2941) );
  XNOR2_X2 U2217 ( .A(n3074), .B(n307), .ZN(n2942) );
  XNOR2_X2 U2218 ( .A(n3075), .B(n307), .ZN(n2943) );
  XNOR2_X2 U2219 ( .A(n3076), .B(n307), .ZN(n2944) );
  XNOR2_X2 U2220 ( .A(n3077), .B(n307), .ZN(n2945) );
  XNOR2_X2 U2221 ( .A(n3078), .B(n307), .ZN(n2946) );
  XNOR2_X2 U2222 ( .A(n3079), .B(n307), .ZN(n2947) );
  XNOR2_X2 U2223 ( .A(n3080), .B(n307), .ZN(n2948) );
  XNOR2_X2 U2224 ( .A(n3081), .B(n307), .ZN(n2949) );
  XNOR2_X2 U2225 ( .A(n3082), .B(n306), .ZN(n2950) );
  XNOR2_X2 U2226 ( .A(n3083), .B(n306), .ZN(n2951) );
  XNOR2_X2 U2227 ( .A(n3084), .B(n306), .ZN(n2952) );
  XNOR2_X2 U2228 ( .A(n3085), .B(n306), .ZN(n2953) );
  XNOR2_X2 U2229 ( .A(n3086), .B(n306), .ZN(n2954) );
  XNOR2_X2 U2230 ( .A(n3087), .B(n306), .ZN(n2955) );
  XNOR2_X2 U2231 ( .A(n3088), .B(n306), .ZN(n2956) );
  XNOR2_X2 U2232 ( .A(n3089), .B(n306), .ZN(n2957) );
  XNOR2_X2 U2233 ( .A(n441), .B(n306), .ZN(n2958) );
  OAI22_X2 U2234 ( .A1(n401), .A2(n3152), .B1(n2992), .B2(n353), .ZN(n2016) );
  OAI22_X2 U2236 ( .A1(n401), .A2(n2962), .B1(n2961), .B2(n353), .ZN(n2436) );
  OAI22_X2 U2237 ( .A1(n401), .A2(n2963), .B1(n2962), .B2(n353), .ZN(n2437) );
  OAI22_X2 U2238 ( .A1(n401), .A2(n2964), .B1(n2963), .B2(n353), .ZN(n2438) );
  OAI22_X2 U2239 ( .A1(n401), .A2(n2965), .B1(n2964), .B2(n353), .ZN(n2439) );
  OAI22_X2 U2240 ( .A1(n401), .A2(n2966), .B1(n2965), .B2(n353), .ZN(n2440) );
  OAI22_X2 U2241 ( .A1(n401), .A2(n2967), .B1(n2966), .B2(n353), .ZN(n2441) );
  OAI22_X2 U2242 ( .A1(n401), .A2(n2968), .B1(n2967), .B2(n353), .ZN(n2442) );
  OAI22_X2 U2243 ( .A1(n401), .A2(n2969), .B1(n2968), .B2(n353), .ZN(n2443) );
  OAI22_X2 U2244 ( .A1(n400), .A2(n2970), .B1(n2969), .B2(n352), .ZN(n2444) );
  OAI22_X2 U2245 ( .A1(n400), .A2(n2971), .B1(n2970), .B2(n352), .ZN(n2445) );
  OAI22_X2 U2246 ( .A1(n400), .A2(n2972), .B1(n2971), .B2(n352), .ZN(n2446) );
  OAI22_X2 U2247 ( .A1(n400), .A2(n2973), .B1(n2972), .B2(n352), .ZN(n2447) );
  OAI22_X2 U2248 ( .A1(n400), .A2(n2974), .B1(n2973), .B2(n352), .ZN(n2448) );
  OAI22_X2 U2249 ( .A1(n400), .A2(n2975), .B1(n2974), .B2(n352), .ZN(n2449) );
  OAI22_X2 U2250 ( .A1(n400), .A2(n2976), .B1(n2975), .B2(n352), .ZN(n2450) );
  OAI22_X2 U2251 ( .A1(n400), .A2(n2977), .B1(n2976), .B2(n352), .ZN(n2451) );
  OAI22_X2 U2252 ( .A1(n400), .A2(n2978), .B1(n2977), .B2(n352), .ZN(n2452) );
  OAI22_X2 U2253 ( .A1(n400), .A2(n2979), .B1(n2978), .B2(n352), .ZN(n2453) );
  OAI22_X2 U2254 ( .A1(n400), .A2(n2980), .B1(n2979), .B2(n352), .ZN(n2454) );
  OAI22_X2 U2255 ( .A1(n399), .A2(n2981), .B1(n2980), .B2(n352), .ZN(n2455) );
  OAI22_X2 U2256 ( .A1(n399), .A2(n2982), .B1(n2981), .B2(n351), .ZN(n2456) );
  OAI22_X2 U2257 ( .A1(n399), .A2(n2983), .B1(n2982), .B2(n351), .ZN(n2457) );
  OAI22_X2 U2258 ( .A1(n399), .A2(n2984), .B1(n2983), .B2(n351), .ZN(n2458) );
  OAI22_X2 U2259 ( .A1(n399), .A2(n2985), .B1(n2984), .B2(n351), .ZN(n2459) );
  OAI22_X2 U2260 ( .A1(n399), .A2(n2986), .B1(n2985), .B2(n351), .ZN(n2460) );
  OAI22_X2 U2261 ( .A1(n399), .A2(n2987), .B1(n2986), .B2(n351), .ZN(n2461) );
  OAI22_X2 U2262 ( .A1(n399), .A2(n2988), .B1(n2987), .B2(n351), .ZN(n2462) );
  OAI22_X2 U2263 ( .A1(n399), .A2(n2989), .B1(n2988), .B2(n351), .ZN(n2463) );
  OAI22_X2 U2264 ( .A1(n399), .A2(n2990), .B1(n2989), .B2(n351), .ZN(n2464) );
  OAI22_X2 U2265 ( .A1(n399), .A2(n2991), .B1(n2990), .B2(n351), .ZN(n2465) );
  XNOR2_X2 U2266 ( .A(n3059), .B(n305), .ZN(n2960) );
  XNOR2_X2 U2267 ( .A(n3060), .B(n305), .ZN(n2961) );
  XNOR2_X2 U2268 ( .A(n3061), .B(n305), .ZN(n2962) );
  XNOR2_X2 U2269 ( .A(n3062), .B(n305), .ZN(n2963) );
  XNOR2_X2 U2270 ( .A(n3063), .B(n305), .ZN(n2964) );
  XNOR2_X2 U2271 ( .A(n3064), .B(n305), .ZN(n2965) );
  XNOR2_X2 U2272 ( .A(n3065), .B(n305), .ZN(n2966) );
  XNOR2_X2 U2273 ( .A(n3066), .B(n305), .ZN(n2967) );
  XNOR2_X2 U2274 ( .A(n3067), .B(n305), .ZN(n2968) );
  XNOR2_X2 U2275 ( .A(n3068), .B(n305), .ZN(n2969) );
  XNOR2_X2 U2276 ( .A(n3069), .B(n305), .ZN(n2970) );
  XNOR2_X2 U2277 ( .A(n3070), .B(n304), .ZN(n2971) );
  XNOR2_X2 U2278 ( .A(n3071), .B(n304), .ZN(n2972) );
  XNOR2_X2 U2279 ( .A(n3072), .B(n304), .ZN(n2973) );
  XNOR2_X2 U2280 ( .A(n3073), .B(n304), .ZN(n2974) );
  XNOR2_X2 U2281 ( .A(n3074), .B(n304), .ZN(n2975) );
  XNOR2_X2 U2282 ( .A(n3075), .B(n304), .ZN(n2976) );
  XNOR2_X2 U2283 ( .A(n3076), .B(n304), .ZN(n2977) );
  XNOR2_X2 U2284 ( .A(n3077), .B(n304), .ZN(n2978) );
  XNOR2_X2 U2285 ( .A(n3078), .B(n304), .ZN(n2979) );
  XNOR2_X2 U2286 ( .A(n3079), .B(n304), .ZN(n2980) );
  XNOR2_X2 U2287 ( .A(n3080), .B(n304), .ZN(n2981) );
  XNOR2_X2 U2288 ( .A(n3081), .B(n304), .ZN(n2982) );
  XNOR2_X2 U2289 ( .A(n3082), .B(n303), .ZN(n2983) );
  XNOR2_X2 U2290 ( .A(n3083), .B(n303), .ZN(n2984) );
  XNOR2_X2 U2291 ( .A(n3084), .B(n303), .ZN(n2985) );
  XNOR2_X2 U2292 ( .A(n3085), .B(n303), .ZN(n2986) );
  XNOR2_X2 U2293 ( .A(n3086), .B(n303), .ZN(n2987) );
  XNOR2_X2 U2294 ( .A(n3087), .B(n303), .ZN(n2988) );
  XNOR2_X2 U2295 ( .A(n3088), .B(n303), .ZN(n2989) );
  XNOR2_X2 U2296 ( .A(n3089), .B(n303), .ZN(n2990) );
  XNOR2_X2 U2297 ( .A(n441), .B(n303), .ZN(n2991) );
  OAI22_X2 U2298 ( .A1(n398), .A2(n3153), .B1(n3025), .B2(n350), .ZN(n2017) );
  OAI22_X2 U2300 ( .A1(n398), .A2(n2995), .B1(n2994), .B2(n350), .ZN(n2468) );
  OAI22_X2 U2301 ( .A1(n398), .A2(n2996), .B1(n2995), .B2(n350), .ZN(n2469) );
  OAI22_X2 U2302 ( .A1(n398), .A2(n2997), .B1(n2996), .B2(n350), .ZN(n2470) );
  OAI22_X2 U2303 ( .A1(n398), .A2(n2998), .B1(n2997), .B2(n350), .ZN(n2471) );
  OAI22_X2 U2304 ( .A1(n398), .A2(n2999), .B1(n2998), .B2(n350), .ZN(n2472) );
  OAI22_X2 U2305 ( .A1(n398), .A2(n3000), .B1(n2999), .B2(n350), .ZN(n2473) );
  OAI22_X2 U2306 ( .A1(n398), .A2(n3001), .B1(n3000), .B2(n350), .ZN(n2474) );
  OAI22_X2 U2307 ( .A1(n398), .A2(n3002), .B1(n3001), .B2(n350), .ZN(n2475) );
  OAI22_X2 U2308 ( .A1(n397), .A2(n3003), .B1(n3002), .B2(n349), .ZN(n2476) );
  OAI22_X2 U2309 ( .A1(n397), .A2(n3004), .B1(n3003), .B2(n349), .ZN(n2477) );
  OAI22_X2 U2310 ( .A1(n397), .A2(n3005), .B1(n3004), .B2(n349), .ZN(n2478) );
  OAI22_X2 U2311 ( .A1(n397), .A2(n3006), .B1(n3005), .B2(n349), .ZN(n2479) );
  OAI22_X2 U2312 ( .A1(n397), .A2(n3007), .B1(n3006), .B2(n349), .ZN(n2480) );
  OAI22_X2 U2313 ( .A1(n397), .A2(n3008), .B1(n3007), .B2(n349), .ZN(n2481) );
  OAI22_X2 U2314 ( .A1(n397), .A2(n3009), .B1(n3008), .B2(n349), .ZN(n2482) );
  OAI22_X2 U2315 ( .A1(n397), .A2(n3010), .B1(n3009), .B2(n349), .ZN(n2483) );
  OAI22_X2 U2316 ( .A1(n397), .A2(n3011), .B1(n3010), .B2(n349), .ZN(n2484) );
  OAI22_X2 U2317 ( .A1(n397), .A2(n3012), .B1(n3011), .B2(n349), .ZN(n2485) );
  OAI22_X2 U2318 ( .A1(n397), .A2(n3013), .B1(n3012), .B2(n349), .ZN(n2486) );
  OAI22_X2 U2319 ( .A1(n396), .A2(n3014), .B1(n3013), .B2(n349), .ZN(n2487) );
  OAI22_X2 U2320 ( .A1(n396), .A2(n3015), .B1(n3014), .B2(n348), .ZN(n2488) );
  OAI22_X2 U2321 ( .A1(n396), .A2(n3016), .B1(n3015), .B2(n348), .ZN(n2489) );
  OAI22_X2 U2322 ( .A1(n396), .A2(n3017), .B1(n3016), .B2(n348), .ZN(n2490) );
  OAI22_X2 U2323 ( .A1(n396), .A2(n3018), .B1(n3017), .B2(n348), .ZN(n2491) );
  OAI22_X2 U2324 ( .A1(n396), .A2(n3019), .B1(n3018), .B2(n348), .ZN(n2492) );
  OAI22_X2 U2325 ( .A1(n396), .A2(n3020), .B1(n3019), .B2(n348), .ZN(n2493) );
  OAI22_X2 U2326 ( .A1(n396), .A2(n3021), .B1(n3020), .B2(n348), .ZN(n2494) );
  OAI22_X2 U2327 ( .A1(n396), .A2(n3022), .B1(n3021), .B2(n348), .ZN(n2495) );
  OAI22_X2 U2328 ( .A1(n396), .A2(n3023), .B1(n3022), .B2(n348), .ZN(n2496) );
  OAI22_X2 U2329 ( .A1(n396), .A2(n3024), .B1(n3023), .B2(n348), .ZN(n2497) );
  XNOR2_X2 U2330 ( .A(n3059), .B(n302), .ZN(n2993) );
  XNOR2_X2 U2331 ( .A(n3060), .B(n302), .ZN(n2994) );
  XNOR2_X2 U2332 ( .A(n3061), .B(n302), .ZN(n2995) );
  XNOR2_X2 U2333 ( .A(n3062), .B(n302), .ZN(n2996) );
  XNOR2_X2 U2334 ( .A(n3063), .B(n302), .ZN(n2997) );
  XNOR2_X2 U2335 ( .A(n3064), .B(n302), .ZN(n2998) );
  XNOR2_X2 U2336 ( .A(n3065), .B(n302), .ZN(n2999) );
  XNOR2_X2 U2337 ( .A(n3066), .B(n302), .ZN(n3000) );
  XNOR2_X2 U2338 ( .A(n3067), .B(n302), .ZN(n3001) );
  XNOR2_X2 U2339 ( .A(n3068), .B(n302), .ZN(n3002) );
  XNOR2_X2 U2340 ( .A(n3069), .B(n302), .ZN(n3003) );
  XNOR2_X2 U2341 ( .A(n3070), .B(n301), .ZN(n3004) );
  XNOR2_X2 U2342 ( .A(n3071), .B(n301), .ZN(n3005) );
  XNOR2_X2 U2343 ( .A(n3072), .B(n301), .ZN(n3006) );
  XNOR2_X2 U2344 ( .A(n3073), .B(n301), .ZN(n3007) );
  XNOR2_X2 U2345 ( .A(n3074), .B(n301), .ZN(n3008) );
  XNOR2_X2 U2346 ( .A(n3075), .B(n301), .ZN(n3009) );
  XNOR2_X2 U2347 ( .A(n3076), .B(n301), .ZN(n3010) );
  XNOR2_X2 U2348 ( .A(n3077), .B(n301), .ZN(n3011) );
  XNOR2_X2 U2349 ( .A(n3078), .B(n301), .ZN(n3012) );
  XNOR2_X2 U2350 ( .A(n3079), .B(n301), .ZN(n3013) );
  XNOR2_X2 U2351 ( .A(n3080), .B(n301), .ZN(n3014) );
  XNOR2_X2 U2352 ( .A(n3081), .B(n301), .ZN(n3015) );
  XNOR2_X2 U2353 ( .A(n3082), .B(n300), .ZN(n3016) );
  XNOR2_X2 U2354 ( .A(n3083), .B(n300), .ZN(n3017) );
  XNOR2_X2 U2355 ( .A(n3084), .B(n300), .ZN(n3018) );
  XNOR2_X2 U2356 ( .A(n3085), .B(n300), .ZN(n3019) );
  XNOR2_X2 U2357 ( .A(n3086), .B(n300), .ZN(n3020) );
  XNOR2_X2 U2358 ( .A(n3087), .B(n300), .ZN(n3021) );
  XNOR2_X2 U2359 ( .A(n3088), .B(n300), .ZN(n3022) );
  XNOR2_X2 U2360 ( .A(n3089), .B(n300), .ZN(n3023) );
  XNOR2_X2 U2361 ( .A(n441), .B(n300), .ZN(n3024) );
  OAI22_X2 U2362 ( .A1(n395), .A2(n3154), .B1(n3058), .B2(n347), .ZN(n2018) );
  OAI22_X2 U2363 ( .A1(n395), .A2(n3027), .B1(n3026), .B2(n347), .ZN(n2500) );
  OAI22_X2 U2364 ( .A1(n395), .A2(n3028), .B1(n3027), .B2(n347), .ZN(n2501) );
  OAI22_X2 U2365 ( .A1(n395), .A2(n3029), .B1(n3028), .B2(n347), .ZN(n2502) );
  OAI22_X2 U2366 ( .A1(n395), .A2(n3030), .B1(n3029), .B2(n347), .ZN(n2503) );
  OAI22_X2 U2367 ( .A1(n395), .A2(n3031), .B1(n3030), .B2(n347), .ZN(n2504) );
  OAI22_X2 U2368 ( .A1(n395), .A2(n3032), .B1(n3031), .B2(n347), .ZN(n2505) );
  OAI22_X2 U2369 ( .A1(n395), .A2(n3033), .B1(n3032), .B2(n347), .ZN(n2506) );
  OAI22_X2 U2370 ( .A1(n395), .A2(n3034), .B1(n3033), .B2(n347), .ZN(n2507) );
  OAI22_X2 U2371 ( .A1(n395), .A2(n3035), .B1(n3034), .B2(n347), .ZN(n2508) );
  OAI22_X2 U2372 ( .A1(n394), .A2(n3036), .B1(n3035), .B2(n346), .ZN(n2509) );
  OAI22_X2 U2373 ( .A1(n394), .A2(n3037), .B1(n3036), .B2(n346), .ZN(n2510) );
  OAI22_X2 U2374 ( .A1(n394), .A2(n3038), .B1(n3037), .B2(n346), .ZN(n2511) );
  OAI22_X2 U2375 ( .A1(n394), .A2(n3039), .B1(n3038), .B2(n346), .ZN(n2512) );
  OAI22_X2 U2376 ( .A1(n394), .A2(n3040), .B1(n3039), .B2(n346), .ZN(n2513) );
  OAI22_X2 U2377 ( .A1(n394), .A2(n3041), .B1(n3040), .B2(n346), .ZN(n2514) );
  OAI22_X2 U2378 ( .A1(n394), .A2(n3042), .B1(n3041), .B2(n346), .ZN(n2515) );
  OAI22_X2 U2379 ( .A1(n394), .A2(n3043), .B1(n3042), .B2(n346), .ZN(n2516) );
  OAI22_X2 U2380 ( .A1(n394), .A2(n3044), .B1(n3043), .B2(n346), .ZN(n2517) );
  OAI22_X2 U2381 ( .A1(n394), .A2(n3045), .B1(n3044), .B2(n346), .ZN(n2518) );
  OAI22_X2 U2382 ( .A1(n394), .A2(n3046), .B1(n3045), .B2(n346), .ZN(n2519) );
  OAI22_X2 U2383 ( .A1(n393), .A2(n3047), .B1(n3046), .B2(n346), .ZN(n2520) );
  OAI22_X2 U2384 ( .A1(n393), .A2(n3048), .B1(n3047), .B2(n345), .ZN(n2521) );
  OAI22_X2 U2385 ( .A1(n393), .A2(n3049), .B1(n3048), .B2(n345), .ZN(n2522) );
  OAI22_X2 U2386 ( .A1(n393), .A2(n3050), .B1(n3049), .B2(n345), .ZN(n2523) );
  OAI22_X2 U2387 ( .A1(n393), .A2(n3051), .B1(n3050), .B2(n345), .ZN(n2524) );
  OAI22_X2 U2388 ( .A1(n393), .A2(n3052), .B1(n3051), .B2(n345), .ZN(n2525) );
  OAI22_X2 U2389 ( .A1(n393), .A2(n3053), .B1(n3052), .B2(n345), .ZN(n2526) );
  OAI22_X2 U2390 ( .A1(n393), .A2(n3054), .B1(n3053), .B2(n345), .ZN(n2527) );
  OAI22_X2 U2391 ( .A1(n393), .A2(n3055), .B1(n3054), .B2(n345), .ZN(n2528) );
  OAI22_X2 U2392 ( .A1(n393), .A2(n3056), .B1(n3055), .B2(n345), .ZN(n2529) );
  OAI22_X2 U2393 ( .A1(n393), .A2(n3057), .B1(n3056), .B2(n345), .ZN(n2530) );
  XNOR2_X2 U2394 ( .A(n3059), .B(n299), .ZN(n3026) );
  XNOR2_X2 U2395 ( .A(n3060), .B(n299), .ZN(n3027) );
  XNOR2_X2 U2396 ( .A(n3061), .B(n299), .ZN(n3028) );
  XNOR2_X2 U2397 ( .A(n3062), .B(n299), .ZN(n3029) );
  XNOR2_X2 U2398 ( .A(n3063), .B(n299), .ZN(n3030) );
  XNOR2_X2 U2399 ( .A(n3064), .B(n299), .ZN(n3031) );
  XNOR2_X2 U2400 ( .A(n3065), .B(n299), .ZN(n3032) );
  XNOR2_X2 U2401 ( .A(n3066), .B(n299), .ZN(n3033) );
  XNOR2_X2 U2402 ( .A(n3067), .B(n299), .ZN(n3034) );
  XNOR2_X2 U2403 ( .A(n3068), .B(n299), .ZN(n3035) );
  XNOR2_X2 U2404 ( .A(n3069), .B(n299), .ZN(n3036) );
  XNOR2_X2 U2405 ( .A(n3070), .B(n298), .ZN(n3037) );
  XNOR2_X2 U2406 ( .A(n3071), .B(n298), .ZN(n3038) );
  XNOR2_X2 U2407 ( .A(n3072), .B(n298), .ZN(n3039) );
  XNOR2_X2 U2408 ( .A(n3073), .B(n298), .ZN(n3040) );
  XNOR2_X2 U2409 ( .A(n3074), .B(n298), .ZN(n3041) );
  XNOR2_X2 U2410 ( .A(n3075), .B(n298), .ZN(n3042) );
  XNOR2_X2 U2411 ( .A(n3076), .B(n298), .ZN(n3043) );
  XNOR2_X2 U2412 ( .A(n3077), .B(n298), .ZN(n3044) );
  XNOR2_X2 U2413 ( .A(n3078), .B(n298), .ZN(n3045) );
  XNOR2_X2 U2414 ( .A(n3079), .B(n298), .ZN(n3046) );
  XNOR2_X2 U2415 ( .A(n3080), .B(n298), .ZN(n3047) );
  XNOR2_X2 U2416 ( .A(n3081), .B(n298), .ZN(n3048) );
  XNOR2_X2 U2417 ( .A(n3082), .B(n297), .ZN(n3049) );
  XNOR2_X2 U2418 ( .A(n3083), .B(n297), .ZN(n3050) );
  XNOR2_X2 U2419 ( .A(n3084), .B(n297), .ZN(n3051) );
  XNOR2_X2 U2420 ( .A(n3085), .B(n297), .ZN(n3052) );
  XNOR2_X2 U2421 ( .A(n3086), .B(n297), .ZN(n3053) );
  XNOR2_X2 U2422 ( .A(n3087), .B(n297), .ZN(n3054) );
  XNOR2_X2 U2423 ( .A(n3088), .B(n297), .ZN(n3055) );
  XNOR2_X2 U2424 ( .A(n3089), .B(n297), .ZN(n3056) );
  XNOR2_X2 U2425 ( .A(n441), .B(n297), .ZN(n3057) );
  BUF_X4 U2426 ( .A(b[31]), .Z(n3059) );
  BUF_X4 U2427 ( .A(b[30]), .Z(n3060) );
  BUF_X4 U2428 ( .A(b[29]), .Z(n3061) );
  BUF_X4 U2429 ( .A(b[28]), .Z(n3062) );
  BUF_X4 U2430 ( .A(b[27]), .Z(n3063) );
  BUF_X4 U2431 ( .A(b[26]), .Z(n3064) );
  BUF_X4 U2432 ( .A(b[25]), .Z(n3065) );
  BUF_X4 U2433 ( .A(b[24]), .Z(n3066) );
  BUF_X4 U2434 ( .A(b[23]), .Z(n3067) );
  BUF_X4 U2435 ( .A(b[22]), .Z(n3068) );
  BUF_X4 U2436 ( .A(b[21]), .Z(n3069) );
  BUF_X4 U2437 ( .A(b[20]), .Z(n3070) );
  BUF_X4 U2438 ( .A(b[19]), .Z(n3071) );
  BUF_X4 U2439 ( .A(b[18]), .Z(n3072) );
  BUF_X4 U2440 ( .A(b[17]), .Z(n3073) );
  BUF_X4 U2441 ( .A(b[16]), .Z(n3074) );
  BUF_X4 U2442 ( .A(b[15]), .Z(n3075) );
  BUF_X4 U2443 ( .A(b[14]), .Z(n3076) );
  BUF_X4 U2444 ( .A(b[13]), .Z(n3077) );
  BUF_X4 U2445 ( .A(b[12]), .Z(n3078) );
  BUF_X4 U2446 ( .A(b[11]), .Z(n3079) );
  BUF_X4 U2447 ( .A(b[10]), .Z(n3080) );
  BUF_X4 U2448 ( .A(b[9]), .Z(n3081) );
  BUF_X4 U2449 ( .A(b[8]), .Z(n3082) );
  BUF_X4 U2450 ( .A(b[7]), .Z(n3083) );
  BUF_X4 U2451 ( .A(b[6]), .Z(n3084) );
  BUF_X4 U2452 ( .A(b[5]), .Z(n3085) );
  BUF_X4 U2453 ( .A(b[4]), .Z(n3086) );
  BUF_X4 U2454 ( .A(b[3]), .Z(n3087) );
  BUF_X4 U2455 ( .A(b[2]), .Z(n3088) );
  BUF_X4 U2456 ( .A(b[1]), .Z(n3089) );
  INV_X32 U2457 ( .A(n342), .ZN(n3139) );
  INV_X32 U2458 ( .A(n339), .ZN(n3140) );
  BUF_X4 U2459 ( .A(a[29]), .Z(n3156) );
  INV_X32 U2460 ( .A(n336), .ZN(n3141) );
  BUF_X4 U2461 ( .A(a[27]), .Z(n3157) );
  INV_X32 U2462 ( .A(n333), .ZN(n3142) );
  BUF_X4 U2463 ( .A(a[25]), .Z(n3158) );
  INV_X32 U2464 ( .A(n330), .ZN(n3143) );
  BUF_X4 U2465 ( .A(a[23]), .Z(n3159) );
  INV_X32 U2466 ( .A(n327), .ZN(n3144) );
  BUF_X4 U2467 ( .A(a[21]), .Z(n3160) );
  INV_X32 U2468 ( .A(n324), .ZN(n3145) );
  BUF_X4 U2469 ( .A(a[19]), .Z(n3161) );
  INV_X32 U2470 ( .A(n321), .ZN(n3146) );
  BUF_X4 U2471 ( .A(a[17]), .Z(n3162) );
  INV_X32 U2472 ( .A(n318), .ZN(n3147) );
  BUF_X4 U2473 ( .A(a[15]), .Z(n3163) );
  INV_X32 U2474 ( .A(n315), .ZN(n3148) );
  BUF_X4 U2475 ( .A(a[13]), .Z(n3164) );
  INV_X32 U2476 ( .A(n312), .ZN(n3149) );
  BUF_X4 U2477 ( .A(a[11]), .Z(n3165) );
  INV_X32 U2478 ( .A(n309), .ZN(n3150) );
  BUF_X4 U2479 ( .A(a[9]), .Z(n3166) );
  INV_X32 U2480 ( .A(n306), .ZN(n3151) );
  BUF_X4 U2481 ( .A(a[7]), .Z(n3167) );
  INV_X32 U2482 ( .A(n303), .ZN(n3152) );
  BUF_X4 U2483 ( .A(a[5]), .Z(n3168) );
  INV_X32 U2484 ( .A(n300), .ZN(n3153) );
  BUF_X4 U2485 ( .A(a[3]), .Z(n3169) );
  INV_X32 U2486 ( .A(n297), .ZN(n3154) );
  BUF_X4 U2487 ( .A(a[1]), .Z(n3170) );
  XOR2_X2 U2489 ( .A(a[30]), .B(a[31]), .Z(n3091) );
  XOR2_X2 U2492 ( .A(a[28]), .B(a[29]), .Z(n3092) );
  XOR2_X2 U2495 ( .A(a[26]), .B(a[27]), .Z(n3093) );
  XOR2_X2 U2498 ( .A(a[24]), .B(a[25]), .Z(n3094) );
  XOR2_X2 U2501 ( .A(a[22]), .B(a[23]), .Z(n3095) );
  XOR2_X2 U2504 ( .A(a[20]), .B(a[21]), .Z(n3096) );
  XOR2_X2 U2507 ( .A(a[18]), .B(a[19]), .Z(n3097) );
  XOR2_X2 U2510 ( .A(a[16]), .B(a[17]), .Z(n3098) );
  XOR2_X2 U2513 ( .A(a[14]), .B(a[15]), .Z(n3099) );
  XOR2_X2 U2516 ( .A(a[12]), .B(a[13]), .Z(n3100) );
  XOR2_X2 U2519 ( .A(a[10]), .B(a[11]), .Z(n3101) );
  XOR2_X2 U2522 ( .A(a[8]), .B(a[9]), .Z(n3102) );
  XOR2_X2 U2525 ( .A(a[6]), .B(a[7]), .Z(n3103) );
  XOR2_X2 U2528 ( .A(a[4]), .B(a[5]), .Z(n3104) );
  XOR2_X2 U2531 ( .A(a[2]), .B(a[3]), .Z(n3105) );
  NAND2_X4 U2533 ( .A1(n3106), .A2(n3138), .ZN(n3122) );
  XOR2_X2 U2534 ( .A(a[0]), .B(a[1]), .Z(n3106) );
  INV_X32 U2535 ( .A(a[0]), .ZN(n3138) );
  OAI22_X4 U2538 ( .A1(n431), .A2(n2631), .B1(n2630), .B2(n383), .ZN(n1103) );
  BUF_X1 U2539 ( .A(n3110), .Z(n431) );
  OAI22_X4 U2540 ( .A1(n416), .A2(n2796), .B1(n2795), .B2(n368), .ZN(n1233) );
  BUF_X1 U2541 ( .A(n3115), .Z(n416) );
  OAI22_X4 U2542 ( .A1(n413), .A2(n2829), .B1(n2828), .B2(n365), .ZN(n1271) );
  BUF_X1 U2543 ( .A(n3116), .Z(n413) );
  OAI22_X4 U2544 ( .A1(n404), .A2(n2928), .B1(n2927), .B2(n356), .ZN(n1409) );
  BUF_X1 U2545 ( .A(n3119), .Z(n404) );
  OAI22_X4 U2546 ( .A1(n410), .A2(n2862), .B1(n2861), .B2(n362), .ZN(n1313) );
  BUF_X1 U2547 ( .A(n3117), .Z(n410) );
  OAI22_X4 U2548 ( .A1(n437), .A2(n2565), .B1(n2564), .B2(n389), .ZN(n1079) );
  BUF_X1 U2549 ( .A(n3108), .Z(n437) );
  OAI22_X4 U2550 ( .A1(n434), .A2(n2598), .B1(n2597), .B2(n386), .ZN(n1089) );
  BUF_X1 U2551 ( .A(n3109), .Z(n434) );
  OAI22_X4 U2552 ( .A1(n428), .A2(n2664), .B1(n2663), .B2(n380), .ZN(n1121) );
  BUF_X1 U2553 ( .A(n3111), .Z(n428) );
  OAI22_X4 U2554 ( .A1(n401), .A2(n2961), .B1(n2960), .B2(n353), .ZN(n1463) );
  BUF_X1 U2555 ( .A(n3120), .Z(n401) );
  OAI22_X4 U2556 ( .A1(n422), .A2(n2730), .B1(n2729), .B2(n374), .ZN(n1169) );
  BUF_X1 U2557 ( .A(n3113), .Z(n422) );
  OAI22_X4 U2558 ( .A1(n419), .A2(n2763), .B1(n2762), .B2(n371), .ZN(n1199) );
  BUF_X1 U2559 ( .A(n3114), .Z(n419) );
  OAI22_X4 U2560 ( .A1(n398), .A2(n2994), .B1(n2993), .B2(n350), .ZN(n1521) );
  BUF_X1 U2561 ( .A(n3121), .Z(n398) );
  OAI22_X4 U2562 ( .A1(n425), .A2(n2697), .B1(n2696), .B2(n377), .ZN(n1143) );
  BUF_X1 U2563 ( .A(n3112), .Z(n425) );
  OAI22_X4 U2564 ( .A1(n407), .A2(n2895), .B1(n2894), .B2(n359), .ZN(n1359) );
  BUF_X1 U2565 ( .A(n3118), .Z(n407) );
  OAI22_X4 U2566 ( .A1(n440), .A2(n2532), .B1(n2531), .B2(n392), .ZN(n1073) );
  BUF_X1 U2567 ( .A(n3107), .Z(n440) );
  BUF_X1 U2568 ( .A(n3129), .Z(n372) );
  BUF_X1 U2569 ( .A(n3129), .Z(n373) );
  BUF_X1 U2570 ( .A(n3129), .Z(n374) );
  NAND2_X2 U2571 ( .A1(n3097), .A2(n3129), .ZN(n3113) );
  XNOR2_X1 U2572 ( .A(a[18]), .B(a[17]), .ZN(n3129) );
  BUF_X1 U2573 ( .A(n3133), .Z(n360) );
  BUF_X1 U2574 ( .A(n3133), .Z(n361) );
  BUF_X1 U2575 ( .A(n3133), .Z(n362) );
  NAND2_X2 U2576 ( .A1(n3101), .A2(n3133), .ZN(n3117) );
  XNOR2_X1 U2577 ( .A(a[10]), .B(a[9]), .ZN(n3133) );
  BUF_X1 U2578 ( .A(n3128), .Z(n375) );
  BUF_X1 U2579 ( .A(n3128), .Z(n376) );
  BUF_X1 U2580 ( .A(n3128), .Z(n377) );
  NAND2_X2 U2581 ( .A1(n3096), .A2(n3128), .ZN(n3112) );
  XNOR2_X1 U2582 ( .A(a[20]), .B(a[19]), .ZN(n3128) );
  BUF_X1 U2583 ( .A(n3132), .Z(n363) );
  BUF_X1 U2584 ( .A(n3132), .Z(n364) );
  BUF_X1 U2585 ( .A(n3132), .Z(n365) );
  NAND2_X2 U2586 ( .A1(n3100), .A2(n3132), .ZN(n3116) );
  XNOR2_X1 U2587 ( .A(a[12]), .B(a[11]), .ZN(n3132) );
  BUF_X1 U2588 ( .A(n3131), .Z(n366) );
  BUF_X1 U2589 ( .A(n3131), .Z(n367) );
  BUF_X1 U2590 ( .A(n3131), .Z(n368) );
  NAND2_X2 U2591 ( .A1(n3099), .A2(n3131), .ZN(n3115) );
  XNOR2_X1 U2592 ( .A(a[14]), .B(a[13]), .ZN(n3131) );
  BUF_X1 U2593 ( .A(n3130), .Z(n369) );
  BUF_X1 U2594 ( .A(n3130), .Z(n370) );
  BUF_X1 U2595 ( .A(n3130), .Z(n371) );
  NAND2_X2 U2596 ( .A1(n3098), .A2(n3130), .ZN(n3114) );
  XNOR2_X1 U2597 ( .A(a[16]), .B(a[15]), .ZN(n3130) );
  BUF_X1 U2598 ( .A(n3127), .Z(n378) );
  BUF_X1 U2599 ( .A(n3127), .Z(n379) );
  BUF_X1 U2600 ( .A(n3127), .Z(n380) );
  NAND2_X2 U2601 ( .A1(n3095), .A2(n3127), .ZN(n3111) );
  XNOR2_X1 U2602 ( .A(a[22]), .B(a[21]), .ZN(n3127) );
  BUF_X1 U2603 ( .A(n3125), .Z(n384) );
  BUF_X1 U2604 ( .A(n3125), .Z(n385) );
  BUF_X1 U2605 ( .A(n3125), .Z(n386) );
  NAND2_X2 U2606 ( .A1(n3093), .A2(n3125), .ZN(n3109) );
  XNOR2_X1 U2607 ( .A(a[26]), .B(a[25]), .ZN(n3125) );
  BUF_X1 U2608 ( .A(n3126), .Z(n381) );
  BUF_X1 U2609 ( .A(n3126), .Z(n382) );
  BUF_X1 U2610 ( .A(n3126), .Z(n383) );
  NAND2_X2 U2611 ( .A1(n3094), .A2(n3126), .ZN(n3110) );
  XNOR2_X1 U2612 ( .A(a[24]), .B(a[23]), .ZN(n3126) );
  BUF_X1 U2613 ( .A(n3124), .Z(n389) );
  BUF_X1 U2614 ( .A(n3124), .Z(n388) );
  BUF_X1 U2615 ( .A(n3124), .Z(n387) );
  NAND2_X2 U2616 ( .A1(n3092), .A2(n3124), .ZN(n3108) );
  XNOR2_X1 U2617 ( .A(a[28]), .B(a[27]), .ZN(n3124) );
  BUF_X1 U2618 ( .A(n3137), .Z(n350) );
  BUF_X1 U2619 ( .A(n3137), .Z(n348) );
  BUF_X1 U2620 ( .A(n3137), .Z(n349) );
  NAND2_X2 U2621 ( .A1(n3105), .A2(n3137), .ZN(n3121) );
  XNOR2_X1 U2622 ( .A(a[2]), .B(a[1]), .ZN(n3137) );
  BUF_X1 U2623 ( .A(n3136), .Z(n351) );
  BUF_X1 U2624 ( .A(n3136), .Z(n352) );
  BUF_X1 U2625 ( .A(n3136), .Z(n353) );
  NAND2_X2 U2626 ( .A1(n3104), .A2(n3136), .ZN(n3120) );
  XNOR2_X1 U2627 ( .A(a[4]), .B(a[3]), .ZN(n3136) );
  BUF_X1 U2628 ( .A(n3135), .Z(n354) );
  BUF_X1 U2629 ( .A(n3135), .Z(n355) );
  BUF_X1 U2630 ( .A(n3135), .Z(n356) );
  NAND2_X2 U2631 ( .A1(n3103), .A2(n3135), .ZN(n3119) );
  XNOR2_X1 U2632 ( .A(a[6]), .B(a[5]), .ZN(n3135) );
  BUF_X1 U2633 ( .A(n3134), .Z(n357) );
  BUF_X1 U2634 ( .A(n3134), .Z(n358) );
  BUF_X1 U2635 ( .A(n3134), .Z(n359) );
  NAND2_X2 U2636 ( .A1(n3102), .A2(n3134), .ZN(n3118) );
  XNOR2_X1 U2637 ( .A(a[8]), .B(a[7]), .ZN(n3134) );
  BUF_X1 U2638 ( .A(n3123), .Z(n390) );
  BUF_X1 U2639 ( .A(n3123), .Z(n391) );
  BUF_X1 U2640 ( .A(n3123), .Z(n392) );
  NAND2_X2 U2641 ( .A1(n3091), .A2(n3123), .ZN(n3107) );
  XNOR2_X1 U2642 ( .A(a[30]), .B(a[29]), .ZN(n3123) );
endmodule


module up_island_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[26] ,
         \carry[23] , \carry[22] , \carry[21] , \carry[20] , \carry[19] ,
         \carry[18] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[4] ,
         \carry[3] , \carry[2] , \carry[1] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163;

  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  NAND2_X1 U1 ( .A1(A[12]), .A2(B[12]), .ZN(n49) );
  NAND2_X1 U2 ( .A1(A[6]), .A2(B[6]), .ZN(n158) );
  INV_X1 U3 ( .A(n44), .ZN(n38) );
  INV_X1 U4 ( .A(n123), .ZN(n50) );
  INV_X1 U5 ( .A(n108), .ZN(n99) );
  INV_X1 U6 ( .A(n136), .ZN(n51) );
  NAND3_X2 U7 ( .A1(n91), .A2(n93), .A3(n92), .ZN(\carry[16] ) );
  NAND3_X2 U8 ( .A1(n40), .A2(n42), .A3(n41), .ZN(\carry[12] ) );
  NAND3_X2 U9 ( .A1(n111), .A2(n113), .A3(n112), .ZN(\carry[29] ) );
  NAND3_X2 U10 ( .A1(n47), .A2(n49), .A3(n48), .ZN(\carry[13] ) );
  BUF_X1 U11 ( .A(n141), .Z(n1) );
  NAND3_X2 U12 ( .A1(n54), .A2(n56), .A3(n55), .ZN(\carry[14] ) );
  BUF_X1 U13 ( .A(n77), .Z(n2) );
  XNOR2_X1 U14 ( .A(\carry[29] ), .B(n3), .ZN(SUM[29]) );
  XNOR2_X1 U15 ( .A(A[29]), .B(B[29]), .ZN(n3) );
  BUF_X1 U16 ( .A(n5), .Z(n4) );
  NAND3_X1 U17 ( .A1(n21), .A2(n23), .A3(n22), .ZN(n5) );
  NAND3_X1 U18 ( .A1(n21), .A2(n23), .A3(n22), .ZN(\carry[2] ) );
  BUF_X1 U19 ( .A(n109), .Z(n6) );
  NAND2_X1 U20 ( .A1(n66), .A2(A[6]), .ZN(n7) );
  NAND3_X1 U21 ( .A1(n159), .A2(n158), .A3(n7), .ZN(n8) );
  NAND3_X1 U22 ( .A1(n73), .A2(n75), .A3(n74), .ZN(\carry[15] ) );
  NAND3_X1 U23 ( .A1(n7), .A2(n159), .A3(n158), .ZN(\carry[7] ) );
  NAND2_X1 U24 ( .A1(n10), .A2(B[5]), .ZN(n9) );
  NAND3_X1 U25 ( .A1(n87), .A2(n88), .A3(n86), .ZN(n10) );
  AND3_X1 U26 ( .A1(n145), .A2(n147), .A3(n146), .ZN(n11) );
  NAND3_X1 U27 ( .A1(n87), .A2(n88), .A3(n86), .ZN(\carry[5] ) );
  NAND3_X1 U28 ( .A1(n27), .A2(n29), .A3(n28), .ZN(n12) );
  NAND3_X1 U29 ( .A1(n1), .A2(n143), .A3(n142), .ZN(n13) );
  NAND2_X1 U30 ( .A1(\carry[29] ), .A2(A[29]), .ZN(n14) );
  NAND3_X1 U31 ( .A1(n141), .A2(n143), .A3(n142), .ZN(n131) );
  BUF_X1 U32 ( .A(n101), .Z(n15) );
  BUF_X1 U33 ( .A(n119), .Z(n16) );
  BUF_X1 U34 ( .A(n105), .Z(n17) );
  NAND3_X1 U35 ( .A1(n68), .A2(n70), .A3(n69), .ZN(n18) );
  AND2_X2 U36 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
  BUF_X1 U37 ( .A(n106), .Z(n19) );
  XOR2_X1 U38 ( .A(B[1]), .B(A[1]), .Z(n20) );
  XOR2_X1 U39 ( .A(\carry[1] ), .B(n20), .Z(SUM[1]) );
  NAND2_X1 U40 ( .A1(\carry[1] ), .A2(B[1]), .ZN(n21) );
  NAND2_X1 U41 ( .A1(\carry[1] ), .A2(A[1]), .ZN(n22) );
  NAND2_X1 U42 ( .A1(B[1]), .A2(A[1]), .ZN(n23) );
  NAND2_X1 U43 ( .A1(\carry[29] ), .A2(A[29]), .ZN(n59) );
  NAND2_X1 U44 ( .A1(n10), .A2(A[5]), .ZN(n24) );
  BUF_X1 U45 ( .A(n125), .Z(n25) );
  XOR2_X1 U46 ( .A(B[2]), .B(A[2]), .Z(n26) );
  XOR2_X1 U47 ( .A(n4), .B(n26), .Z(SUM[2]) );
  NAND2_X1 U48 ( .A1(n5), .A2(B[2]), .ZN(n27) );
  NAND2_X1 U49 ( .A1(\carry[2] ), .A2(A[2]), .ZN(n28) );
  NAND2_X1 U50 ( .A1(B[2]), .A2(A[2]), .ZN(n29) );
  NAND3_X1 U51 ( .A1(n27), .A2(n29), .A3(n28), .ZN(\carry[3] ) );
  NAND3_X1 U52 ( .A1(n14), .A2(n58), .A3(n60), .ZN(n30) );
  NAND3_X1 U53 ( .A1(n59), .A2(n58), .A3(n60), .ZN(\carry[30] ) );
  NAND2_X1 U54 ( .A1(\carry[26] ), .A2(B[26]), .ZN(n125) );
  BUF_X1 U55 ( .A(n8), .Z(n31) );
  BUF_X1 U56 ( .A(n12), .Z(n32) );
  BUF_X1 U57 ( .A(\carry[11] ), .Z(n33) );
  BUF_X1 U58 ( .A(\carry[13] ), .Z(n34) );
  BUF_X1 U59 ( .A(\carry[14] ), .Z(n35) );
  BUF_X1 U60 ( .A(\carry[12] ), .Z(n36) );
  INV_X1 U61 ( .A(n11), .ZN(n37) );
  XNOR2_X1 U62 ( .A(n43), .B(n38), .ZN(SUM[28]) );
  XOR2_X1 U63 ( .A(A[11]), .B(B[11]), .Z(n39) );
  XOR2_X1 U64 ( .A(n33), .B(n39), .Z(SUM[11]) );
  NAND2_X1 U65 ( .A1(\carry[11] ), .A2(A[11]), .ZN(n40) );
  NAND2_X1 U66 ( .A1(\carry[11] ), .A2(B[11]), .ZN(n41) );
  NAND2_X1 U67 ( .A1(A[11]), .A2(B[11]), .ZN(n42) );
  AND3_X1 U68 ( .A1(n137), .A2(n139), .A3(n138), .ZN(n43) );
  XNOR2_X1 U69 ( .A(A[28]), .B(B[28]), .ZN(n44) );
  NAND2_X1 U70 ( .A1(n37), .A2(A[26]), .ZN(n45) );
  XOR2_X1 U71 ( .A(A[12]), .B(B[12]), .Z(n46) );
  XOR2_X1 U72 ( .A(n36), .B(n46), .Z(SUM[12]) );
  NAND2_X1 U73 ( .A1(\carry[12] ), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U74 ( .A1(\carry[12] ), .A2(B[12]), .ZN(n48) );
  XNOR2_X1 U75 ( .A(n52), .B(n50), .ZN(SUM[26]) );
  XNOR2_X1 U76 ( .A(n96), .B(n51), .ZN(SUM[27]) );
  BUF_X1 U77 ( .A(n37), .Z(n52) );
  XOR2_X1 U78 ( .A(A[13]), .B(B[13]), .Z(n53) );
  XOR2_X1 U79 ( .A(n34), .B(n53), .Z(SUM[13]) );
  NAND2_X1 U80 ( .A1(\carry[13] ), .A2(A[13]), .ZN(n54) );
  NAND2_X1 U81 ( .A1(\carry[13] ), .A2(B[13]), .ZN(n55) );
  NAND2_X1 U82 ( .A1(A[13]), .A2(B[13]), .ZN(n56) );
  BUF_X1 U83 ( .A(n18), .Z(n57) );
  NAND2_X1 U84 ( .A1(A[29]), .A2(B[29]), .ZN(n58) );
  NAND2_X1 U85 ( .A1(B[29]), .A2(n65), .ZN(n60) );
  XOR2_X1 U86 ( .A(A[30]), .B(B[30]), .Z(n61) );
  XOR2_X1 U87 ( .A(n30), .B(n61), .Z(SUM[30]) );
  NAND2_X1 U88 ( .A1(A[30]), .A2(B[30]), .ZN(n62) );
  NAND2_X1 U89 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n63) );
  NAND2_X1 U90 ( .A1(\carry[30] ), .A2(B[30]), .ZN(n64) );
  NAND3_X1 U91 ( .A1(n63), .A2(n64), .A3(n62), .ZN(\carry[31] ) );
  NAND3_X1 U92 ( .A1(n111), .A2(n113), .A3(n112), .ZN(n65) );
  NAND3_X1 U93 ( .A1(n128), .A2(n130), .A3(n129), .ZN(n66) );
  XOR2_X1 U94 ( .A(A[3]), .B(B[3]), .Z(n67) );
  XOR2_X1 U95 ( .A(n32), .B(n67), .Z(SUM[3]) );
  NAND2_X1 U96 ( .A1(n12), .A2(A[3]), .ZN(n68) );
  NAND2_X1 U97 ( .A1(\carry[3] ), .A2(B[3]), .ZN(n69) );
  NAND2_X1 U98 ( .A1(A[3]), .A2(B[3]), .ZN(n70) );
  NAND3_X1 U99 ( .A1(n68), .A2(n70), .A3(n69), .ZN(\carry[4] ) );
  BUF_X1 U100 ( .A(\carry[15] ), .Z(n71) );
  XOR2_X1 U101 ( .A(A[14]), .B(B[14]), .Z(n72) );
  XOR2_X1 U102 ( .A(n35), .B(n72), .Z(SUM[14]) );
  NAND2_X1 U103 ( .A1(\carry[14] ), .A2(A[14]), .ZN(n73) );
  NAND2_X1 U104 ( .A1(\carry[14] ), .A2(B[14]), .ZN(n74) );
  NAND2_X1 U105 ( .A1(A[14]), .A2(B[14]), .ZN(n75) );
  BUF_X1 U106 ( .A(\carry[21] ), .Z(n76) );
  NAND3_X1 U107 ( .A1(n82), .A2(n84), .A3(n83), .ZN(n77) );
  BUF_X1 U108 ( .A(n10), .Z(n78) );
  NAND3_X1 U109 ( .A1(n115), .A2(n117), .A3(n116), .ZN(n79) );
  NAND3_X1 U110 ( .A1(n16), .A2(n121), .A3(n120), .ZN(n80) );
  XOR2_X1 U111 ( .A(A[21]), .B(B[21]), .Z(n81) );
  XOR2_X1 U112 ( .A(n76), .B(n81), .Z(SUM[21]) );
  NAND2_X1 U113 ( .A1(\carry[21] ), .A2(A[21]), .ZN(n82) );
  NAND2_X1 U114 ( .A1(\carry[21] ), .A2(B[21]), .ZN(n83) );
  NAND2_X1 U115 ( .A1(A[21]), .A2(B[21]), .ZN(n84) );
  NAND3_X1 U116 ( .A1(n82), .A2(n84), .A3(n83), .ZN(\carry[22] ) );
  XOR2_X1 U117 ( .A(B[4]), .B(A[4]), .Z(n85) );
  XOR2_X1 U118 ( .A(n57), .B(n85), .Z(SUM[4]) );
  NAND2_X1 U119 ( .A1(\carry[4] ), .A2(B[4]), .ZN(n86) );
  NAND2_X1 U120 ( .A1(n18), .A2(A[4]), .ZN(n87) );
  NAND2_X1 U121 ( .A1(B[4]), .A2(A[4]), .ZN(n88) );
  NAND3_X1 U122 ( .A1(n17), .A2(n107), .A3(n19), .ZN(n89) );
  XOR2_X1 U123 ( .A(A[15]), .B(B[15]), .Z(n90) );
  XOR2_X1 U124 ( .A(n71), .B(n90), .Z(SUM[15]) );
  NAND2_X1 U125 ( .A1(\carry[15] ), .A2(A[15]), .ZN(n91) );
  NAND2_X1 U126 ( .A1(\carry[15] ), .A2(B[15]), .ZN(n92) );
  NAND2_X1 U127 ( .A1(A[15]), .A2(B[15]), .ZN(n93) );
  BUF_X1 U128 ( .A(\carry[16] ), .Z(n94) );
  NAND2_X1 U129 ( .A1(\carry[26] ), .A2(A[26]), .ZN(n124) );
  NAND3_X1 U130 ( .A1(n45), .A2(n126), .A3(n25), .ZN(n96) );
  NAND3_X1 U131 ( .A1(n125), .A2(n126), .A3(n124), .ZN(n95) );
  BUF_X1 U132 ( .A(n66), .Z(n97) );
  NAND3_X1 U133 ( .A1(n15), .A2(n103), .A3(n102), .ZN(n98) );
  XNOR2_X1 U134 ( .A(\carry[31] ), .B(n99), .ZN(SUM[31]) );
  XOR2_X1 U135 ( .A(A[22]), .B(B[22]), .Z(n100) );
  XOR2_X1 U136 ( .A(n2), .B(n100), .Z(SUM[22]) );
  NAND2_X1 U137 ( .A1(n77), .A2(A[22]), .ZN(n101) );
  NAND2_X1 U138 ( .A1(\carry[22] ), .A2(B[22]), .ZN(n102) );
  NAND2_X1 U139 ( .A1(A[22]), .A2(B[22]), .ZN(n103) );
  NAND3_X1 U140 ( .A1(n101), .A2(n103), .A3(n102), .ZN(\carry[23] ) );
  XOR2_X1 U141 ( .A(A[16]), .B(B[16]), .Z(n104) );
  XOR2_X1 U142 ( .A(n94), .B(n104), .Z(SUM[16]) );
  NAND2_X1 U143 ( .A1(\carry[16] ), .A2(A[16]), .ZN(n105) );
  NAND2_X1 U144 ( .A1(\carry[16] ), .A2(B[16]), .ZN(n106) );
  NAND2_X1 U145 ( .A1(A[16]), .A2(B[16]), .ZN(n107) );
  NAND3_X1 U146 ( .A1(n105), .A2(n107), .A3(n106), .ZN(\carry[17] ) );
  XOR2_X1 U147 ( .A(A[31]), .B(B[31]), .Z(n108) );
  NAND3_X1 U148 ( .A1(n115), .A2(n117), .A3(n116), .ZN(n109) );
  NAND3_X1 U149 ( .A1(n133), .A2(n135), .A3(n134), .ZN(n110) );
  NAND3_X1 U150 ( .A1(n145), .A2(n147), .A3(n146), .ZN(\carry[26] ) );
  NAND2_X1 U151 ( .A1(\carry[28] ), .A2(A[28]), .ZN(n111) );
  NAND2_X1 U152 ( .A1(\carry[28] ), .A2(B[28]), .ZN(n112) );
  NAND2_X1 U153 ( .A1(A[28]), .A2(B[28]), .ZN(n113) );
  XOR2_X1 U154 ( .A(A[23]), .B(B[23]), .Z(n114) );
  XOR2_X1 U155 ( .A(n98), .B(n114), .Z(SUM[23]) );
  NAND2_X1 U156 ( .A1(\carry[23] ), .A2(A[23]), .ZN(n115) );
  NAND2_X1 U157 ( .A1(\carry[23] ), .A2(B[23]), .ZN(n116) );
  NAND2_X1 U158 ( .A1(A[23]), .A2(B[23]), .ZN(n117) );
  XOR2_X1 U159 ( .A(A[17]), .B(B[17]), .Z(n118) );
  XOR2_X1 U160 ( .A(n89), .B(n118), .Z(SUM[17]) );
  NAND2_X1 U161 ( .A1(\carry[17] ), .A2(A[17]), .ZN(n119) );
  NAND2_X1 U162 ( .A1(\carry[17] ), .A2(B[17]), .ZN(n120) );
  NAND2_X1 U163 ( .A1(A[17]), .A2(B[17]), .ZN(n121) );
  NAND3_X1 U164 ( .A1(n119), .A2(n121), .A3(n120), .ZN(\carry[18] ) );
  NAND3_X1 U165 ( .A1(n150), .A2(n152), .A3(n151), .ZN(n122) );
  XOR2_X1 U166 ( .A(A[26]), .B(B[26]), .Z(n123) );
  NAND2_X1 U167 ( .A1(A[26]), .A2(B[26]), .ZN(n126) );
  XOR2_X1 U168 ( .A(A[5]), .B(B[5]), .Z(n127) );
  XOR2_X1 U169 ( .A(n78), .B(n127), .Z(SUM[5]) );
  NAND2_X1 U170 ( .A1(\carry[5] ), .A2(A[5]), .ZN(n128) );
  NAND2_X1 U171 ( .A1(\carry[5] ), .A2(B[5]), .ZN(n129) );
  NAND2_X1 U172 ( .A1(A[5]), .A2(B[5]), .ZN(n130) );
  NAND3_X1 U173 ( .A1(n24), .A2(n130), .A3(n9), .ZN(\carry[6] ) );
  XOR2_X1 U174 ( .A(A[18]), .B(B[18]), .Z(n132) );
  XOR2_X1 U175 ( .A(n80), .B(n132), .Z(SUM[18]) );
  NAND2_X1 U176 ( .A1(\carry[18] ), .A2(A[18]), .ZN(n133) );
  NAND2_X1 U177 ( .A1(\carry[18] ), .A2(B[18]), .ZN(n134) );
  NAND2_X1 U178 ( .A1(A[18]), .A2(B[18]), .ZN(n135) );
  NAND3_X1 U179 ( .A1(n133), .A2(n135), .A3(n134), .ZN(\carry[19] ) );
  XOR2_X1 U180 ( .A(A[27]), .B(B[27]), .Z(n136) );
  NAND2_X1 U181 ( .A1(n95), .A2(A[27]), .ZN(n137) );
  NAND2_X1 U182 ( .A1(n95), .A2(B[27]), .ZN(n138) );
  NAND2_X1 U183 ( .A1(A[27]), .A2(B[27]), .ZN(n139) );
  NAND3_X1 U184 ( .A1(n137), .A2(n138), .A3(n139), .ZN(\carry[28] ) );
  XOR2_X1 U185 ( .A(A[24]), .B(B[24]), .Z(n140) );
  XOR2_X1 U186 ( .A(n6), .B(n140), .Z(SUM[24]) );
  NAND2_X1 U187 ( .A1(n79), .A2(A[24]), .ZN(n141) );
  NAND2_X1 U188 ( .A1(n109), .A2(B[24]), .ZN(n142) );
  NAND2_X1 U189 ( .A1(A[24]), .A2(B[24]), .ZN(n143) );
  XOR2_X1 U190 ( .A(A[25]), .B(B[25]), .Z(n144) );
  XOR2_X1 U191 ( .A(n13), .B(n144), .Z(SUM[25]) );
  NAND2_X1 U192 ( .A1(n131), .A2(A[25]), .ZN(n145) );
  NAND2_X1 U193 ( .A1(n131), .A2(B[25]), .ZN(n146) );
  NAND2_X1 U194 ( .A1(A[25]), .A2(B[25]), .ZN(n147) );
  BUF_X1 U195 ( .A(B[0]), .Z(n148) );
  XOR2_X1 U196 ( .A(A[19]), .B(B[19]), .Z(n149) );
  XOR2_X1 U197 ( .A(n110), .B(n149), .Z(SUM[19]) );
  NAND2_X1 U198 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n150) );
  NAND2_X1 U199 ( .A1(\carry[19] ), .A2(B[19]), .ZN(n151) );
  NAND2_X1 U200 ( .A1(A[19]), .A2(B[19]), .ZN(n152) );
  NAND3_X1 U201 ( .A1(n150), .A2(n152), .A3(n151), .ZN(\carry[20] ) );
  XOR2_X1 U202 ( .A(A[20]), .B(B[20]), .Z(n153) );
  XOR2_X1 U203 ( .A(n122), .B(n153), .Z(SUM[20]) );
  NAND2_X1 U204 ( .A1(\carry[20] ), .A2(A[20]), .ZN(n154) );
  NAND2_X1 U205 ( .A1(\carry[20] ), .A2(B[20]), .ZN(n155) );
  NAND2_X1 U206 ( .A1(A[20]), .A2(B[20]), .ZN(n156) );
  NAND3_X1 U207 ( .A1(n154), .A2(n156), .A3(n155), .ZN(\carry[21] ) );
  XOR2_X1 U208 ( .A(A[6]), .B(B[6]), .Z(n157) );
  XOR2_X1 U209 ( .A(n157), .B(n97), .Z(SUM[6]) );
  NAND2_X1 U210 ( .A1(B[6]), .A2(\carry[6] ), .ZN(n159) );
  XOR2_X1 U211 ( .A(A[7]), .B(B[7]), .Z(n160) );
  XOR2_X1 U212 ( .A(n160), .B(n31), .Z(SUM[7]) );
  NAND2_X1 U213 ( .A1(A[7]), .A2(B[7]), .ZN(n161) );
  NAND2_X1 U214 ( .A1(A[7]), .A2(\carry[7] ), .ZN(n162) );
  NAND2_X1 U215 ( .A1(n8), .A2(B[7]), .ZN(n163) );
  NAND3_X1 U216 ( .A1(n162), .A2(n163), .A3(n161), .ZN(\carry[8] ) );
  XOR2_X1 U217 ( .A(n148), .B(A[0]), .Z(SUM[0]) );
endmodule


module up_island_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] , \B_not[28] ,
         \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] , \B_not[23] ,
         \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] , \B_not[18] ,
         \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] , \B_not[13] ,
         \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] , \B_not[8] ,
         \B_not[7] , \B_not[6] , \B_not[5] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178;

  FA_X1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  FA_X1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  NAND2_X1 U1 ( .A1(\B_not[9] ), .A2(A[9]), .ZN(n109) );
  NAND2_X1 U2 ( .A1(\B_not[10] ), .A2(A[10]), .ZN(n113) );
  NAND2_X1 U3 ( .A1(A[22]), .A2(\B_not[22] ), .ZN(n34) );
  NAND2_X1 U4 ( .A1(\B_not[23] ), .A2(A[23]), .ZN(n169) );
  NAND2_X1 U5 ( .A1(\B_not[8] ), .A2(A[8]), .ZN(n160) );
  NAND2_X1 U6 ( .A1(\B_not[16] ), .A2(A[16]), .ZN(n80) );
  NAND2_X1 U7 ( .A1(\B_not[17] ), .A2(A[17]), .ZN(n173) );
  NAND2_X1 U8 ( .A1(\B_not[7] ), .A2(A[7]), .ZN(n164) );
  NAND2_X1 U9 ( .A1(\B_not[14] ), .A2(A[14]), .ZN(n156) );
  NAND2_X1 U10 ( .A1(\B_not[13] ), .A2(A[13]), .ZN(n148) );
  NAND2_X1 U11 ( .A1(\B_not[11] ), .A2(A[11]), .ZN(n105) );
  NAND2_X1 U12 ( .A1(\B_not[12] ), .A2(A[12]), .ZN(n140) );
  NAND2_X1 U13 ( .A1(A[24]), .A2(\B_not[24] ), .ZN(n123) );
  NAND2_X1 U14 ( .A1(\B_not[6] ), .A2(A[6]), .ZN(n144) );
  INV_X1 U15 ( .A(n118), .ZN(n72) );
  INV_X1 U16 ( .A(n134), .ZN(n46) );
  NAND2_X1 U17 ( .A1(n64), .A2(\B_not[12] ), .ZN(n1) );
  NAND2_X2 U18 ( .A1(n71), .A2(\B_not[24] ), .ZN(n125) );
  NAND2_X1 U19 ( .A1(\carry[24] ), .A2(A[24]), .ZN(n2) );
  NAND2_X1 U20 ( .A1(\carry[24] ), .A2(A[24]), .ZN(n124) );
  NAND3_X1 U21 ( .A1(n2), .A2(n123), .A3(n125), .ZN(n3) );
  BUF_X1 U22 ( .A(n2), .Z(n4) );
  BUF_X1 U23 ( .A(A[1]), .Z(n5) );
  NAND3_X2 U24 ( .A1(n163), .A2(n164), .A3(n162), .ZN(\carry[8] ) );
  NAND2_X1 U25 ( .A1(\carry[13] ), .A2(A[13]), .ZN(n147) );
  NAND3_X1 U26 ( .A1(n101), .A2(n102), .A3(n100), .ZN(\carry[6] ) );
  INV_X1 U27 ( .A(n165), .ZN(n6) );
  NAND2_X1 U28 ( .A1(\carry[11] ), .A2(A[11]), .ZN(n7) );
  NAND2_X1 U29 ( .A1(n29), .A2(\B_not[11] ), .ZN(n8) );
  NAND2_X2 U30 ( .A1(n87), .A2(\B_not[13] ), .ZN(n146) );
  NAND3_X2 U31 ( .A1(n108), .A2(n109), .A3(n107), .ZN(\carry[10] ) );
  NAND3_X1 U32 ( .A1(n159), .A2(n160), .A3(n158), .ZN(n9) );
  BUF_X1 U33 ( .A(n48), .Z(n10) );
  BUF_X1 U34 ( .A(n49), .Z(n11) );
  NAND2_X1 U35 ( .A1(n21), .A2(A[3]), .ZN(n12) );
  BUF_X1 U36 ( .A(n64), .Z(n13) );
  NAND3_X1 U37 ( .A1(n147), .A2(n148), .A3(n146), .ZN(n14) );
  BUF_X1 U38 ( .A(n90), .Z(n15) );
  NAND3_X1 U39 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n16) );
  BUF_X1 U40 ( .A(\carry[10] ), .Z(n17) );
  BUF_X1 U41 ( .A(n26), .Z(n18) );
  BUF_X1 U42 ( .A(n128), .Z(n19) );
  BUF_X1 U43 ( .A(\carry[19] ), .Z(n20) );
  NAND3_X2 U44 ( .A1(n32), .A2(n34), .A3(n33), .ZN(\carry[23] ) );
  NAND3_X1 U45 ( .A1(n159), .A2(n158), .A3(n160), .ZN(\carry[9] ) );
  NAND3_X1 U46 ( .A1(n132), .A2(n131), .A3(n133), .ZN(n21) );
  NAND3_X1 U47 ( .A1(n132), .A2(n131), .A3(n133), .ZN(\carry[3] ) );
  BUF_X1 U48 ( .A(n74), .Z(n22) );
  NAND2_X1 U49 ( .A1(n15), .A2(\B_not[25] ), .ZN(n23) );
  BUF_X1 U50 ( .A(n75), .Z(n24) );
  BUF_X1 U51 ( .A(\carry[24] ), .Z(n25) );
  NAND3_X1 U52 ( .A1(n92), .A2(n93), .A3(n94), .ZN(n26) );
  NAND3_X1 U53 ( .A1(n96), .A2(n97), .A3(n98), .ZN(n27) );
  NAND3_X1 U54 ( .A1(n92), .A2(n94), .A3(n93), .ZN(\carry[22] ) );
  NAND3_X2 U55 ( .A1(n58), .A2(n60), .A3(n59), .ZN(\carry[5] ) );
  NAND3_X1 U56 ( .A1(n12), .A2(n117), .A3(n115), .ZN(n28) );
  NAND3_X1 U57 ( .A1(n112), .A2(n113), .A3(n111), .ZN(n29) );
  BUF_X1 U58 ( .A(\carry[16] ), .Z(n30) );
  XOR2_X1 U59 ( .A(A[22]), .B(\B_not[22] ), .Z(n31) );
  XOR2_X1 U60 ( .A(n18), .B(n31), .Z(DIFF[22]) );
  NAND2_X1 U61 ( .A1(n26), .A2(A[22]), .ZN(n32) );
  NAND2_X1 U62 ( .A1(\carry[22] ), .A2(\B_not[22] ), .ZN(n33) );
  NAND3_X1 U63 ( .A1(n10), .A2(n50), .A3(n11), .ZN(n35) );
  INV_X4 U64 ( .A(B[22]), .ZN(\B_not[22] ) );
  AND3_X1 U65 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n40) );
  NAND2_X1 U66 ( .A1(n64), .A2(\B_not[12] ), .ZN(n36) );
  NAND3_X1 U67 ( .A1(n112), .A2(n111), .A3(n113), .ZN(\carry[11] ) );
  NAND2_X1 U68 ( .A1(\carry[10] ), .A2(\B_not[10] ), .ZN(n111) );
  XNOR2_X1 U69 ( .A(\carry[31] ), .B(n45), .ZN(DIFF[31]) );
  BUF_X1 U70 ( .A(\carry[23] ), .Z(n37) );
  BUF_X1 U71 ( .A(\carry[4] ), .Z(n38) );
  NAND3_X1 U72 ( .A1(n116), .A2(n117), .A3(n115), .ZN(\carry[4] ) );
  XNOR2_X1 U73 ( .A(n40), .B(n39), .ZN(DIFF[30]) );
  INV_X32 U74 ( .A(n46), .ZN(n39) );
  BUF_X1 U75 ( .A(n16), .Z(n41) );
  BUF_X1 U76 ( .A(n147), .Z(n42) );
  BUF_X1 U77 ( .A(n79), .Z(n43) );
  XNOR2_X1 U78 ( .A(n44), .B(n81), .ZN(DIFF[28]) );
  AND3_X1 U79 ( .A1(n119), .A2(n120), .A3(n121), .ZN(n44) );
  XNOR2_X1 U80 ( .A(A[31]), .B(\B_not[31] ), .ZN(n45) );
  XOR2_X1 U81 ( .A(A[19]), .B(\B_not[19] ), .Z(n47) );
  XOR2_X1 U82 ( .A(n20), .B(n47), .Z(DIFF[19]) );
  NAND2_X1 U83 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n48) );
  NAND2_X1 U84 ( .A1(\carry[19] ), .A2(\B_not[19] ), .ZN(n49) );
  NAND2_X1 U85 ( .A1(A[19]), .A2(\B_not[19] ), .ZN(n50) );
  NAND3_X1 U86 ( .A1(n48), .A2(n49), .A3(n50), .ZN(\carry[20] ) );
  BUF_X1 U87 ( .A(\carry[6] ), .Z(n51) );
  BUF_X1 U88 ( .A(\carry[5] ), .Z(n52) );
  NAND3_X1 U89 ( .A1(n19), .A2(n127), .A3(n23), .ZN(n53) );
  NAND3_X1 U90 ( .A1(n43), .A2(n80), .A3(n78), .ZN(n54) );
  BUF_X1 U91 ( .A(\carry[13] ), .Z(n55) );
  NAND3_X1 U92 ( .A1(n143), .A2(n144), .A3(n142), .ZN(n56) );
  XOR2_X1 U93 ( .A(A[4]), .B(n174), .Z(n57) );
  XOR2_X1 U94 ( .A(n38), .B(n57), .Z(DIFF[4]) );
  NAND2_X1 U95 ( .A1(\carry[4] ), .A2(A[4]), .ZN(n58) );
  NAND2_X1 U96 ( .A1(n28), .A2(n174), .ZN(n59) );
  NAND2_X1 U97 ( .A1(A[4]), .A2(n174), .ZN(n60) );
  NAND3_X1 U98 ( .A1(n82), .A2(n84), .A3(n83), .ZN(n61) );
  NAND3_X1 U99 ( .A1(n78), .A2(n80), .A3(n79), .ZN(\carry[17] ) );
  BUF_X1 U100 ( .A(\carry[9] ), .Z(n62) );
  BUF_X1 U101 ( .A(\carry[8] ), .Z(n63) );
  NAND3_X1 U102 ( .A1(n8), .A2(n105), .A3(n7), .ZN(n64) );
  BUF_X1 U103 ( .A(n29), .Z(n65) );
  XOR2_X1 U104 ( .A(A[26]), .B(\B_not[26] ), .Z(n66) );
  XOR2_X1 U105 ( .A(n53), .B(n66), .Z(DIFF[26]) );
  NAND2_X1 U106 ( .A1(\carry[26] ), .A2(A[26]), .ZN(n67) );
  NAND2_X1 U107 ( .A1(\carry[26] ), .A2(\B_not[26] ), .ZN(n68) );
  NAND2_X1 U108 ( .A1(A[26]), .A2(\B_not[26] ), .ZN(n69) );
  NAND3_X1 U109 ( .A1(n67), .A2(n69), .A3(n68), .ZN(\carry[27] ) );
  NAND3_X1 U110 ( .A1(n22), .A2(n76), .A3(n24), .ZN(n70) );
  NAND3_X1 U111 ( .A1(n167), .A2(n169), .A3(n168), .ZN(n71) );
  NAND3_X1 U112 ( .A1(n104), .A2(n105), .A3(n7), .ZN(\carry[12] ) );
  XNOR2_X1 U113 ( .A(n41), .B(n72), .ZN(DIFF[27]) );
  XOR2_X1 U114 ( .A(A[20]), .B(\B_not[20] ), .Z(n73) );
  XOR2_X1 U115 ( .A(n35), .B(n73), .Z(DIFF[20]) );
  NAND2_X1 U116 ( .A1(\carry[20] ), .A2(A[20]), .ZN(n74) );
  NAND2_X1 U117 ( .A1(\carry[20] ), .A2(\B_not[20] ), .ZN(n75) );
  NAND2_X1 U118 ( .A1(A[20]), .A2(\B_not[20] ), .ZN(n76) );
  NAND3_X1 U119 ( .A1(n74), .A2(n75), .A3(n76), .ZN(\carry[21] ) );
  XOR2_X1 U120 ( .A(\B_not[16] ), .B(A[16]), .Z(n77) );
  XOR2_X1 U121 ( .A(n30), .B(n77), .Z(DIFF[16]) );
  NAND2_X1 U122 ( .A1(\carry[16] ), .A2(\B_not[16] ), .ZN(n78) );
  NAND2_X1 U123 ( .A1(\carry[16] ), .A2(A[16]), .ZN(n79) );
  XOR2_X1 U124 ( .A(A[28]), .B(\B_not[28] ), .Z(n81) );
  NAND2_X1 U125 ( .A1(\carry[28] ), .A2(A[28]), .ZN(n82) );
  NAND2_X1 U126 ( .A1(\carry[28] ), .A2(\B_not[28] ), .ZN(n83) );
  NAND2_X1 U127 ( .A1(A[28]), .A2(\B_not[28] ), .ZN(n84) );
  NAND3_X1 U128 ( .A1(n82), .A2(n83), .A3(n84), .ZN(\carry[29] ) );
  BUF_X1 U129 ( .A(n27), .Z(n85) );
  BUF_X1 U130 ( .A(n21), .Z(n86) );
  NAND3_X1 U131 ( .A1(n139), .A2(n140), .A3(n1), .ZN(n87) );
  NAND3_X1 U132 ( .A1(n146), .A2(n148), .A3(n42), .ZN(n88) );
  BUF_X1 U133 ( .A(n56), .Z(n89) );
  NAND3_X1 U134 ( .A1(n4), .A2(n123), .A3(n125), .ZN(n90) );
  XOR2_X1 U135 ( .A(A[21]), .B(\B_not[21] ), .Z(n91) );
  XOR2_X1 U136 ( .A(n70), .B(n91), .Z(DIFF[21]) );
  NAND2_X1 U137 ( .A1(\carry[21] ), .A2(A[21]), .ZN(n92) );
  NAND2_X1 U138 ( .A1(\carry[21] ), .A2(\B_not[21] ), .ZN(n93) );
  NAND2_X1 U139 ( .A1(A[21]), .A2(\B_not[21] ), .ZN(n94) );
  XOR2_X1 U140 ( .A(n177), .B(n5), .Z(n95) );
  XOR2_X1 U141 ( .A(\carry[1] ), .B(n95), .Z(DIFF[1]) );
  NAND2_X1 U142 ( .A1(\carry[1] ), .A2(n177), .ZN(n96) );
  NAND2_X1 U143 ( .A1(\carry[1] ), .A2(A[1]), .ZN(n97) );
  NAND2_X1 U144 ( .A1(n177), .A2(A[1]), .ZN(n98) );
  NAND3_X1 U145 ( .A1(n97), .A2(n98), .A3(n96), .ZN(\carry[2] ) );
  NAND3_X1 U146 ( .A1(n36), .A2(n139), .A3(n140), .ZN(\carry[13] ) );
  NAND3_X1 U147 ( .A1(n147), .A2(n148), .A3(n146), .ZN(\carry[14] ) );
  NAND3_X1 U148 ( .A1(n143), .A2(n144), .A3(n142), .ZN(\carry[7] ) );
  NAND3_X1 U149 ( .A1(n124), .A2(n123), .A3(n125), .ZN(\carry[25] ) );
  INV_X8 U150 ( .A(B[21]), .ZN(\B_not[21] ) );
  OR2_X2 U151 ( .A1(n165), .A2(A[0]), .ZN(\carry[1] ) );
  NAND2_X1 U152 ( .A1(\carry[7] ), .A2(\B_not[7] ), .ZN(n162) );
  XOR2_X1 U153 ( .A(\B_not[5] ), .B(A[5]), .Z(n99) );
  XOR2_X1 U154 ( .A(n52), .B(n99), .Z(DIFF[5]) );
  NAND2_X1 U155 ( .A1(\carry[5] ), .A2(\B_not[5] ), .ZN(n100) );
  NAND2_X1 U156 ( .A1(\carry[5] ), .A2(A[5]), .ZN(n101) );
  NAND2_X1 U157 ( .A1(\B_not[5] ), .A2(A[5]), .ZN(n102) );
  XOR2_X1 U158 ( .A(\B_not[11] ), .B(A[11]), .Z(n103) );
  XOR2_X1 U159 ( .A(n65), .B(n103), .Z(DIFF[11]) );
  NAND2_X1 U160 ( .A1(n29), .A2(\B_not[11] ), .ZN(n104) );
  INV_X2 U161 ( .A(B[11]), .ZN(\B_not[11] ) );
  XOR2_X1 U162 ( .A(\B_not[9] ), .B(A[9]), .Z(n106) );
  XOR2_X1 U163 ( .A(n62), .B(n106), .Z(DIFF[9]) );
  NAND2_X1 U164 ( .A1(n9), .A2(\B_not[9] ), .ZN(n107) );
  NAND2_X1 U165 ( .A1(\carry[9] ), .A2(A[9]), .ZN(n108) );
  XOR2_X1 U166 ( .A(\B_not[10] ), .B(A[10]), .Z(n110) );
  XOR2_X1 U167 ( .A(n17), .B(n110), .Z(DIFF[10]) );
  NAND2_X1 U168 ( .A1(\carry[10] ), .A2(A[10]), .ZN(n112) );
  XOR2_X1 U169 ( .A(n175), .B(A[3]), .Z(n114) );
  XOR2_X1 U170 ( .A(n86), .B(n114), .Z(DIFF[3]) );
  NAND2_X1 U171 ( .A1(\carry[3] ), .A2(n175), .ZN(n115) );
  NAND2_X1 U172 ( .A1(n21), .A2(A[3]), .ZN(n116) );
  NAND2_X1 U173 ( .A1(n175), .A2(A[3]), .ZN(n117) );
  XOR2_X1 U174 ( .A(A[27]), .B(\B_not[27] ), .Z(n118) );
  NAND2_X1 U175 ( .A1(\carry[27] ), .A2(A[27]), .ZN(n119) );
  NAND2_X1 U176 ( .A1(n16), .A2(\B_not[27] ), .ZN(n120) );
  NAND2_X1 U177 ( .A1(A[27]), .A2(\B_not[27] ), .ZN(n121) );
  NAND3_X1 U178 ( .A1(n119), .A2(n120), .A3(n121), .ZN(\carry[28] ) );
  XOR2_X1 U179 ( .A(A[24]), .B(\B_not[24] ), .Z(n122) );
  XOR2_X1 U180 ( .A(n25), .B(n122), .Z(DIFF[24]) );
  XOR2_X1 U181 ( .A(A[25]), .B(\B_not[25] ), .Z(n126) );
  XOR2_X1 U182 ( .A(n126), .B(n90), .Z(DIFF[25]) );
  NAND2_X1 U183 ( .A1(A[25]), .A2(\B_not[25] ), .ZN(n127) );
  NAND2_X1 U184 ( .A1(\carry[25] ), .A2(A[25]), .ZN(n128) );
  NAND2_X1 U185 ( .A1(n3), .A2(\B_not[25] ), .ZN(n129) );
  NAND3_X1 U186 ( .A1(n128), .A2(n127), .A3(n129), .ZN(\carry[26] ) );
  XOR2_X1 U187 ( .A(n176), .B(A[2]), .Z(n130) );
  XOR2_X1 U188 ( .A(n85), .B(n130), .Z(DIFF[2]) );
  NAND2_X1 U189 ( .A1(\carry[2] ), .A2(n176), .ZN(n131) );
  NAND2_X1 U190 ( .A1(n27), .A2(A[2]), .ZN(n132) );
  NAND2_X1 U191 ( .A1(n176), .A2(A[2]), .ZN(n133) );
  XOR2_X1 U192 ( .A(A[30]), .B(\B_not[30] ), .Z(n134) );
  NAND2_X1 U193 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n135) );
  NAND2_X1 U194 ( .A1(\carry[30] ), .A2(\B_not[30] ), .ZN(n136) );
  NAND2_X1 U195 ( .A1(A[30]), .A2(\B_not[30] ), .ZN(n137) );
  NAND3_X1 U196 ( .A1(n135), .A2(n136), .A3(n137), .ZN(\carry[31] ) );
  XOR2_X1 U197 ( .A(\B_not[12] ), .B(A[12]), .Z(n138) );
  XOR2_X1 U198 ( .A(n13), .B(n138), .Z(DIFF[12]) );
  NAND2_X1 U199 ( .A1(\carry[12] ), .A2(A[12]), .ZN(n139) );
  XOR2_X1 U200 ( .A(\B_not[6] ), .B(A[6]), .Z(n141) );
  XOR2_X1 U201 ( .A(n51), .B(n141), .Z(DIFF[6]) );
  NAND2_X1 U202 ( .A1(\carry[6] ), .A2(\B_not[6] ), .ZN(n142) );
  NAND2_X1 U203 ( .A1(\carry[6] ), .A2(A[6]), .ZN(n143) );
  INV_X8 U204 ( .A(B[30]), .ZN(\B_not[30] ) );
  XOR2_X1 U205 ( .A(\B_not[13] ), .B(A[13]), .Z(n145) );
  XOR2_X1 U206 ( .A(n55), .B(n145), .Z(DIFF[13]) );
  XOR2_X1 U207 ( .A(A[29]), .B(\B_not[29] ), .Z(n149) );
  XOR2_X1 U208 ( .A(n61), .B(n149), .Z(DIFF[29]) );
  NAND2_X1 U209 ( .A1(\carry[29] ), .A2(A[29]), .ZN(n150) );
  NAND2_X1 U210 ( .A1(\carry[29] ), .A2(\B_not[29] ), .ZN(n151) );
  NAND2_X1 U211 ( .A1(A[29]), .A2(\B_not[29] ), .ZN(n152) );
  NAND3_X1 U212 ( .A1(n150), .A2(n151), .A3(n152), .ZN(\carry[30] ) );
  XOR2_X1 U213 ( .A(\B_not[14] ), .B(A[14]), .Z(n153) );
  XOR2_X1 U214 ( .A(n88), .B(n153), .Z(DIFF[14]) );
  NAND2_X1 U215 ( .A1(n14), .A2(\B_not[14] ), .ZN(n154) );
  NAND2_X1 U216 ( .A1(\carry[14] ), .A2(A[14]), .ZN(n155) );
  NAND3_X1 U217 ( .A1(n155), .A2(n156), .A3(n154), .ZN(\carry[15] ) );
  XOR2_X1 U218 ( .A(\B_not[8] ), .B(A[8]), .Z(n157) );
  XOR2_X1 U219 ( .A(n63), .B(n157), .Z(DIFF[8]) );
  NAND2_X1 U220 ( .A1(\carry[8] ), .A2(\B_not[8] ), .ZN(n158) );
  NAND2_X1 U221 ( .A1(\carry[8] ), .A2(A[8]), .ZN(n159) );
  XOR2_X1 U222 ( .A(\B_not[7] ), .B(A[7]), .Z(n161) );
  XOR2_X1 U223 ( .A(n89), .B(n161), .Z(DIFF[7]) );
  NAND2_X1 U224 ( .A1(n56), .A2(A[7]), .ZN(n163) );
  INV_X8 U225 ( .A(B[29]), .ZN(\B_not[29] ) );
  INV_X1 U226 ( .A(B[0]), .ZN(n165) );
  XOR2_X1 U227 ( .A(\B_not[23] ), .B(A[23]), .Z(n166) );
  XOR2_X1 U228 ( .A(n37), .B(n166), .Z(DIFF[23]) );
  NAND2_X1 U229 ( .A1(\carry[23] ), .A2(\B_not[23] ), .ZN(n167) );
  NAND2_X1 U230 ( .A1(\carry[23] ), .A2(A[23]), .ZN(n168) );
  NAND3_X1 U231 ( .A1(n168), .A2(n167), .A3(n169), .ZN(\carry[24] ) );
  XOR2_X1 U232 ( .A(\B_not[17] ), .B(A[17]), .Z(n170) );
  XOR2_X1 U233 ( .A(n54), .B(n170), .Z(DIFF[17]) );
  NAND2_X1 U234 ( .A1(\carry[17] ), .A2(\B_not[17] ), .ZN(n171) );
  NAND2_X1 U235 ( .A1(\carry[17] ), .A2(A[17]), .ZN(n172) );
  NAND3_X1 U236 ( .A1(n172), .A2(n171), .A3(n173), .ZN(\carry[18] ) );
  INV_X1 U237 ( .A(B[4]), .ZN(n174) );
  INV_X1 U238 ( .A(B[3]), .ZN(n175) );
  INV_X1 U239 ( .A(B[2]), .ZN(n176) );
  INV_X1 U240 ( .A(B[1]), .ZN(n177) );
  INV_X1 U241 ( .A(n6), .ZN(n178) );
  XNOR2_X1 U242 ( .A(A[0]), .B(n178), .ZN(DIFF[0]) );
  INV_X1 U243 ( .A(B[9]), .ZN(\B_not[9] ) );
  INV_X1 U244 ( .A(B[8]), .ZN(\B_not[8] ) );
  INV_X1 U245 ( .A(B[7]), .ZN(\B_not[7] ) );
  INV_X1 U246 ( .A(B[6]), .ZN(\B_not[6] ) );
  INV_X1 U247 ( .A(B[5]), .ZN(\B_not[5] ) );
  INV_X1 U248 ( .A(B[31]), .ZN(\B_not[31] ) );
  INV_X1 U249 ( .A(B[28]), .ZN(\B_not[28] ) );
  INV_X1 U250 ( .A(B[27]), .ZN(\B_not[27] ) );
  INV_X1 U251 ( .A(B[26]), .ZN(\B_not[26] ) );
  INV_X1 U252 ( .A(B[25]), .ZN(\B_not[25] ) );
  INV_X1 U253 ( .A(B[24]), .ZN(\B_not[24] ) );
  INV_X1 U254 ( .A(B[23]), .ZN(\B_not[23] ) );
  INV_X1 U255 ( .A(B[20]), .ZN(\B_not[20] ) );
  INV_X1 U256 ( .A(B[19]), .ZN(\B_not[19] ) );
  INV_X1 U257 ( .A(B[18]), .ZN(\B_not[18] ) );
  INV_X1 U258 ( .A(B[17]), .ZN(\B_not[17] ) );
  INV_X1 U259 ( .A(B[16]), .ZN(\B_not[16] ) );
  INV_X1 U260 ( .A(B[15]), .ZN(\B_not[15] ) );
  INV_X1 U261 ( .A(B[14]), .ZN(\B_not[14] ) );
  INV_X1 U262 ( .A(B[13]), .ZN(\B_not[13] ) );
  INV_X1 U263 ( .A(B[12]), .ZN(\B_not[12] ) );
  INV_X1 U264 ( .A(B[10]), .ZN(\B_not[10] ) );
endmodule


module up_island_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  AND4_X2 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(n6) );
  AND4_X1 U2 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(n1) );
  AND4_X1 U3 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n2) );
  AND4_X1 U4 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n3) );
  AND4_X1 U5 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n4) );
  INV_X1 U6 ( .A(NE), .ZN(EQ) );
  NAND2_X1 U7 ( .A1(n5), .A2(n6), .ZN(NE) );
  XNOR2_X1 U8 ( .A(B[11]), .B(A[11]), .ZN(n10) );
  XNOR2_X1 U9 ( .A(B[12]), .B(A[12]), .ZN(n9) );
  XNOR2_X1 U10 ( .A(B[13]), .B(A[13]), .ZN(n8) );
  XNOR2_X1 U11 ( .A(B[14]), .B(A[14]), .ZN(n7) );
  XNOR2_X1 U12 ( .A(B[7]), .B(A[7]), .ZN(n14) );
  XNOR2_X1 U13 ( .A(B[8]), .B(A[8]), .ZN(n13) );
  XNOR2_X1 U14 ( .A(B[9]), .B(A[9]), .ZN(n12) );
  XNOR2_X1 U15 ( .A(B[10]), .B(A[10]), .ZN(n11) );
  XNOR2_X1 U16 ( .A(B[3]), .B(A[3]), .ZN(n18) );
  XNOR2_X1 U17 ( .A(B[4]), .B(A[4]), .ZN(n17) );
  XNOR2_X1 U18 ( .A(B[5]), .B(A[5]), .ZN(n16) );
  XNOR2_X1 U19 ( .A(B[6]), .B(A[6]), .ZN(n15) );
  OAI22_X1 U20 ( .A1(n23), .A2(n24), .B1(B[1]), .B2(n23), .ZN(n22) );
  INV_X1 U21 ( .A(A[1]), .ZN(n24) );
  AND2_X1 U22 ( .A1(B[0]), .A2(n25), .ZN(n23) );
  OAI22_X1 U23 ( .A1(A[1]), .A2(n26), .B1(n26), .B2(n27), .ZN(n21) );
  INV_X1 U24 ( .A(B[1]), .ZN(n27) );
  NOR2_X1 U25 ( .A1(n25), .A2(B[0]), .ZN(n26) );
  INV_X1 U26 ( .A(A[0]), .ZN(n25) );
  XNOR2_X1 U27 ( .A(B[31]), .B(A[31]), .ZN(n20) );
  XNOR2_X1 U28 ( .A(B[2]), .B(A[2]), .ZN(n19) );
  NOR4_X1 U29 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n5) );
  NAND4_X1 U30 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XNOR2_X1 U31 ( .A(B[27]), .B(A[27]), .ZN(n35) );
  XNOR2_X1 U32 ( .A(B[28]), .B(A[28]), .ZN(n34) );
  XNOR2_X1 U33 ( .A(B[29]), .B(A[29]), .ZN(n33) );
  XNOR2_X1 U34 ( .A(B[30]), .B(A[30]), .ZN(n32) );
  NAND4_X1 U35 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XNOR2_X1 U36 ( .A(B[23]), .B(A[23]), .ZN(n39) );
  XNOR2_X1 U37 ( .A(B[24]), .B(A[24]), .ZN(n38) );
  XNOR2_X1 U38 ( .A(B[25]), .B(A[25]), .ZN(n37) );
  XNOR2_X1 U39 ( .A(B[26]), .B(A[26]), .ZN(n36) );
  NAND4_X1 U40 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XNOR2_X1 U41 ( .A(B[19]), .B(A[19]), .ZN(n43) );
  XNOR2_X1 U42 ( .A(B[20]), .B(A[20]), .ZN(n42) );
  XNOR2_X1 U43 ( .A(B[21]), .B(A[21]), .ZN(n41) );
  XNOR2_X1 U44 ( .A(B[22]), .B(A[22]), .ZN(n40) );
  NAND4_X1 U45 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XNOR2_X1 U46 ( .A(B[15]), .B(A[15]), .ZN(n47) );
  XNOR2_X1 U47 ( .A(B[16]), .B(A[16]), .ZN(n46) );
  XNOR2_X1 U48 ( .A(B[17]), .B(A[17]), .ZN(n45) );
  XNOR2_X1 U49 ( .A(B[18]), .B(A[18]), .ZN(n44) );
endmodule


module up_island_DW01_add_2 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] ;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X2 U1 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X2 U2 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X2 U3 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X2 U4 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X2 U5 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X2 U6 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U7 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  AND2_X1 U8 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U9 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U10 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U11 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U12 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  XOR2_X1 U13 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  AND2_X1 U14 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U15 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  XOR2_X1 U16 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  AND2_X1 U17 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U18 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  XOR2_X1 U19 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  AND2_X1 U20 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  XOR2_X1 U21 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  XOR2_X1 U23 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  AND2_X1 U24 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  XOR2_X1 U25 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  AND2_X1 U26 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  XOR2_X1 U27 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  AND2_X1 U28 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  XOR2_X1 U29 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  AND2_X1 U30 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  XOR2_X1 U31 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  AND2_X1 U32 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  XOR2_X1 U33 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  AND2_X1 U34 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  XOR2_X1 U35 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  AND2_X1 U36 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  XOR2_X1 U37 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  AND2_X1 U38 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  XOR2_X1 U39 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  AND2_X1 U40 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  XOR2_X1 U41 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  INV_X1 U42 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module up_island_DW01_add_1 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \carry[23] , \carry[22] , \carry[21] , \carry[20] , \carry[19] ,
         \carry[18] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[4] ,
         \carry[3] , \carry[2] , \carry[1] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40;

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .S(SUM[23]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  NAND3_X1 U1 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n2) );
  BUF_X1 U3 ( .A(B[0]), .Z(n3) );
  NAND3_X1 U4 ( .A1(n18), .A2(n19), .A3(n20), .ZN(\carry[10] ) );
  XOR2_X1 U5 ( .A(A[20]), .B(B[20]), .Z(n4) );
  XOR2_X1 U6 ( .A(n4), .B(\carry[20] ), .Z(SUM[20]) );
  NAND2_X2 U7 ( .A1(A[20]), .A2(B[20]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(A[20]), .A2(\carry[20] ), .ZN(n6) );
  NAND2_X1 U9 ( .A1(B[20]), .A2(\carry[20] ), .ZN(n7) );
  NAND3_X2 U10 ( .A1(n5), .A2(n6), .A3(n7), .ZN(\carry[21] ) );
  XOR2_X1 U11 ( .A(A[21]), .B(B[21]), .Z(n8) );
  XOR2_X1 U12 ( .A(n8), .B(\carry[21] ), .Z(SUM[21]) );
  NAND2_X1 U13 ( .A1(A[21]), .A2(B[21]), .ZN(n9) );
  NAND2_X1 U14 ( .A1(A[21]), .A2(\carry[21] ), .ZN(n10) );
  NAND2_X1 U15 ( .A1(B[21]), .A2(\carry[21] ), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n9), .A2(n10), .A3(n11), .ZN(\carry[22] ) );
  BUF_X1 U17 ( .A(n2), .Z(n12) );
  NAND3_X1 U18 ( .A1(n26), .A2(n27), .A3(n28), .ZN(\carry[15] ) );
  XOR2_X1 U19 ( .A(B[22]), .B(A[22]), .Z(n13) );
  XOR2_X1 U20 ( .A(\carry[22] ), .B(n13), .Z(SUM[22]) );
  NAND2_X1 U21 ( .A1(\carry[22] ), .A2(B[22]), .ZN(n14) );
  NAND2_X1 U22 ( .A1(\carry[22] ), .A2(A[22]), .ZN(n15) );
  NAND2_X1 U23 ( .A1(B[22]), .A2(A[22]), .ZN(n16) );
  NAND3_X1 U24 ( .A1(n14), .A2(n16), .A3(n15), .ZN(\carry[23] ) );
  XOR2_X1 U25 ( .A(A[9]), .B(B[9]), .Z(n17) );
  XOR2_X1 U26 ( .A(n17), .B(\carry[9] ), .Z(SUM[9]) );
  NAND2_X2 U27 ( .A1(A[9]), .A2(B[9]), .ZN(n18) );
  NAND2_X1 U28 ( .A1(A[9]), .A2(\carry[9] ), .ZN(n19) );
  NAND2_X1 U29 ( .A1(B[9]), .A2(\carry[9] ), .ZN(n20) );
  XOR2_X1 U30 ( .A(A[10]), .B(B[10]), .Z(n21) );
  XOR2_X1 U31 ( .A(n21), .B(n1), .Z(SUM[10]) );
  NAND2_X1 U32 ( .A1(A[10]), .A2(B[10]), .ZN(n22) );
  NAND2_X1 U33 ( .A1(A[10]), .A2(n1), .ZN(n23) );
  NAND2_X1 U34 ( .A1(B[10]), .A2(\carry[10] ), .ZN(n24) );
  NAND3_X1 U35 ( .A1(n22), .A2(n23), .A3(n24), .ZN(\carry[11] ) );
  AND2_X2 U36 ( .A1(B[0]), .A2(A[0]), .ZN(\carry[1] ) );
  XOR2_X1 U37 ( .A(A[14]), .B(B[14]), .Z(n25) );
  XOR2_X1 U38 ( .A(n25), .B(\carry[14] ), .Z(SUM[14]) );
  NAND2_X2 U39 ( .A1(A[14]), .A2(B[14]), .ZN(n26) );
  NAND2_X1 U40 ( .A1(A[14]), .A2(\carry[14] ), .ZN(n27) );
  NAND2_X1 U41 ( .A1(B[14]), .A2(\carry[14] ), .ZN(n28) );
  XOR2_X1 U42 ( .A(A[15]), .B(B[15]), .Z(n29) );
  XOR2_X1 U43 ( .A(n29), .B(n12), .Z(SUM[15]) );
  NAND2_X1 U44 ( .A1(A[15]), .A2(B[15]), .ZN(n30) );
  NAND2_X1 U45 ( .A1(A[15]), .A2(\carry[15] ), .ZN(n31) );
  NAND2_X1 U46 ( .A1(B[15]), .A2(n2), .ZN(n32) );
  NAND3_X1 U47 ( .A1(n32), .A2(n31), .A3(n30), .ZN(\carry[16] ) );
  XOR2_X1 U48 ( .A(A[1]), .B(B[1]), .Z(n33) );
  XOR2_X1 U49 ( .A(n33), .B(\carry[1] ), .Z(SUM[1]) );
  NAND2_X1 U50 ( .A1(A[1]), .A2(B[1]), .ZN(n34) );
  NAND2_X1 U51 ( .A1(A[1]), .A2(\carry[1] ), .ZN(n35) );
  NAND2_X1 U52 ( .A1(B[1]), .A2(\carry[1] ), .ZN(n36) );
  NAND3_X2 U53 ( .A1(n34), .A2(n35), .A3(n36), .ZN(\carry[2] ) );
  XOR2_X1 U54 ( .A(A[2]), .B(B[2]), .Z(n37) );
  XOR2_X1 U55 ( .A(n37), .B(\carry[2] ), .Z(SUM[2]) );
  NAND2_X1 U56 ( .A1(A[2]), .A2(B[2]), .ZN(n38) );
  NAND2_X1 U57 ( .A1(A[2]), .A2(\carry[2] ), .ZN(n39) );
  NAND2_X1 U58 ( .A1(B[2]), .A2(\carry[2] ), .ZN(n40) );
  NAND3_X1 U59 ( .A1(n38), .A2(n39), .A3(n40), .ZN(\carry[3] ) );
  XOR2_X1 U60 ( .A(n3), .B(A[0]), .Z(SUM[0]) );
endmodule


module up_island_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   \carry[60] , \carry[58] , \carry[57] , \carry[56] , \carry[48] ,
         \carry[47] , \carry[46] , \carry[45] , \carry[30] , \carry[29] ,
         \carry[20] , \carry[19] , \carry[15] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[1] , net55603, net55599, net55595, net55592,
         net55587, net55583, net55579, net55571, net55691, net55689, net55683,
         net55682, net55681, net55674, net55673, net55672, net55837, net55836,
         net55832, net55830, net55826, net55822, net55819, net55817, net55816,
         net55812, net55808, net55936, net55927, net55925, net55923, net55976,
         net55967, net55966, net55965, net55964, net55962, net56025, net56022,
         net56020, net56069, net56060, net56056, net56052, net56048, net56044,
         net56040, net56036, net56158, net56154, net56152, net56150, net56148,
         net56140, net56210, net56209, net56227, net56226, net56225, net56261,
         net56313, net56309, net56341, net56336, net56332, net56368, net56366,
         net56363, net56400, net56405, net56437, net56435, net56433, net56431,
         net56428, net56427, net56471, net56470, net56468, net56467, net56481,
         net56477, net56476, net56540, net56545, net56549, net56561, net56571,
         net56562, net56598, net56630, net56628, net56651, net56650, net56649,
         net56639, net56744, net56739, net56755, net56753, net56793, net56808,
         net56856, net56862, net56887, net56883, net56880, net56901, net56933,
         net56931, net57004, net57006, net57011, net57022, net57025, net57024,
         net57031, net57045, net57059, net57069, net57085, net57089, net57091,
         net57097, net57100, net58078, net58076, net58059, net58056, net58054,
         net58040, net58037, net58121, net58125, net58242, net58243, net58244,
         net58238, net58236, net58228, net58227, net58226, net58222, net58210,
         net58282, net58292, net58315, net58323, net58329, net58351, net58422,
         net58405, net58404, net58399, net58389, net58441, net58447, net59519,
         net59517, net60649, net60647, net60691, net60754, net60758, net60823,
         net60821, net60815, net60813, net60809, net60808, net60804, net60803,
         net60800, net60796, net60794, net60771, net60770, net60767, net60835,
         net60854, net60856, net60880, net60886, net62145, net62141, net62140,
         net62139, net62138, net62132, net62131, net62130, net62129, net62117,
         net62111, net62110, net62177, net62194, net62200, net62205, net62212,
         net62218, net62273, net62290, net62338, net62309, net59538, net59537,
         net56047, net56045, net64022, net64020, net64053, net64059, net65124,
         net65126, net65225, net65221, net65219, net65201, net65199, net65196,
         net65192, net65188, net65160, net65159, net65153, net65144, net65234,
         net65272, net65290, net65299, net65309, net65321, net65637, net65638,
         net65704, net65702, net65688, net65684, net65683, net67391, net67389,
         net67385, net67373, net67370, net67368, net67360, net67359, net67357,
         net67355, net67423, net67429, net67433, net67457, net67466, net60799,
         net69139, net69132, net69126, net69124, net69119, net69117, net69094,
         net69089, net69168, net69188, net69202, net69203, net70500, net70495,
         net70488, net70487, net70483, net70482, net70480, net70474, net70465,
         net70464, net70460, net70456, net70443, net70524, net70527, net72097,
         net72087, net72085, net65288, net65181, net65179, net73498, net73494,
         net73492, net73491, net73490, net73489, net73488, net73487, net73473,
         net73472, net73468, net73519, net73518, net73528, net73527, net73526,
         net73525, net73524, net73562, net73570, net73589, net73634, net73656,
         net73660, net73669, net73675, net65183, net65687, net65686, net65680,
         net65675, net57080, net56371, net56370, net75678, net75759, net75757,
         net75743, net75734, net75725, net75723, net75720, net75718, net75699,
         net75831, net75842, net75844, net56859, net77806, net77785, net77776,
         net77768, net77766, net77765, net77748, net77818, net77817, net77826,
         net77831, net56041, net58038, net56817, net56144, net79856, net79855,
         net79851, net79849, net79844, net79836, net79832, net79866, net79893,
         net79896, net79904, net79930, net79929, net79928, net79933, net73596,
         net62137, net62289, net57103, net57061, net56791, net56335, net56334,
         net56333, net73577, net73566, net73564, net65215, net64058,
         \carry[39] , net67379, \carry[17] , \carry[28] , \carry[27] ,
         net82439, net82430, net82429, net82427, net82423, net82419, net82413,
         net82412, net82405, net82402, net82394, net82391, net82387, net82385,
         net82384, net82383, net82381, net82377, net82373, net82369, net82367,
         net82365, net82363, net82355, net82338, net82333, net82494, net82504,
         net82508, net82510, net82512, net82511, net82516, net82522, net82542,
         net82565, net84135, net84131, net84129, net84122, net84109, net84105,
         net84099, net73663, net73561, net73557, net73554, net65191, net64019,
         net64012, net64010, net57019, net62344, net62332, net62326, net62307,
         net56569, net56054, net69164, net65709, net65697, net65693, net65691,
         net65685, net65679, net65678, net65677, net65673, net65671, net65659,
         net65658, \carry[32] , net58409, net58206, net58069, net58061,
         net58055, net84167, net84166, net75846, net82410, net82409, net82378,
         net73517, net58450, net58449, net58424, net58326, net58321, net58320,
         net58289, net58066, net58064, net58063, net58060, net58057, net56855,
         net56147, net56142, \carry[53] , net70458, net69072, net67456,
         net67421, net55937, net67465, net67462, net57116, net56888,
         \carry[18] , net82548, net82523, net82375, net70489, net69130,
         net69110, net84123, net84111, net75750, net75745, net75736, net75726,
         net75707, net75705, net55680, net58440, net58419, net58417, net58394,
         net58393, net58385, net58384, net58327, net65682, net59514,
         \carry[3] , net79932, net79914, net73580, net79908, net75853,
         net60817, net60810, net60805, net60798, net60797, net60779, net60768,
         net57039, net55833, net87602, net87601, net87597, net87594, net87578,
         net87623, net73567, net73556, net65251, net65202, net65200, net65197,
         net65184, net75735, net75731, net62181, \carry[43] , n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395;

  NOR2_X2 net58124 ( .A1(net58404), .A2(net58405), .ZN(net58315) );
  NAND3_X1 net57010 ( .A1(net62110), .A2(net62111), .A3(n297), .ZN(net56158)
         );
  NAND2_X2 net62274 ( .A1(net62309), .A2(net60815), .ZN(net60808) );
  NAND2_X2 net62276 ( .A1(B[24]), .A2(net60813), .ZN(net60809) );
  NAND2_X2 net65122 ( .A1(net65144), .A2(n288), .ZN(net55817) );
  NAND2_X2 syn338 ( .A1(net56481), .A2(B[12]), .ZN(net69094) );
  NAND3_X1 net56885 ( .A1(net69089), .A2(net55925), .A3(n279), .ZN(net56020)
         );
  NAND2_X2 net70438 ( .A1(n270), .A2(net70443), .ZN(net69132) );
  INV_X2 syn301 ( .A(n265), .ZN(net56753) );
  INV_X2 syn271 ( .A(net73468), .ZN(net73490) );
  INV_X2 syn44 ( .A(B[8]), .ZN(n262) );
  INV_X2 syn371 ( .A(net75757), .ZN(net56336) );
  NAND2_X2 net58346 ( .A1(B[50]), .A2(A[50]), .ZN(net56041) );
  NAND2_X2 syn194 ( .A1(A[39]), .A2(B[39]), .ZN(net79844) );
  INV_X2 syn454 ( .A(n223), .ZN(n222) );
  NAND3_X1 net56021 ( .A1(net67355), .A2(net67391), .A3(net67357), .ZN(
        net55976) );
  MUX2_X1 syn755 ( .A(net82338), .B(n203), .S(n200), .Z(n181) );
  NAND2_X2 syn753 ( .A1(A[11]), .A2(net82367), .ZN(n203) );
  XNOR2_X2 syn751 ( .A(n199), .B(net82367), .ZN(n201) );
  INV_X2 syn750 ( .A(n202), .ZN(net55967) );
  XNOR2_X2 syn749 ( .A(B[10]), .B(A[10]), .ZN(n202) );
  NAND2_X2 syn747 ( .A1(n201), .A2(net82365), .ZN(n182) );
  INV_X2 syn721 ( .A(net82383), .ZN(net82427) );
  NAND2_X2 syn717 ( .A1(net82381), .A2(net82384), .ZN(n192) );
  INV_X2 syn704 ( .A(net82381), .ZN(net82387) );
  NAND2_X2 syn687 ( .A1(net82419), .A2(net70500), .ZN(n195) );
  NAND2_X2 syn649 ( .A1(net82367), .A2(net82365), .ZN(net82377) );
  INV_X2 syn643 ( .A(net82338), .ZN(net82419) );
  INV_X2 syn640 ( .A(n199), .ZN(n200) );
  OAI21_X2 syn638 ( .B1(net82413), .B2(net82363), .A(n198), .ZN(n199) );
  NAND2_X2 syn636 ( .A1(A[10]), .A2(net77826), .ZN(n198) );
  INV_X2 syn633 ( .A(net82412), .ZN(net82413) );
  AND3_X2 syn502 ( .A1(n196), .A2(n195), .A3(n194), .ZN(n185) );
  NAND2_X2 syn245 ( .A1(net82384), .A2(net70500), .ZN(net82383) );
  INV_X2 syn25 ( .A(net56025), .ZN(net82355) );
  NAND2_X2 net82294 ( .A1(n181), .A2(n182), .ZN(SUM[11]) );
  NAND3_X1 net75835 ( .A1(net56333), .A2(n62), .A3(n166), .ZN(net75831) );
  NAND2_X2 net84066 ( .A1(n162), .A2(net84105), .ZN(net75743) );
  NAND2_X2 net84042 ( .A1(net57045), .A2(n161), .ZN(net56476) );
  NAND2_X2 net84068 ( .A1(net75725), .A2(n160), .ZN(net75757) );
  AOI21_X2 net65125 ( .B1(net65159), .B2(net65160), .A(n153), .ZN(net65126) );
  NAND2_X2 net62260 ( .A1(net60770), .A2(net60771), .ZN(net60647) );
  INV_X2 syn19 ( .A(B[31]), .ZN(net65673) );
  NAND2_X2 syn40 ( .A1(net65673), .A2(net65671), .ZN(net65679) );
  NAND2_X2 net58373 ( .A1(net56041), .A2(net58399), .ZN(net58236) );
  NAND3_X1 net56627 ( .A1(net58076), .A2(net56041), .A3(net58078), .ZN(
        net57006) );
  OAI21_X2 net73459 ( .B1(A[7]), .B2(B[7]), .A(net73468), .ZN(net72087) );
  AOI21_X2 net70423 ( .B1(net70456), .B2(net69094), .A(net70458), .ZN(net56808) );
  NAND2_X2 syn745 ( .A1(net82375), .A2(net82423), .ZN(net82391) );
  NOR2_X2 syn498 ( .A1(n105), .A2(net82369), .ZN(net82394) );
  NOR2_X2 syn520 ( .A1(net82373), .A2(n105), .ZN(net82402) );
  NAND2_X2 net70430 ( .A1(B[14]), .A2(net70443), .ZN(net69110) );
  NAND2_X2 syn515 ( .A1(net82384), .A2(net70489), .ZN(n108) );
  NAND2_X2 net55972 ( .A1(B[11]), .A2(A[11]), .ZN(net82338) );
  NAND3_X1 syn632 ( .A1(n49), .A2(net82387), .A3(net82510), .ZN(net82412) );
  NAND3_X1 syn737 ( .A1(net82548), .A2(net82510), .A3(net82387), .ZN(net82430)
         );
  NAND3_X1 syn739 ( .A1(net82523), .A2(n3), .A3(n111), .ZN(net82405) );
  INV_X2 syn653 ( .A(net82375), .ZN(n111) );
  NAND3_X1 syn689 ( .A1(net82523), .A2(net82439), .A3(n111), .ZN(n110) );
  NOR2_X2 syn510 ( .A1(n104), .A2(n105), .ZN(n107) );
  NAND2_X2 net84036 ( .A1(net75726), .A2(net84111), .ZN(\carry[45] ) );
  NAND2_X2 net84060 ( .A1(n103), .A2(net84109), .ZN(net75725) );
  NOR2_X2 syn164 ( .A1(A[43]), .A2(net75745), .ZN(net84123) );
  INV_X2 net84067 ( .A(net75726), .ZN(net75745) );
  NAND3_X1 net58376 ( .A1(B[49]), .A2(A[49]), .A3(net58389), .ZN(net58242) );
  NAND2_X2 net58374 ( .A1(net58384), .A2(net58385), .ZN(net58238) );
  NAND3_X1 net65644 ( .A1(net59514), .A2(net65704), .A3(net69164), .ZN(
        net56628) );
  OAI21_X2 net60751 ( .B1(net60823), .B2(net60767), .A(net60768), .ZN(net56471) );
  INV_X2 net62278 ( .A(net60770), .ZN(net60810) );
  AND2_X2 net60757 ( .A1(n72), .A2(n73), .ZN(net60758) );
  NAND2_X2 net62247 ( .A1(B[24]), .A2(A[24]), .ZN(net55833) );
  NOR2_X2 net62259 ( .A1(n75), .A2(net60779), .ZN(net57039) );
  NAND2_X2 syn223 ( .A1(net87602), .A2(net87601), .ZN(net87578) );
  INV_X2 syn28 ( .A(net56540), .ZN(net87594) );
  INV_X2 net65132 ( .A(A[37]), .ZN(net64012) );
  INV_X2 net65131 ( .A(B[37]), .ZN(net64010) );
  OAI21_X2 net65134 ( .B1(A[37]), .B2(B[37]), .A(net65153), .ZN(net64020) );
  NAND3_X1 net84034 ( .A1(net62181), .A2(net84167), .A3(net56333), .ZN(
        \carry[43] ) );
  INV_X2 net84062 ( .A(net75723), .ZN(net75731) );
  INV_X2 syn283 ( .A(n35), .ZN(n22) );
  NAND2_X2 syn282 ( .A1(n34), .A2(n33), .ZN(n35) );
  NAND2_X2 syn274 ( .A1(net87578), .A2(A[61]), .ZN(n34) );
  NAND2_X2 syn272 ( .A1(net87578), .A2(B[61]), .ZN(n33) );
  NAND2_X2 syn263 ( .A1(A[62]), .A2(B[62]), .ZN(n26) );
  NAND3_X1 syn261 ( .A1(n27), .A2(n26), .A3(net56649), .ZN(n31) );
  INV_X2 syn236 ( .A(net87594), .ZN(n29) );
  NAND3_X1 syn234 ( .A1(B[62]), .A2(A[62]), .A3(n29), .ZN(n28) );
  OAI21_X2 syn197 ( .B1(n19), .B2(n20), .A(n28), .ZN(n17) );
  NOR2_X2 syn190 ( .A1(A[62]), .A2(B[62]), .ZN(n27) );
  NAND3_X1 syn189 ( .A1(n20), .A2(n26), .A3(net56649), .ZN(n25) );
  XNOR2_X2 syn182 ( .A(A[62]), .B(n18), .ZN(net56477) );
  XNOR2_X2 syn172 ( .A(B[61]), .B(A[61]), .ZN(net87597) );
  NOR2_X2 syn146 ( .A1(B[61]), .A2(A[61]), .ZN(n23) );
  NOR2_X2 syn142 ( .A1(B[61]), .A2(A[61]), .ZN(n21) );
  NAND3_X1 syn141 ( .A1(net56226), .A2(net56225), .A3(net56227), .ZN(net87623)
         );
  NAND2_X2 syn69 ( .A1(B[61]), .A2(A[61]), .ZN(n20) );
  INV_X2 syn46 ( .A(net87578), .ZN(n19) );
  INV_X2 syn22 ( .A(B[62]), .ZN(n18) );
  NOR2_X2 net88854 ( .A1(n16), .A2(n17), .ZN(net56650) );
  NAND2_X2 net88860 ( .A1(net56540), .A2(B[62]), .ZN(net87602) );
  NAND2_X2 net88859 ( .A1(net56540), .A2(A[62]), .ZN(net87601) );
  INV_X1 U1 ( .A(net62131), .ZN(net73561) );
  INV_X1 U2 ( .A(net62131), .ZN(net62137) );
  INV_X1 U3 ( .A(n359), .ZN(n58) );
  BUF_X1 U4 ( .A(n176), .Z(n1) );
  NAND2_X1 U5 ( .A1(net82430), .A2(n2), .ZN(n180) );
  AND2_X1 U6 ( .A1(net82384), .A2(net70488), .ZN(n2) );
  BUF_X1 U7 ( .A(net73517), .Z(n3) );
  NAND2_X1 U8 ( .A1(n118), .A2(B[17]), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n118), .A2(B[17]), .ZN(net57116) );
  AND3_X2 U10 ( .A1(net62138), .A2(net62139), .A3(net62137), .ZN(n5) );
  NAND3_X1 U11 ( .A1(n247), .A2(n246), .A3(n245), .ZN(n6) );
  NAND3_X1 U12 ( .A1(net56888), .A2(n114), .A3(n115), .ZN(n116) );
  NAND3_X1 U13 ( .A1(net55680), .A2(net55681), .A3(net55682), .ZN(\carry[46] )
         );
  NOR2_X1 U14 ( .A1(net65680), .A2(net56435), .ZN(n7) );
  NAND2_X1 U15 ( .A1(n61), .A2(B[47]), .ZN(n8) );
  NAND3_X1 U16 ( .A1(n390), .A2(n389), .A3(n388), .ZN(n9) );
  NAND2_X2 U17 ( .A1(n321), .A2(A[56]), .ZN(n389) );
  NAND3_X1 U18 ( .A1(net55962), .A2(n369), .A3(n368), .ZN(n337) );
  NOR2_X1 U19 ( .A1(net65680), .A2(net56435), .ZN(net65684) );
  NAND3_X1 U20 ( .A1(n113), .A2(net57116), .A3(n112), .ZN(n10) );
  NOR2_X2 U21 ( .A1(n41), .A2(net65309), .ZN(net65290) );
  BUF_X2 U22 ( .A(net73517), .Z(net82439) );
  BUF_X1 U23 ( .A(net73517), .Z(net82548) );
  AND3_X2 U24 ( .A1(net62138), .A2(net62139), .A3(net62137), .ZN(net73596) );
  NOR2_X1 U25 ( .A1(n36), .A2(n23), .ZN(n24) );
  NAND2_X1 U26 ( .A1(\carry[1] ), .A2(n81), .ZN(n11) );
  NAND2_X1 U27 ( .A1(\carry[1] ), .A2(n81), .ZN(n89) );
  NAND3_X1 U28 ( .A1(n86), .A2(n95), .A3(n88), .ZN(n12) );
  NAND2_X2 U29 ( .A1(n94), .A2(n93), .ZN(n88) );
  NAND2_X2 U30 ( .A1(n146), .A2(n145), .ZN(net73517) );
  NOR2_X1 U31 ( .A1(n37), .A2(n22), .ZN(n16) );
  BUF_X1 U32 ( .A(n357), .Z(n13) );
  NAND2_X1 U33 ( .A1(\carry[46] ), .A2(B[46]), .ZN(n14) );
  NAND3_X1 U34 ( .A1(net56261), .A2(n353), .A3(n354), .ZN(n15) );
  AND3_X2 U35 ( .A1(net56226), .A2(net56227), .A3(net56225), .ZN(n36) );
  OAI21_X1 U36 ( .B1(n21), .B2(n36), .A(n20), .ZN(n32) );
  XNOR2_X1 U37 ( .A(n32), .B(net56598), .ZN(SUM[62]) );
  OAI21_X1 U38 ( .B1(n24), .B2(n25), .A(n31), .ZN(n30) );
  INV_X1 U39 ( .A(n30), .ZN(net56651) );
  INV_X1 U40 ( .A(net87623), .ZN(n37) );
  NOR2_X1 U41 ( .A1(n40), .A2(n39), .ZN(net75735) );
  AOI21_X2 U42 ( .B1(net75735), .B2(net75736), .A(net75707), .ZN(net55680) );
  NOR2_X1 U43 ( .A1(\carry[43] ), .A2(B[43]), .ZN(n40) );
  NAND2_X2 U44 ( .A1(net75731), .A2(B[45]), .ZN(n39) );
  NOR2_X1 U45 ( .A1(n38), .A2(n39), .ZN(net75705) );
  NAND2_X1 U46 ( .A1(net84135), .A2(net75731), .ZN(net84111) );
  NOR2_X1 U47 ( .A1(\carry[43] ), .A2(B[43]), .ZN(n38) );
  NAND2_X1 U48 ( .A1(net79932), .A2(B[42]), .ZN(net62181) );
  NAND2_X2 U49 ( .A1(net75723), .A2(net75726), .ZN(net84122) );
  NAND2_X1 U50 ( .A1(net82512), .A2(A[42]), .ZN(net84167) );
  NAND2_X1 U51 ( .A1(net79932), .A2(B[42]), .ZN(net84166) );
  OAI21_X1 U52 ( .B1(n46), .B2(n43), .A(n44), .ZN(n41) );
  NAND2_X2 U53 ( .A1(net65202), .A2(B[38]), .ZN(n44) );
  INV_X1 U54 ( .A(net65153), .ZN(net65202) );
  NAND2_X1 U55 ( .A1(net65197), .A2(net65196), .ZN(n46) );
  NAND2_X2 U56 ( .A1(B[38]), .A2(net65192), .ZN(n43) );
  INV_X2 U57 ( .A(n43), .ZN(net65225) );
  NAND2_X2 U58 ( .A1(B[37]), .A2(A[37]), .ZN(net65153) );
  NAND2_X1 U59 ( .A1(net73596), .A2(n45), .ZN(net65197) );
  BUF_X1 U60 ( .A(net65197), .Z(net73669) );
  INV_X1 U61 ( .A(net65251), .ZN(n45) );
  AND2_X1 U62 ( .A1(n45), .A2(net65153), .ZN(net73567) );
  AND2_X1 U63 ( .A1(n45), .A2(net73557), .ZN(net73556) );
  NAND2_X1 U64 ( .A1(net65201), .A2(net65184), .ZN(net65251) );
  INV_X1 U65 ( .A(A[36]), .ZN(net65184) );
  AOI21_X2 U66 ( .B1(net65200), .B2(net65201), .A(n42), .ZN(net65196) );
  INV_X2 U67 ( .A(B[36]), .ZN(n42) );
  NOR2_X2 U68 ( .A1(A[36]), .A2(net65183), .ZN(net65200) );
  INV_X2 U69 ( .A(net65192), .ZN(net65215) );
  NAND2_X1 U70 ( .A1(n5), .A2(net73556), .ZN(net73554) );
  NAND2_X1 U71 ( .A1(n5), .A2(net73567), .ZN(net73564) );
  XNOR2_X2 U72 ( .A(B[36]), .B(A[36]), .ZN(net64022) );
  NAND2_X2 U73 ( .A1(net65183), .A2(net65124), .ZN(net65144) );
  NAND2_X2 U74 ( .A1(A[36]), .A2(net65183), .ZN(net65191) );
  NAND2_X1 U75 ( .A1(n165), .A2(net84099), .ZN(n47) );
  NOR2_X1 U76 ( .A1(net75745), .A2(B[43]), .ZN(net84099) );
  OAI21_X1 U77 ( .B1(net79908), .B2(net60805), .A(net60817), .ZN(net60797) );
  NAND3_X1 U78 ( .A1(n228), .A2(n177), .A3(net79844), .ZN(n48) );
  NAND3_X1 U79 ( .A1(n228), .A2(n177), .A3(net79844), .ZN(net73577) );
  AND3_X2 U80 ( .A1(n185), .A2(n184), .A3(n183), .ZN(net70460) );
  INV_X1 U81 ( .A(net82542), .ZN(n49) );
  NAND2_X1 U82 ( .A1(\carry[48] ), .A2(A[48]), .ZN(n50) );
  NAND2_X1 U83 ( .A1(n48), .A2(net79856), .ZN(n51) );
  OAI21_X1 U84 ( .B1(net73494), .B2(net73489), .A(net73468), .ZN(n264) );
  AND2_X2 U85 ( .A1(n51), .A2(net79849), .ZN(net79904) );
  AND2_X1 U86 ( .A1(n77), .A2(n78), .ZN(n52) );
  AND2_X1 U87 ( .A1(n77), .A2(n78), .ZN(net73580) );
  NAND2_X1 U88 ( .A1(\carry[53] ), .A2(B[53]), .ZN(n53) );
  NAND2_X1 U89 ( .A1(\carry[47] ), .A2(A[47]), .ZN(n54) );
  NAND2_X1 U90 ( .A1(net57103), .A2(B[42]), .ZN(n55) );
  NAND2_X1 U91 ( .A1(n333), .A2(A[46]), .ZN(n56) );
  NAND2_X1 U92 ( .A1(n333), .A2(A[46]), .ZN(n393) );
  NAND2_X1 U93 ( .A1(n373), .A2(B[55]), .ZN(n57) );
  XNOR2_X1 U94 ( .A(n58), .B(n350), .ZN(SUM[60]) );
  NAND2_X1 U95 ( .A1(n229), .A2(A[42]), .ZN(n59) );
  AND2_X2 U96 ( .A1(net79933), .A2(net79849), .ZN(net79914) );
  NAND2_X1 U97 ( .A1(net67359), .A2(net67360), .ZN(n60) );
  NAND3_X1 U98 ( .A1(n56), .A2(n14), .A3(n392), .ZN(n61) );
  BUF_X1 U99 ( .A(n59), .Z(n62) );
  NOR2_X1 U100 ( .A1(net82385), .A2(n188), .ZN(n183) );
  BUF_X1 U101 ( .A(net79836), .Z(n63) );
  INV_X1 U102 ( .A(n1), .ZN(n64) );
  NAND2_X1 U103 ( .A1(net82423), .A2(net70500), .ZN(n65) );
  NAND2_X1 U104 ( .A1(net82429), .A2(n66), .ZN(n196) );
  INV_X1 U105 ( .A(n65), .ZN(n66) );
  NAND2_X1 U106 ( .A1(net70480), .A2(net70474), .ZN(net70500) );
  INV_X1 U107 ( .A(n105), .ZN(net82423) );
  AOI21_X1 U108 ( .B1(net75705), .B2(net75736), .A(net75707), .ZN(net56880) );
  NAND2_X1 U109 ( .A1(n6), .A2(B[48]), .ZN(n67) );
  NAND2_X1 U110 ( .A1(n317), .A2(B[26]), .ZN(n68) );
  AOI21_X2 U111 ( .B1(n110), .B2(n107), .A(n106), .ZN(n109) );
  XNOR2_X1 U112 ( .A(net87623), .B(net87597), .ZN(SUM[61]) );
  AND2_X1 U113 ( .A1(n197), .A2(n180), .ZN(n69) );
  NAND3_X1 U114 ( .A1(net57039), .A2(n71), .A3(net55833), .ZN(n70) );
  NAND2_X1 U115 ( .A1(n70), .A2(A[25]), .ZN(net60691) );
  NAND2_X1 U116 ( .A1(n70), .A2(A[25]), .ZN(net55689) );
  NAND2_X1 U117 ( .A1(net60797), .A2(n74), .ZN(n71) );
  AND2_X1 U118 ( .A1(n73), .A2(A[24]), .ZN(n74) );
  INV_X2 U119 ( .A(net60798), .ZN(net60817) );
  OAI21_X1 U120 ( .B1(net69202), .B2(net60804), .A(net60817), .ZN(net69203) );
  OAI21_X1 U121 ( .B1(net62289), .B2(net60804), .A(net60817), .ZN(net60796) );
  OAI21_X2 U122 ( .B1(net60823), .B2(net60803), .A(net60817), .ZN(n72) );
  NAND2_X2 U123 ( .A1(net60768), .A2(net60794), .ZN(net60798) );
  NOR2_X2 U124 ( .A1(A[22]), .A2(B[22]), .ZN(net60805) );
  NAND2_X2 U125 ( .A1(net60808), .A2(net60809), .ZN(net60779) );
  NOR2_X1 U126 ( .A1(net75853), .A2(net62307), .ZN(n75) );
  AND3_X1 U127 ( .A1(net62344), .A2(n151), .A3(net62332), .ZN(net75853) );
  NAND3_X1 U128 ( .A1(net82516), .A2(net55832), .A3(net55833), .ZN(net82511)
         );
  NAND3_X1 U129 ( .A1(net60754), .A2(net65321), .A3(net55833), .ZN(net60880)
         );
  NAND3_X1 U130 ( .A1(net60886), .A2(net55832), .A3(net55833), .ZN(net56862)
         );
  NAND2_X2 U131 ( .A1(net60810), .A2(net60794), .ZN(n73) );
  AND2_X1 U132 ( .A1(n73), .A2(A[24]), .ZN(net60854) );
  XNOR2_X2 U133 ( .A(B[24]), .B(A[24]), .ZN(net62338) );
  AND3_X2 U134 ( .A1(net56054), .A2(net62344), .A3(net62332), .ZN(net79908) );
  NOR2_X1 U135 ( .A1(net79908), .A2(net62307), .ZN(net60799) );
  NAND2_X2 U136 ( .A1(A[22]), .A2(B[22]), .ZN(net60768) );
  INV_X2 U137 ( .A(net60768), .ZN(net60815) );
  NAND3_X1 U138 ( .A1(net73580), .A2(net79914), .A3(net56371), .ZN(net79932)
         );
  BUF_X1 U139 ( .A(n52), .Z(net56791) );
  NAND3_X1 U140 ( .A1(n52), .A2(net79904), .A3(net56371), .ZN(net57103) );
  OR2_X1 U141 ( .A1(n79), .A2(net79832), .ZN(n78) );
  INV_X1 U142 ( .A(A[41]), .ZN(n79) );
  NAND2_X1 U143 ( .A1(net79836), .A2(n80), .ZN(n77) );
  AND2_X1 U144 ( .A1(net79855), .A2(A[41]), .ZN(n80) );
  BUF_X1 U145 ( .A(net79904), .Z(net57061) );
  NAND2_X1 U146 ( .A1(B[41]), .A2(A[41]), .ZN(net56371) );
  OR2_X1 U147 ( .A1(net79929), .A2(net79832), .ZN(net79928) );
  NAND2_X1 U148 ( .A1(n76), .A2(net79832), .ZN(net56630) );
  INV_X2 U149 ( .A(net79832), .ZN(net79851) );
  NAND2_X1 U150 ( .A1(n63), .A2(net79855), .ZN(n76) );
  AND2_X1 U151 ( .A1(net79855), .A2(A[41]), .ZN(net79930) );
  NAND2_X1 U152 ( .A1(n82), .A2(n83), .ZN(\carry[3] ) );
  NAND2_X1 U153 ( .A1(\carry[3] ), .A2(B[3]), .ZN(net62205) );
  BUF_X1 U154 ( .A(\carry[3] ), .Z(net56405) );
  NAND2_X1 U155 ( .A1(\carry[3] ), .A2(B[3]), .ZN(net69168) );
  NAND2_X1 U156 ( .A1(n92), .A2(n96), .ZN(n83) );
  INV_X1 U157 ( .A(n99), .ZN(n96) );
  AND2_X1 U158 ( .A1(A[3]), .A2(n96), .ZN(net77765) );
  XNOR2_X1 U159 ( .A(n96), .B(A[2]), .ZN(net77785) );
  INV_X1 U160 ( .A(B[2]), .ZN(n99) );
  NAND3_X1 U161 ( .A1(n90), .A2(n89), .A3(n91), .ZN(n92) );
  NAND2_X1 U162 ( .A1(n87), .A2(A[2]), .ZN(n82) );
  INV_X1 U163 ( .A(B[2]), .ZN(n98) );
  INV_X1 U164 ( .A(B[2]), .ZN(n85) );
  NAND2_X1 U165 ( .A1(net57022), .A2(n97), .ZN(n90) );
  NAND3_X1 U166 ( .A1(n90), .A2(n11), .A3(n91), .ZN(net77776) );
  BUF_X2 U167 ( .A(B[1]), .Z(n97) );
  NAND2_X1 U168 ( .A1(n97), .A2(n81), .ZN(n91) );
  BUF_X1 U169 ( .A(n97), .Z(net77831) );
  NAND2_X1 U170 ( .A1(net57022), .A2(n97), .ZN(n95) );
  BUF_X2 U171 ( .A(A[1]), .Z(n81) );
  BUF_X1 U172 ( .A(n81), .Z(net77806) );
  NAND2_X1 U173 ( .A1(net57022), .A2(n81), .ZN(n86) );
  NAND3_X1 U174 ( .A1(n88), .A2(n95), .A3(n86), .ZN(n87) );
  NAND2_X1 U175 ( .A1(n12), .A2(net77766), .ZN(net77768) );
  NAND2_X1 U176 ( .A1(n85), .A2(n84), .ZN(n93) );
  INV_X1 U177 ( .A(A[1]), .ZN(n84) );
  NAND2_X1 U178 ( .A1(n98), .A2(net77748), .ZN(n94) );
  INV_X1 U179 ( .A(B[1]), .ZN(net77748) );
  NOR2_X1 U180 ( .A1(n101), .A2(net65682), .ZN(n100) );
  AOI21_X1 U181 ( .B1(n100), .B2(net65697), .A(net65659), .ZN(\carry[32] ) );
  AND2_X2 U182 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n101) );
  NOR2_X1 U183 ( .A1(n101), .A2(net65682), .ZN(net65685) );
  BUF_X1 U184 ( .A(n101), .Z(net65702) );
  NAND2_X2 U185 ( .A1(net65677), .A2(net59514), .ZN(net65682) );
  NOR2_X1 U186 ( .A1(net65682), .A2(net65702), .ZN(net65658) );
  NAND2_X1 U187 ( .A1(\carry[30] ), .A2(A[30]), .ZN(net56435) );
  XNOR2_X2 U188 ( .A(A[30]), .B(B[30]), .ZN(net59517) );
  NAND2_X1 U189 ( .A1(A[30]), .A2(B[30]), .ZN(net59514) );
  NAND2_X2 U190 ( .A1(net65691), .A2(net65677), .ZN(net65693) );
  NOR2_X2 U191 ( .A1(net65675), .A2(net65677), .ZN(net65678) );
  NOR2_X2 U192 ( .A1(net65680), .A2(net59514), .ZN(net65683) );
  NAND2_X1 U193 ( .A1(n102), .A2(net58393), .ZN(net58327) );
  NAND2_X1 U194 ( .A1(net58327), .A2(net58326), .ZN(net58057) );
  NAND2_X1 U195 ( .A1(net58327), .A2(net58409), .ZN(net58449) );
  NAND2_X1 U196 ( .A1(net58327), .A2(net58409), .ZN(net58321) );
  NAND2_X1 U197 ( .A1(net58440), .A2(net58384), .ZN(n102) );
  NAND2_X2 U198 ( .A1(A[49]), .A2(B[49]), .ZN(net58393) );
  NAND2_X1 U199 ( .A1(net58394), .A2(net58393), .ZN(net79896) );
  NAND2_X1 U200 ( .A1(net58394), .A2(net58393), .ZN(net56147) );
  NAND3_X1 U201 ( .A1(net58227), .A2(net56152), .A3(net58226), .ZN(net58440)
         );
  NAND2_X1 U202 ( .A1(net58440), .A2(net58384), .ZN(net58394) );
  NAND2_X1 U203 ( .A1(net58417), .A2(net58419), .ZN(net58384) );
  INV_X1 U204 ( .A(net58384), .ZN(net58222) );
  INV_X2 U205 ( .A(A[49]), .ZN(net58419) );
  INV_X2 U206 ( .A(B[49]), .ZN(net58417) );
  NAND2_X2 U207 ( .A1(A[49]), .A2(B[49]), .ZN(net58385) );
  AND3_X2 U208 ( .A1(n67), .A2(n50), .A3(net58226), .ZN(net58329) );
  INV_X2 U209 ( .A(net75750), .ZN(net75707) );
  NAND2_X2 U210 ( .A1(net75745), .A2(B[45]), .ZN(net75750) );
  NAND2_X1 U211 ( .A1(net75846), .A2(n103), .ZN(net75736) );
  INV_X2 U212 ( .A(A[43]), .ZN(n103) );
  NAND3_X1 U213 ( .A1(net75726), .A2(n103), .A3(net84131), .ZN(net84105) );
  NAND2_X2 U214 ( .A1(A[44]), .A2(B[44]), .ZN(net75726) );
  NAND2_X1 U215 ( .A1(net75846), .A2(net84123), .ZN(net84129) );
  BUF_X1 U216 ( .A(net75846), .Z(net75844) );
  INV_X2 U217 ( .A(A[44]), .ZN(net75720) );
  XNOR2_X2 U218 ( .A(A[44]), .B(B[44]), .ZN(net75759) );
  INV_X2 U219 ( .A(B[44]), .ZN(net75718) );
  OAI21_X1 U220 ( .B1(net82410), .B2(n108), .A(n109), .ZN(net82409) );
  NOR2_X2 U221 ( .A1(n104), .A2(net82338), .ZN(n106) );
  INV_X2 U222 ( .A(net70489), .ZN(n104) );
  NAND2_X1 U223 ( .A1(net82439), .A2(n111), .ZN(net82429) );
  NOR2_X1 U224 ( .A1(net82383), .A2(n3), .ZN(net82385) );
  AND2_X2 U225 ( .A1(A[12]), .A2(net69130), .ZN(net70489) );
  NAND2_X1 U226 ( .A1(net70464), .A2(net70489), .ZN(net70527) );
  INV_X2 U227 ( .A(net69110), .ZN(net69130) );
  NAND2_X1 U228 ( .A1(net69126), .A2(net69130), .ZN(net69117) );
  AND2_X2 U229 ( .A1(net69130), .A2(B[12]), .ZN(net70488) );
  NAND2_X2 U230 ( .A1(net82377), .A2(A[10]), .ZN(n105) );
  AND2_X2 U231 ( .A1(net73525), .A2(net73526), .ZN(net82523) );
  BUF_X1 U232 ( .A(n64), .Z(net82504) );
  NAND2_X2 U233 ( .A1(net73518), .A2(net56025), .ZN(net82375) );
  NOR2_X1 U234 ( .A1(net82508), .A2(net82375), .ZN(net82333) );
  NAND2_X1 U235 ( .A1(n116), .A2(B[19]), .ZN(net57091) );
  NAND2_X1 U236 ( .A1(n116), .A2(B[19]), .ZN(net55962) );
  BUF_X1 U237 ( .A(n116), .Z(net57085) );
  NAND2_X1 U238 ( .A1(\carry[18] ), .A2(A[18]), .ZN(n114) );
  NAND2_X1 U239 ( .A1(n117), .A2(B[18]), .ZN(net56888) );
  NAND2_X1 U240 ( .A1(B[18]), .A2(A[18]), .ZN(n115) );
  NAND3_X1 U241 ( .A1(net67465), .A2(n120), .A3(n115), .ZN(\carry[19] ) );
  NAND3_X1 U242 ( .A1(n119), .A2(net67462), .A3(n112), .ZN(\carry[18] ) );
  NAND2_X1 U243 ( .A1(\carry[18] ), .A2(A[18]), .ZN(n120) );
  NAND2_X1 U244 ( .A1(n60), .A2(A[17]), .ZN(net67462) );
  NAND2_X1 U245 ( .A1(n121), .A2(B[17]), .ZN(n119) );
  NAND2_X1 U246 ( .A1(net67421), .A2(net67379), .ZN(n121) );
  XOR2_X1 U247 ( .A(B[18]), .B(A[18]), .Z(net56887) );
  NAND3_X1 U248 ( .A1(n4), .A2(n113), .A3(n112), .ZN(n117) );
  NAND2_X1 U249 ( .A1(n10), .A2(B[18]), .ZN(net67465) );
  BUF_X1 U250 ( .A(n10), .Z(net57100) );
  NAND2_X1 U251 ( .A1(net67421), .A2(net67379), .ZN(n118) );
  NAND2_X1 U252 ( .A1(\carry[17] ), .A2(A[17]), .ZN(n113) );
  NAND2_X1 U253 ( .A1(A[17]), .A2(B[17]), .ZN(n112) );
  XOR2_X1 U254 ( .A(A[17]), .B(B[17]), .Z(net55603) );
  AND2_X2 U255 ( .A1(n127), .A2(n126), .ZN(net67421) );
  INV_X1 U256 ( .A(n123), .ZN(n126) );
  AND2_X2 U257 ( .A1(net67385), .A2(n126), .ZN(net67359) );
  OAI21_X1 U258 ( .B1(n124), .B2(net67355), .A(n125), .ZN(n123) );
  NAND2_X2 U259 ( .A1(B[16]), .A2(A[16]), .ZN(n125) );
  INV_X2 U260 ( .A(net67373), .ZN(n124) );
  NAND2_X1 U261 ( .A1(net55937), .A2(n128), .ZN(n127) );
  INV_X2 U262 ( .A(n122), .ZN(n128) );
  NAND2_X1 U263 ( .A1(net67466), .A2(n128), .ZN(net67360) );
  NAND2_X2 U264 ( .A1(net67373), .A2(B[15]), .ZN(n122) );
  NAND3_X1 U265 ( .A1(net67456), .A2(net69188), .A3(net55837), .ZN(net55937)
         );
  NAND2_X1 U266 ( .A1(net69072), .A2(A[14]), .ZN(net67456) );
  AOI21_X1 U267 ( .B1(net70460), .B2(n129), .A(net70458), .ZN(net69072) );
  INV_X2 U268 ( .A(net70443), .ZN(net70458) );
  AOI21_X1 U269 ( .B1(net82565), .B2(n129), .A(net70458), .ZN(net82522) );
  INV_X2 U270 ( .A(net70482), .ZN(n129) );
  NOR2_X2 U271 ( .A1(net70483), .A2(n129), .ZN(net70465) );
  NAND3_X1 U272 ( .A1(n137), .A2(n134), .A3(net56144), .ZN(n132) );
  NAND2_X1 U273 ( .A1(n132), .A2(B[54]), .ZN(net55819) );
  NAND2_X1 U274 ( .A1(n132), .A2(B[54]), .ZN(net73524) );
  BUF_X1 U275 ( .A(n132), .Z(net57004) );
  NAND2_X1 U276 ( .A1(\carry[53] ), .A2(B[53]), .ZN(n137) );
  NAND3_X1 U277 ( .A1(n53), .A2(n134), .A3(net56144), .ZN(net56431) );
  NAND3_X1 U278 ( .A1(net56855), .A2(net58289), .A3(net56140), .ZN(\carry[53] ) );
  INV_X1 U279 ( .A(net58320), .ZN(net58289) );
  OAI211_X1 U280 ( .C1(net58064), .C2(net58061), .A(n135), .B(net58449), .ZN(
        net58320) );
  NAND2_X1 U281 ( .A1(net79896), .A2(net58206), .ZN(n135) );
  INV_X2 U282 ( .A(net58069), .ZN(net58064) );
  OAI211_X1 U283 ( .C1(net58064), .C2(net58061), .A(net58321), .B(net58066), 
        .ZN(net58063) );
  OAI21_X2 U284 ( .B1(n133), .B2(net58040), .A(A[52]), .ZN(net56855) );
  NAND2_X1 U285 ( .A1(net58060), .A2(net58057), .ZN(n133) );
  NOR2_X2 U286 ( .A1(n136), .A2(net58450), .ZN(net58060) );
  INV_X32 U287 ( .A(net58242), .ZN(net58450) );
  NOR2_X1 U288 ( .A1(net58244), .A2(net58329), .ZN(n136) );
  INV_X2 U289 ( .A(net58424), .ZN(net58326) );
  NAND2_X1 U290 ( .A1(net79896), .A2(net58326), .ZN(net58059) );
  NAND2_X2 U291 ( .A1(B[50]), .A2(net58054), .ZN(net58424) );
  NAND2_X1 U292 ( .A1(n131), .A2(A[53]), .ZN(n134) );
  NAND3_X1 U293 ( .A1(net56142), .A2(n130), .A3(net56140), .ZN(n131) );
  INV_X1 U294 ( .A(net58063), .ZN(net56142) );
  BUF_X1 U295 ( .A(net56142), .Z(net58292) );
  NAND2_X1 U296 ( .A1(net56147), .A2(net58206), .ZN(net58066) );
  NAND2_X1 U297 ( .A1(net56817), .A2(A[52]), .ZN(n130) );
  NAND3_X1 U298 ( .A1(n140), .A2(n139), .A3(n138), .ZN(n141) );
  NAND2_X1 U299 ( .A1(n141), .A2(B[58]), .ZN(net56549) );
  NAND2_X1 U300 ( .A1(n141), .A2(B[58]), .ZN(net56261) );
  BUF_X1 U301 ( .A(n141), .Z(net56400) );
  NAND2_X1 U302 ( .A1(n9), .A2(B[57]), .ZN(n140) );
  NAND3_X1 U303 ( .A1(n139), .A2(n138), .A3(n140), .ZN(\carry[58] ) );
  NAND2_X1 U304 ( .A1(\carry[57] ), .A2(A[57]), .ZN(n139) );
  NAND2_X1 U305 ( .A1(A[57]), .A2(B[57]), .ZN(n138) );
  XOR2_X1 U306 ( .A(A[57]), .B(B[57]), .Z(net55571) );
  INV_X1 U307 ( .A(net73517), .ZN(net82542) );
  AND2_X1 U308 ( .A1(n144), .A2(B[9]), .ZN(n145) );
  NAND3_X1 U309 ( .A1(net56755), .A2(net73488), .A3(net73487), .ZN(n146) );
  BUF_X1 U310 ( .A(n146), .Z(net73656) );
  NAND2_X2 U311 ( .A1(n143), .A2(n142), .ZN(n144) );
  AND2_X1 U312 ( .A1(n144), .A2(A[9]), .ZN(net77818) );
  NAND2_X1 U313 ( .A1(net73656), .A2(n144), .ZN(net73473) );
  AND2_X1 U314 ( .A1(n144), .A2(A[9]), .ZN(net73528) );
  NAND2_X2 U315 ( .A1(net73491), .A2(A[7]), .ZN(n142) );
  NAND2_X2 U316 ( .A1(net73491), .A2(B[7]), .ZN(n143) );
  INV_X1 U317 ( .A(B[9]), .ZN(net73519) );
  NAND2_X1 U318 ( .A1(B[9]), .A2(A[9]), .ZN(net56025) );
  XOR2_X1 U319 ( .A(B[9]), .B(A[9]), .Z(net56022) );
  NAND3_X1 U320 ( .A1(net56755), .A2(net73488), .A3(net73487), .ZN(net56793)
         );
  AOI21_X2 U321 ( .B1(net73490), .B2(net73491), .A(net73492), .ZN(net73472) );
  NAND2_X2 U322 ( .A1(A[7]), .A2(B[7]), .ZN(net73468) );
  NOR2_X2 U323 ( .A1(A[7]), .A2(B[7]), .ZN(net73489) );
  INV_X1 U324 ( .A(net82409), .ZN(net69119) );
  INV_X1 U325 ( .A(net82378), .ZN(net82384) );
  NAND2_X1 U326 ( .A1(net82377), .A2(B[10]), .ZN(net82378) );
  INV_X1 U327 ( .A(net82412), .ZN(net82410) );
  AND3_X2 U328 ( .A1(net84166), .A2(net84167), .A3(net56333), .ZN(net75846) );
  NAND2_X2 U329 ( .A1(n147), .A2(B[52]), .ZN(net58061) );
  NAND2_X2 U330 ( .A1(net58056), .A2(net56041), .ZN(n147) );
  AND3_X2 U331 ( .A1(A[50]), .A2(B[52]), .A3(net58069), .ZN(net58206) );
  AND3_X2 U332 ( .A1(B[50]), .A2(B[52]), .A3(net58069), .ZN(net58409) );
  NAND2_X2 U333 ( .A1(net58055), .A2(net58056), .ZN(net58069) );
  INV_X2 U334 ( .A(net58054), .ZN(net58055) );
  OAI21_X2 U335 ( .B1(net58055), .B2(net56041), .A(net58056), .ZN(net58040) );
  NAND2_X1 U336 ( .A1(\carry[32] ), .A2(B[32]), .ZN(net59537) );
  INV_X2 U337 ( .A(net65693), .ZN(net65659) );
  AOI21_X1 U338 ( .B1(net65658), .B2(net69164), .A(net65659), .ZN(net65638) );
  AOI21_X1 U339 ( .B1(net65685), .B2(net65697), .A(net65659), .ZN(net65637) );
  INV_X2 U340 ( .A(net65679), .ZN(net65691) );
  INV_X1 U341 ( .A(net65709), .ZN(net65697) );
  BUF_X1 U342 ( .A(net65697), .Z(net69164) );
  NAND2_X2 U343 ( .A1(B[31]), .A2(A[31]), .ZN(net65677) );
  NAND2_X2 U344 ( .A1(A[32]), .A2(net65679), .ZN(net65680) );
  INV_X2 U345 ( .A(A[31]), .ZN(net65671) );
  AND2_X2 U346 ( .A1(net57011), .A2(B[30]), .ZN(net65709) );
  AOI21_X2 U347 ( .B1(net65709), .B2(net65687), .A(net65678), .ZN(net65686) );
  XNOR2_X2 U348 ( .A(B[31]), .B(A[31]), .ZN(net59519) );
  BUF_X1 U349 ( .A(net57011), .Z(net56468) );
  NAND2_X2 U350 ( .A1(n149), .A2(net60770), .ZN(net62307) );
  NOR2_X1 U351 ( .A1(net69202), .A2(net62307), .ZN(net62273) );
  NOR2_X2 U352 ( .A1(n148), .A2(net62326), .ZN(n149) );
  INV_X2 U353 ( .A(B[24]), .ZN(net62326) );
  NOR2_X2 U354 ( .A1(B[22]), .A2(A[22]), .ZN(n148) );
  NAND2_X1 U355 ( .A1(net56569), .A2(B[21]), .ZN(net62344) );
  NAND3_X1 U356 ( .A1(net55966), .A2(net55965), .A3(net55964), .ZN(net56569)
         );
  NAND2_X1 U357 ( .A1(n152), .A2(A[21]), .ZN(net56054) );
  NAND2_X2 U358 ( .A1(A[21]), .A2(B[21]), .ZN(net62332) );
  AND3_X1 U359 ( .A1(n150), .A2(n151), .A3(net62332), .ZN(net62289) );
  AND3_X2 U360 ( .A1(n150), .A2(net56054), .A3(net62332), .ZN(net69202) );
  AND2_X2 U361 ( .A1(net60770), .A2(B[24]), .ZN(net62309) );
  NAND2_X1 U362 ( .A1(net65234), .A2(B[21]), .ZN(n150) );
  XNOR2_X2 U363 ( .A(A[21]), .B(B[21]), .ZN(net60821) );
  NAND3_X1 U364 ( .A1(net55966), .A2(net55965), .A3(net55964), .ZN(net65234)
         );
  NAND3_X1 U365 ( .A1(net56901), .A2(net57089), .A3(net55964), .ZN(n152) );
  NAND2_X1 U366 ( .A1(n152), .A2(A[21]), .ZN(n151) );
  AOI21_X1 U367 ( .B1(n154), .B2(n155), .A(n153), .ZN(net57019) );
  NAND2_X1 U368 ( .A1(net57019), .A2(A[38]), .ZN(net65272) );
  INV_X2 U369 ( .A(n157), .ZN(n153) );
  NAND2_X2 U370 ( .A1(net65153), .A2(n156), .ZN(n157) );
  INV_X2 U371 ( .A(net64019), .ZN(n156) );
  NAND2_X2 U372 ( .A1(net64012), .A2(net64010), .ZN(net64019) );
  NAND2_X2 U373 ( .A1(net64012), .A2(net64010), .ZN(net65192) );
  NAND2_X1 U374 ( .A1(n159), .A2(net65221), .ZN(n155) );
  INV_X2 U375 ( .A(net65191), .ZN(net65221) );
  NAND2_X1 U376 ( .A1(net73570), .A2(net73663), .ZN(n159) );
  AND2_X1 U377 ( .A1(net73562), .A2(net73561), .ZN(net73663) );
  AND2_X2 U378 ( .A1(net73562), .A2(net73561), .ZN(net62117) );
  NAND2_X1 U379 ( .A1(net73554), .A2(n158), .ZN(n154) );
  OR2_X1 U380 ( .A1(net65199), .A2(net65196), .ZN(n158) );
  INV_X1 U381 ( .A(net65199), .ZN(net73557) );
  INV_X2 U382 ( .A(B[43]), .ZN(net84109) );
  AND2_X2 U383 ( .A1(n47), .A2(net84122), .ZN(n162) );
  INV_X2 U384 ( .A(net75699), .ZN(n163) );
  INV_X2 U385 ( .A(net57080), .ZN(net84131) );
  NAND2_X2 U386 ( .A1(A[43]), .A2(B[43]), .ZN(n160) );
  NAND2_X2 U387 ( .A1(A[43]), .A2(n163), .ZN(n161) );
  NAND2_X2 U388 ( .A1(A[43]), .A2(B[43]), .ZN(n164) );
  NAND4_X1 U389 ( .A1(n55), .A2(n164), .A3(n59), .A4(net56333), .ZN(net84135)
         );
  AND3_X2 U390 ( .A1(net75734), .A2(net84129), .A3(net84122), .ZN(net75678) );
  AND3_X2 U391 ( .A1(net56335), .A2(net56334), .A3(net56333), .ZN(n165) );
  BUF_X1 U392 ( .A(n55), .Z(n166) );
  NAND2_X1 U393 ( .A1(n165), .A2(net84099), .ZN(net75734) );
  NAND3_X1 U394 ( .A1(n178), .A2(net79844), .A3(n168), .ZN(n167) );
  NAND2_X1 U395 ( .A1(\carry[39] ), .A2(A[39]), .ZN(n168) );
  NAND2_X2 U396 ( .A1(n169), .A2(n170), .ZN(net70464) );
  AND4_X2 U397 ( .A1(n190), .A2(n189), .A3(n191), .A4(net82338), .ZN(n169) );
  AND3_X2 U398 ( .A1(net82391), .A2(n192), .A3(n193), .ZN(n170) );
  AND3_X1 U399 ( .A1(n185), .A2(n184), .A3(n183), .ZN(net82565) );
  NAND3_X1 U400 ( .A1(net55819), .A2(n376), .A3(n375), .ZN(n171) );
  NAND2_X1 U401 ( .A1(net82384), .A2(n172), .ZN(n189) );
  NAND2_X1 U402 ( .A1(n240), .A2(n241), .ZN(n172) );
  NAND2_X1 U403 ( .A1(n207), .A2(B[27]), .ZN(n173) );
  NAND2_X1 U404 ( .A1(\carry[27] ), .A2(A[27]), .ZN(n174) );
  NAND2_X1 U405 ( .A1(net82522), .A2(A[14]), .ZN(n175) );
  NOR2_X1 U406 ( .A1(net60799), .A2(net60800), .ZN(net82516) );
  NOR2_X1 U407 ( .A1(net60799), .A2(net60800), .ZN(net60886) );
  NAND3_X1 U408 ( .A1(net79914), .A2(net56370), .A3(net56371), .ZN(net82512)
         );
  AND2_X2 U409 ( .A1(n240), .A2(n241), .ZN(net82510) );
  BUF_X1 U410 ( .A(net82542), .Z(net82508) );
  NAND2_X1 U411 ( .A1(net73525), .A2(net73526), .ZN(n176) );
  NAND2_X1 U412 ( .A1(net82542), .A2(net82384), .ZN(n190) );
  NAND2_X1 U413 ( .A1(net82542), .A2(net82423), .ZN(n193) );
  NAND2_X1 U414 ( .A1(n176), .A2(net82423), .ZN(n191) );
  NAND2_X1 U415 ( .A1(n176), .A2(net82394), .ZN(n194) );
  NAND2_X1 U416 ( .A1(net82333), .A2(net82504), .ZN(net77826) );
  NAND2_X1 U417 ( .A1(\carry[39] ), .A2(A[39]), .ZN(n177) );
  BUF_X1 U418 ( .A(net67360), .Z(net82494) );
  NAND2_X1 U419 ( .A1(net56856), .A2(B[39]), .ZN(n178) );
  NAND2_X1 U420 ( .A1(\carry[28] ), .A2(B[28]), .ZN(n179) );
  AOI21_X1 U421 ( .B1(net82405), .B2(net82402), .A(n186), .ZN(n197) );
  NAND2_X1 U422 ( .A1(net82427), .A2(n172), .ZN(n184) );
  AOI21_X2 U423 ( .B1(net70464), .B2(n271), .A(net70465), .ZN(net55836) );
  INV_X2 U424 ( .A(B[10]), .ZN(net82363) );
  INV_X2 U425 ( .A(A[11]), .ZN(net82365) );
  INV_X2 U426 ( .A(B[11]), .ZN(net82367) );
  INV_X2 U427 ( .A(net70500), .ZN(net82369) );
  INV_X2 U428 ( .A(net70488), .ZN(net82373) );
  NOR2_X2 U429 ( .A1(net82373), .A2(net82338), .ZN(n186) );
  NAND2_X2 U430 ( .A1(n187), .A2(net73518), .ZN(net82381) );
  NOR2_X2 U431 ( .A1(net82383), .A2(net82387), .ZN(n188) );
  NOR2_X2 U432 ( .A1(A[10]), .A2(net82355), .ZN(n187) );
  NAND3_X1 U433 ( .A1(n215), .A2(n206), .A3(n205), .ZN(n208) );
  NAND2_X1 U434 ( .A1(n208), .A2(B[29]), .ZN(net62177) );
  BUF_X1 U435 ( .A(n208), .Z(net56209) );
  NAND2_X1 U436 ( .A1(n209), .A2(A[28]), .ZN(n206) );
  NAND3_X1 U437 ( .A1(n174), .A2(n173), .A3(n204), .ZN(n209) );
  NAND2_X1 U438 ( .A1(\carry[28] ), .A2(B[28]), .ZN(n215) );
  NAND3_X1 U439 ( .A1(n210), .A2(n179), .A3(n205), .ZN(\carry[29] ) );
  NAND3_X1 U440 ( .A1(n211), .A2(n214), .A3(n204), .ZN(\carry[28] ) );
  NAND2_X1 U441 ( .A1(n217), .A2(A[27]), .ZN(n214) );
  NAND3_X1 U442 ( .A1(net57097), .A2(net60856), .A3(net55592), .ZN(n217) );
  NAND2_X1 U443 ( .A1(n213), .A2(B[27]), .ZN(n211) );
  NAND2_X1 U444 ( .A1(A[28]), .A2(B[28]), .ZN(n205) );
  XOR2_X1 U445 ( .A(A[28]), .B(B[28]), .Z(net56060) );
  NAND2_X1 U446 ( .A1(net62212), .A2(A[28]), .ZN(n210) );
  NAND2_X1 U447 ( .A1(\carry[27] ), .A2(A[27]), .ZN(n212) );
  NAND3_X1 U448 ( .A1(n212), .A2(n216), .A3(n204), .ZN(net62212) );
  NAND3_X1 U449 ( .A1(net57097), .A2(net60856), .A3(net55592), .ZN(\carry[27] ) );
  NAND2_X1 U450 ( .A1(n207), .A2(B[27]), .ZN(n216) );
  NAND3_X1 U451 ( .A1(net73589), .A2(n68), .A3(net55592), .ZN(n207) );
  NAND2_X1 U452 ( .A1(A[27]), .A2(B[27]), .ZN(n204) );
  XOR2_X1 U453 ( .A(A[27]), .B(B[27]), .Z(net55595) );
  NAND3_X1 U454 ( .A1(net73589), .A2(n68), .A3(net55592), .ZN(n213) );
  BUF_X1 U455 ( .A(n213), .Z(net55673) );
  NAND2_X1 U456 ( .A1(net70524), .A2(n218), .ZN(net67379) );
  AND2_X1 U457 ( .A1(A[15]), .A2(net67373), .ZN(n218) );
  NAND2_X1 U458 ( .A1(net67359), .A2(net67360), .ZN(\carry[17] ) );
  XNOR2_X2 U459 ( .A(B[16]), .B(A[16]), .ZN(net67389) );
  INV_X2 U460 ( .A(B[16]), .ZN(net67370) );
  NAND2_X1 U461 ( .A1(net73577), .A2(net79856), .ZN(net79933) );
  BUF_X1 U462 ( .A(n48), .Z(net56744) );
  NAND2_X1 U463 ( .A1(net56856), .A2(B[39]), .ZN(n228) );
  NAND3_X1 U464 ( .A1(n178), .A2(n168), .A3(net79844), .ZN(net79836) );
  NAND3_X1 U465 ( .A1(net65272), .A2(n219), .A3(net56739), .ZN(\carry[39] ) );
  NAND2_X1 U466 ( .A1(net64058), .A2(B[38]), .ZN(n219) );
  AOI21_X1 U467 ( .B1(n220), .B2(n221), .A(n222), .ZN(net64058) );
  NAND2_X2 U468 ( .A1(net65215), .A2(net65153), .ZN(n223) );
  NAND2_X1 U469 ( .A1(net73564), .A2(n224), .ZN(n221) );
  OR2_X1 U470 ( .A1(net73566), .A2(net65196), .ZN(n224) );
  INV_X1 U471 ( .A(net65153), .ZN(net73566) );
  NAND2_X1 U472 ( .A1(n225), .A2(n226), .ZN(n220) );
  OR2_X1 U473 ( .A1(n227), .A2(net65221), .ZN(n226) );
  INV_X1 U474 ( .A(net65188), .ZN(n227) );
  NAND2_X1 U475 ( .A1(net62117), .A2(net73675), .ZN(n225) );
  NAND2_X1 U476 ( .A1(net57103), .A2(B[42]), .ZN(net56335) );
  NAND2_X1 U477 ( .A1(n229), .A2(A[42]), .ZN(net56334) );
  NAND2_X1 U478 ( .A1(A[42]), .A2(B[42]), .ZN(net56333) );
  XOR2_X1 U479 ( .A(A[42]), .B(B[42]), .Z(net56332) );
  NAND3_X1 U480 ( .A1(net79904), .A2(net56370), .A3(net56371), .ZN(n229) );
  NAND3_X1 U481 ( .A1(net56791), .A2(net56371), .A3(net57061), .ZN(net56427)
         );
  AND2_X2 U482 ( .A1(n230), .A2(net79928), .ZN(net56370) );
  NAND2_X1 U483 ( .A1(n167), .A2(net79930), .ZN(n230) );
  INV_X1 U484 ( .A(A[41]), .ZN(net79929) );
  BUF_X1 U485 ( .A(net56630), .Z(net79893) );
  BUF_X1 U486 ( .A(net56856), .Z(net79866) );
  INV_X2 U487 ( .A(A[40]), .ZN(n231) );
  INV_X2 U488 ( .A(B[40]), .ZN(n232) );
  NAND2_X2 U489 ( .A1(A[40]), .A2(B[40]), .ZN(net79832) );
  NAND2_X2 U490 ( .A1(B[41]), .A2(A[40]), .ZN(n233) );
  NAND2_X2 U491 ( .A1(B[41]), .A2(B[40]), .ZN(n234) );
  NAND2_X2 U492 ( .A1(net79851), .A2(B[41]), .ZN(net79849) );
  NAND2_X2 U493 ( .A1(n232), .A2(n231), .ZN(net79855) );
  NAND2_X2 U494 ( .A1(n234), .A2(n233), .ZN(net79856) );
  XNOR2_X2 U495 ( .A(A[39]), .B(B[39]), .ZN(n235) );
  INV_X2 U496 ( .A(n235), .ZN(net56639) );
  XNOR2_X2 U497 ( .A(A[40]), .B(B[40]), .ZN(n236) );
  INV_X2 U498 ( .A(n236), .ZN(net56562) );
  NAND2_X1 U499 ( .A1(n237), .A2(net58059), .ZN(net56817) );
  AND2_X2 U500 ( .A1(net58447), .A2(n238), .ZN(n237) );
  AND2_X1 U501 ( .A1(net58038), .A2(net58242), .ZN(n238) );
  INV_X2 U502 ( .A(net58040), .ZN(net58038) );
  NAND2_X1 U503 ( .A1(net58037), .A2(net58038), .ZN(net58121) );
  NAND2_X1 U504 ( .A1(A[53]), .A2(B[53]), .ZN(net56144) );
  BUF_X1 U505 ( .A(net79896), .Z(net58351) );
  INV_X2 U506 ( .A(B[50]), .ZN(net58405) );
  AND2_X2 U507 ( .A1(net77768), .A2(n243), .ZN(n239) );
  NAND2_X1 U508 ( .A1(net56793), .A2(net77818), .ZN(n240) );
  OR2_X1 U509 ( .A1(net77817), .A2(net73472), .ZN(n241) );
  INV_X1 U510 ( .A(A[9]), .ZN(net77817) );
  AND2_X2 U511 ( .A1(A[2]), .A2(A[3]), .ZN(net77766) );
  INV_X2 U512 ( .A(net77785), .ZN(net55812) );
  INV_X2 U513 ( .A(n244), .ZN(net55808) );
  XNOR2_X1 U514 ( .A(net77806), .B(net77831), .ZN(n244) );
  NOR2_X1 U515 ( .A1(\carry[1] ), .A2(net77806), .ZN(n242) );
  OAI21_X1 U516 ( .B1(net77748), .B2(n242), .A(net56561), .ZN(net56545) );
  BUF_X1 U517 ( .A(\carry[1] ), .Z(net57059) );
  NAND2_X1 U518 ( .A1(net77765), .A2(net77776), .ZN(n243) );
  NAND3_X1 U519 ( .A1(n246), .A2(n247), .A3(n245), .ZN(net56859) );
  NAND2_X1 U520 ( .A1(net56859), .A2(B[48]), .ZN(net58227) );
  BUF_X1 U521 ( .A(n6), .Z(net56883) );
  NAND2_X1 U522 ( .A1(n61), .A2(B[47]), .ZN(n247) );
  NAND3_X1 U523 ( .A1(n8), .A2(n54), .A3(n245), .ZN(\carry[48] ) );
  NAND2_X1 U524 ( .A1(\carry[47] ), .A2(A[47]), .ZN(n246) );
  NAND2_X1 U525 ( .A1(A[47]), .A2(B[47]), .ZN(n245) );
  XOR2_X1 U526 ( .A(A[47]), .B(B[47]), .Z(net55579) );
  BUF_X1 U527 ( .A(net75678), .Z(net75842) );
  NOR2_X1 U528 ( .A1(net65684), .A2(net65683), .ZN(n248) );
  NOR2_X1 U529 ( .A1(n7), .A2(net65683), .ZN(net65688) );
  NAND2_X1 U530 ( .A1(net75842), .A2(A[45]), .ZN(n249) );
  INV_X1 U531 ( .A(net75844), .ZN(net57080) );
  NAND2_X2 U532 ( .A1(n250), .A2(net75725), .ZN(net75723) );
  INV_X2 U533 ( .A(net75743), .ZN(net57069) );
  NAND2_X2 U534 ( .A1(net75720), .A2(net75718), .ZN(n250) );
  INV_X2 U535 ( .A(net75759), .ZN(net55822) );
  NOR2_X1 U536 ( .A1(net75831), .A2(B[43]), .ZN(net75699) );
  AND2_X2 U537 ( .A1(net70524), .A2(A[15]), .ZN(net67433) );
  AND2_X1 U538 ( .A1(net67373), .A2(A[15]), .ZN(net67429) );
  XOR2_X1 U539 ( .A(B[41]), .B(A[41]), .Z(net56368) );
  AND2_X2 U540 ( .A1(n248), .A2(net65686), .ZN(net59538) );
  AND2_X1 U541 ( .A1(net65686), .A2(net65688), .ZN(net73660) );
  INV_X2 U542 ( .A(A[32]), .ZN(net65675) );
  INV_X2 U543 ( .A(net65680), .ZN(net65687) );
  XOR2_X1 U544 ( .A(A[32]), .B(B[32]), .Z(net56044) );
  NAND2_X1 U545 ( .A1(A[32]), .A2(B[32]), .ZN(net56045) );
  NAND2_X2 U546 ( .A1(net65181), .A2(net65179), .ZN(net65183) );
  AND2_X2 U547 ( .A1(net73570), .A2(net65188), .ZN(net73675) );
  NAND3_X1 U548 ( .A1(n313), .A2(net60691), .A3(n386), .ZN(n251) );
  INV_X1 U549 ( .A(net73494), .ZN(net73634) );
  BUF_X1 U550 ( .A(n284), .Z(n252) );
  AND2_X1 U551 ( .A1(net56739), .A2(n292), .ZN(n253) );
  NAND2_X1 U552 ( .A1(net65219), .A2(net65225), .ZN(n292) );
  NAND3_X1 U553 ( .A1(net62205), .A2(n239), .A3(n346), .ZN(n254) );
  NAND3_X1 U554 ( .A1(net62205), .A2(n239), .A3(n346), .ZN(n343) );
  NAND2_X1 U555 ( .A1(n251), .A2(A[26]), .ZN(net73589) );
  NAND3_X1 U556 ( .A1(net73660), .A2(net56047), .A3(net56045), .ZN(n255) );
  BUF_X1 U557 ( .A(net56341), .Z(n256) );
  AND2_X1 U558 ( .A1(net73669), .A2(net65196), .ZN(n266) );
  NAND2_X1 U559 ( .A1(net65196), .A2(net73669), .ZN(n257) );
  NAND2_X1 U560 ( .A1(n284), .A2(net62140), .ZN(net73570) );
  NAND2_X1 U561 ( .A1(n268), .A2(n267), .ZN(net73562) );
  NAND3_X1 U562 ( .A1(n332), .A2(n331), .A3(n330), .ZN(n258) );
  NAND2_X1 U563 ( .A1(n254), .A2(B[4]), .ZN(n259) );
  NAND3_X1 U564 ( .A1(n332), .A2(n330), .A3(n331), .ZN(\carry[6] ) );
  NAND2_X1 U565 ( .A1(net70464), .A2(net70488), .ZN(n260) );
  NAND2_X1 U566 ( .A1(net56793), .A2(net73528), .ZN(net73525) );
  OR2_X1 U567 ( .A1(net73527), .A2(net73472), .ZN(net73526) );
  INV_X1 U568 ( .A(A[9]), .ZN(net73527) );
  BUF_X1 U569 ( .A(n258), .Z(n261) );
  OR2_X1 U570 ( .A1(net73519), .A2(net73472), .ZN(net73518) );
  NAND2_X1 U571 ( .A1(net73473), .A2(net73472), .ZN(net56341) );
  INV_X1 U572 ( .A(net73656), .ZN(net73494) );
  NAND2_X1 U573 ( .A1(\carry[6] ), .A2(B[6]), .ZN(net73488) );
  INV_X2 U574 ( .A(A[8]), .ZN(n263) );
  XNOR2_X2 U575 ( .A(A[8]), .B(B[8]), .ZN(net72085) );
  INV_X2 U576 ( .A(n264), .ZN(net72097) );
  NAND2_X2 U577 ( .A1(n263), .A2(n262), .ZN(net73491) );
  NAND2_X2 U578 ( .A1(A[8]), .A2(B[8]), .ZN(net73498) );
  INV_X2 U579 ( .A(net73498), .ZN(net73492) );
  NAND2_X2 U580 ( .A1(A[6]), .A2(B[6]), .ZN(net73487) );
  XNOR2_X2 U581 ( .A(B[6]), .B(A[6]), .ZN(n265) );
  NAND2_X1 U582 ( .A1(net62117), .A2(net73570), .ZN(net65288) );
  BUF_X1 U583 ( .A(net65288), .Z(net65124) );
  INV_X2 U584 ( .A(B[35]), .ZN(net65179) );
  INV_X2 U585 ( .A(A[35]), .ZN(net65181) );
  BUF_X1 U586 ( .A(n266), .Z(net65299) );
  INV_X32 U587 ( .A(n295), .ZN(n267) );
  NAND3_X1 U588 ( .A1(net59537), .A2(net59538), .A3(net56045), .ZN(n268) );
  NAND2_X1 U589 ( .A1(net65637), .A2(B[32]), .ZN(net56047) );
  INV_X2 U590 ( .A(net72085), .ZN(net56313) );
  INV_X2 U591 ( .A(net72087), .ZN(net56309) );
  INV_X2 U592 ( .A(net72097), .ZN(net56366) );
  AND3_X2 U593 ( .A1(n260), .A2(net70527), .A3(n278), .ZN(n269) );
  NAND3_X1 U594 ( .A1(n269), .A2(net55836), .A3(net55837), .ZN(net70524) );
  INV_X2 U595 ( .A(A[12]), .ZN(net70474) );
  INV_X2 U596 ( .A(B[13]), .ZN(n272) );
  INV_X2 U597 ( .A(A[13]), .ZN(n273) );
  INV_X2 U598 ( .A(B[12]), .ZN(net70480) );
  NAND2_X2 U599 ( .A1(net69089), .A2(n270), .ZN(net70482) );
  NAND2_X2 U600 ( .A1(A[14]), .A2(net70443), .ZN(net70483) );
  NOR2_X2 U601 ( .A1(net70483), .A2(net70480), .ZN(n274) );
  NOR2_X2 U602 ( .A1(net70487), .A2(net70474), .ZN(net69139) );
  NAND2_X2 U603 ( .A1(net69089), .A2(n270), .ZN(n275) );
  AOI21_X2 U604 ( .B1(A[12]), .B2(net56481), .A(n275), .ZN(net70456) );
  NAND2_X2 U605 ( .A1(A[13]), .A2(B[13]), .ZN(n270) );
  INV_X2 U606 ( .A(n270), .ZN(net69124) );
  INV_X2 U607 ( .A(net56481), .ZN(net70487) );
  NAND2_X2 U608 ( .A1(n273), .A2(n272), .ZN(net70443) );
  INV_X2 U609 ( .A(net70483), .ZN(net70495) );
  NAND2_X2 U610 ( .A1(net70495), .A2(A[12]), .ZN(n276) );
  INV_X2 U611 ( .A(n274), .ZN(n277) );
  NAND2_X2 U612 ( .A1(n277), .A2(n276), .ZN(n271) );
  BUF_X1 U613 ( .A(net70464), .Z(net56481) );
  AND2_X1 U614 ( .A1(net69117), .A2(n280), .ZN(n278) );
  AND3_X2 U615 ( .A1(net69119), .A2(n69), .A3(n278), .ZN(net69188) );
  NAND2_X1 U616 ( .A1(net69124), .A2(B[14]), .ZN(n280) );
  INV_X1 U617 ( .A(net69139), .ZN(net55925) );
  NAND2_X2 U618 ( .A1(A[12]), .A2(B[12]), .ZN(net69089) );
  NAND2_X2 U619 ( .A1(net56481), .A2(B[12]), .ZN(n279) );
  INV_X2 U620 ( .A(net69089), .ZN(net69126) );
  INV_X2 U621 ( .A(net69132), .ZN(net55927) );
  XNOR2_X2 U622 ( .A(B[12]), .B(A[12]), .ZN(n281) );
  INV_X2 U623 ( .A(n281), .ZN(net55923) );
  NAND2_X1 U624 ( .A1(net56862), .A2(B[25]), .ZN(n282) );
  NAND3_X1 U625 ( .A1(n175), .A2(n269), .A3(net55837), .ZN(net67466) );
  NAND2_X1 U626 ( .A1(n252), .A2(A[33]), .ZN(n297) );
  BUF_X1 U627 ( .A(net67466), .Z(net67457) );
  NAND2_X1 U628 ( .A1(net67457), .A2(B[15]), .ZN(net67357) );
  BUF_X1 U629 ( .A(net67359), .Z(net67423) );
  INV_X2 U630 ( .A(A[16]), .ZN(net67368) );
  NAND2_X2 U631 ( .A1(A[15]), .A2(B[15]), .ZN(net67355) );
  NAND2_X2 U632 ( .A1(net67370), .A2(net67368), .ZN(net67373) );
  XNOR2_X2 U633 ( .A(A[15]), .B(B[15]), .ZN(n283) );
  INV_X2 U634 ( .A(n283), .ZN(net55691) );
  INV_X2 U635 ( .A(net67389), .ZN(net55599) );
  INV_X1 U636 ( .A(net67433), .ZN(net67391) );
  NAND2_X1 U637 ( .A1(\carry[15] ), .A2(net67429), .ZN(net67385) );
  NAND2_X1 U638 ( .A1(net67423), .A2(net82494), .ZN(net55674) );
  NAND3_X1 U639 ( .A1(net56047), .A2(net73660), .A3(net56045), .ZN(n284) );
  NAND2_X1 U640 ( .A1(n343), .A2(B[4]), .ZN(n285) );
  INV_X1 U641 ( .A(net65702), .ZN(net65704) );
  NAND2_X1 U642 ( .A1(net60796), .A2(net60854), .ZN(net65321) );
  NAND2_X1 U643 ( .A1(net69203), .A2(net60854), .ZN(net55832) );
  BUF_X1 U644 ( .A(n294), .Z(n286) );
  NAND2_X1 U645 ( .A1(net65221), .A2(net65124), .ZN(net65160) );
  NAND2_X1 U646 ( .A1(net65221), .A2(net65124), .ZN(n289) );
  NAND2_X1 U647 ( .A1(n291), .A2(n253), .ZN(net65309) );
  BUF_X1 U648 ( .A(n307), .Z(n287) );
  NAND2_X1 U649 ( .A1(A[35]), .A2(B[35]), .ZN(net65201) );
  AND3_X1 U650 ( .A1(net65188), .A2(n257), .A3(n289), .ZN(net64053) );
  NOR2_X1 U651 ( .A1(net65299), .A2(net65199), .ZN(net65159) );
  NAND2_X1 U652 ( .A1(net65290), .A2(net65272), .ZN(net56856) );
  NAND2_X2 U653 ( .A1(A[35]), .A2(B[35]), .ZN(n288) );
  NAND2_X2 U654 ( .A1(n290), .A2(A[36]), .ZN(net65188) );
  NAND2_X2 U655 ( .A1(net65188), .A2(net65153), .ZN(net65199) );
  INV_X2 U656 ( .A(n288), .ZN(n290) );
  INV_X2 U657 ( .A(net65188), .ZN(net65219) );
  NAND3_X1 U658 ( .A1(net65288), .A2(net65225), .A3(net65221), .ZN(n291) );
  XNOR2_X2 U659 ( .A(A[35]), .B(B[35]), .ZN(n293) );
  INV_X2 U660 ( .A(n293), .ZN(net55683) );
  BUF_X1 U661 ( .A(net65234), .Z(net56428) );
  BUF_X1 U662 ( .A(net65638), .Z(net56210) );
  BUF_X1 U663 ( .A(net65126), .Z(net64059) );
  NAND3_X1 U664 ( .A1(net59537), .A2(net59538), .A3(net56045), .ZN(n294) );
  NAND2_X1 U665 ( .A1(B[33]), .A2(n286), .ZN(net62110) );
  NAND2_X1 U666 ( .A1(n294), .A2(net62141), .ZN(net62138) );
  INV_X2 U667 ( .A(net64020), .ZN(net55587) );
  INV_X2 U668 ( .A(net64022), .ZN(net55583) );
  INV_X1 U669 ( .A(net64053), .ZN(net55672) );
  NAND2_X2 U670 ( .A1(net62130), .A2(B[33]), .ZN(n295) );
  INV_X2 U671 ( .A(n295), .ZN(net62141) );
  INV_X2 U672 ( .A(net62130), .ZN(net62132) );
  NAND2_X2 U673 ( .A1(net62130), .A2(A[33]), .ZN(net62129) );
  NAND2_X2 U674 ( .A1(B[33]), .A2(A[33]), .ZN(net62111) );
  XNOR2_X2 U675 ( .A(B[33]), .B(A[33]), .ZN(net62145) );
  INV_X2 U676 ( .A(net62338), .ZN(net55830) );
  BUF_X1 U677 ( .A(net62289), .Z(net62290) );
  BUF_X1 U678 ( .A(net58059), .Z(net62218) );
  NAND2_X1 U679 ( .A1(\carry[4] ), .A2(A[4]), .ZN(n296) );
  BUF_X1 U680 ( .A(net65124), .Z(net62200) );
  NOR2_X2 U681 ( .A1(net62273), .A2(net60800), .ZN(net60754) );
  NAND2_X1 U682 ( .A1(net57080), .A2(B[43]), .ZN(net62194) );
  NAND2_X1 U683 ( .A1(n255), .A2(net62140), .ZN(net62139) );
  INV_X1 U684 ( .A(net62290), .ZN(net56148) );
  OR2_X2 U685 ( .A1(net58329), .A2(net58244), .ZN(net58447) );
  INV_X2 U686 ( .A(B[34]), .ZN(n298) );
  INV_X2 U687 ( .A(A[34]), .ZN(n299) );
  OAI21_X2 U688 ( .B1(net62132), .B2(net62111), .A(n300), .ZN(net62131) );
  NAND2_X2 U689 ( .A1(n299), .A2(n298), .ZN(net62130) );
  NAND2_X2 U690 ( .A1(A[34]), .A2(B[34]), .ZN(n300) );
  INV_X2 U691 ( .A(net62129), .ZN(net62140) );
  INV_X2 U692 ( .A(net62145), .ZN(net56048) );
  XNOR2_X2 U693 ( .A(A[34]), .B(B[34]), .ZN(n301) );
  INV_X2 U694 ( .A(n301), .ZN(net55826) );
  NAND3_X1 U695 ( .A1(net55689), .A2(n282), .A3(n386), .ZN(n302) );
  NAND3_X1 U696 ( .A1(net55689), .A2(n385), .A3(n386), .ZN(n317) );
  NAND2_X1 U697 ( .A1(n251), .A2(A[26]), .ZN(net60856) );
  INV_X1 U698 ( .A(net60823), .ZN(net60835) );
  INV_X2 U699 ( .A(B[23]), .ZN(n303) );
  INV_X2 U700 ( .A(A[23]), .ZN(n304) );
  NAND2_X2 U701 ( .A1(A[23]), .A2(B[23]), .ZN(net60794) );
  NAND2_X2 U702 ( .A1(n303), .A2(n304), .ZN(net60770) );
  NOR2_X2 U703 ( .A1(A[22]), .A2(B[22]), .ZN(net60767) );
  NOR2_X2 U704 ( .A1(A[22]), .A2(B[22]), .ZN(net60803) );
  NOR2_X2 U705 ( .A1(A[22]), .A2(B[22]), .ZN(net60804) );
  XNOR2_X2 U706 ( .A(A[22]), .B(B[22]), .ZN(net60649) );
  NAND2_X2 U707 ( .A1(net60808), .A2(net60809), .ZN(net60800) );
  INV_X2 U708 ( .A(net60794), .ZN(net60813) );
  NAND2_X2 U709 ( .A1(A[23]), .A2(B[23]), .ZN(net60771) );
  INV_X2 U710 ( .A(net60821), .ZN(net56052) );
  INV_X1 U711 ( .A(net56148), .ZN(net60823) );
  INV_X2 U712 ( .A(net60647), .ZN(net56437) );
  INV_X2 U713 ( .A(net60649), .ZN(net56056) );
  BUF_X1 U714 ( .A(net60758), .Z(net56470) );
  INV_X1 U715 ( .A(net58351), .ZN(net58404) );
  INV_X2 U716 ( .A(net59517), .ZN(net56433) );
  INV_X2 U717 ( .A(net59519), .ZN(net56154) );
  AND2_X1 U718 ( .A1(net58447), .A2(net58242), .ZN(n305) );
  BUF_X1 U719 ( .A(net58329), .Z(net58441) );
  INV_X2 U720 ( .A(A[50]), .ZN(net58422) );
  INV_X2 U721 ( .A(net58243), .ZN(net58389) );
  NAND2_X2 U722 ( .A1(net58422), .A2(net58405), .ZN(net58399) );
  INV_X1 U723 ( .A(net58441), .ZN(net58323) );
  BUF_X1 U724 ( .A(\carry[56] ), .Z(n306) );
  NAND2_X1 U725 ( .A1(n171), .A2(A[55]), .ZN(n307) );
  NAND2_X1 U726 ( .A1(n171), .A2(A[55]), .ZN(n381) );
  NAND2_X1 U727 ( .A1(net62218), .A2(n305), .ZN(net58282) );
  INV_X4 U728 ( .A(net58282), .ZN(net58037) );
  NAND2_X1 U729 ( .A1(A[50]), .A2(net58351), .ZN(net58228) );
  AND2_X2 U730 ( .A1(A[50]), .A2(net58054), .ZN(net58210) );
  INV_X2 U731 ( .A(net58228), .ZN(net58125) );
  XNOR2_X2 U732 ( .A(A[48]), .B(B[48]), .ZN(n308) );
  INV_X2 U733 ( .A(n308), .ZN(net56150) );
  INV_X2 U734 ( .A(net58236), .ZN(net56040) );
  INV_X2 U735 ( .A(net58238), .ZN(net56036) );
  NAND2_X1 U736 ( .A1(A[48]), .A2(B[48]), .ZN(net58226) );
  OR2_X1 U737 ( .A1(net58222), .A2(net58243), .ZN(net58244) );
  INV_X1 U738 ( .A(net58210), .ZN(net58243) );
  NAND2_X1 U739 ( .A1(net58121), .A2(A[52]), .ZN(n309) );
  INV_X2 U740 ( .A(B[51]), .ZN(n310) );
  INV_X2 U741 ( .A(A[51]), .ZN(n311) );
  NAND2_X2 U742 ( .A1(n311), .A2(n310), .ZN(net58054) );
  NAND2_X2 U743 ( .A1(A[51]), .A2(B[51]), .ZN(net58056) );
  XNOR2_X2 U744 ( .A(A[51]), .B(B[51]), .ZN(n312) );
  INV_X2 U745 ( .A(n312), .ZN(net56571) );
  INV_X1 U746 ( .A(net58125), .ZN(net58076) );
  INV_X1 U747 ( .A(net58315), .ZN(net58078) );
  NAND2_X1 U748 ( .A1(net60880), .A2(B[25]), .ZN(n313) );
  NAND2_X1 U749 ( .A1(n302), .A2(B[26]), .ZN(net57097) );
  NAND2_X1 U750 ( .A1(\carry[20] ), .A2(A[20]), .ZN(net57089) );
  BUF_X1 U751 ( .A(n316), .Z(n314) );
  NAND2_X1 U752 ( .A1(net75678), .A2(A[45]), .ZN(n315) );
  NAND2_X1 U753 ( .A1(\carry[45] ), .A2(A[45]), .ZN(net55681) );
  NAND2_X1 U754 ( .A1(n15), .A2(A[59]), .ZN(n357) );
  NAND2_X1 U755 ( .A1(net56431), .A2(A[54]), .ZN(n316) );
  NAND2_X1 U756 ( .A1(net56431), .A2(A[54]), .ZN(n375) );
  BUF_X1 U757 ( .A(net62194), .Z(net57045) );
  BUF_X1 U758 ( .A(n56), .Z(n318) );
  NAND2_X1 U759 ( .A1(n306), .A2(B[56]), .ZN(n319) );
  BUF_X1 U760 ( .A(\carry[46] ), .Z(net57031) );
  NAND2_X1 U761 ( .A1(net57031), .A2(B[46]), .ZN(n320) );
  INV_X1 U762 ( .A(net57085), .ZN(net57024) );
  INV_X1 U763 ( .A(net57024), .ZN(net57025) );
  NAND3_X1 U764 ( .A1(n57), .A2(n381), .A3(n382), .ZN(n321) );
  AND2_X2 U765 ( .A1(B[0]), .A2(A[0]), .ZN(net57022) );
  NAND3_X1 U766 ( .A1(n285), .A2(n296), .A3(n348), .ZN(n322) );
  BUF_X1 U767 ( .A(n322), .Z(n323) );
  NAND3_X1 U768 ( .A1(n259), .A2(n348), .A3(n296), .ZN(\carry[5] ) );
  NAND3_X1 U769 ( .A1(net62177), .A2(n365), .A3(n364), .ZN(net57011) );
  BUF_X1 U770 ( .A(net73524), .Z(net56931) );
  BUF_X1 U771 ( .A(net57080), .Z(net56933) );
  NAND2_X1 U772 ( .A1(n337), .A2(B[20]), .ZN(net56901) );
  NAND3_X1 U773 ( .A1(net62177), .A2(n365), .A3(n364), .ZN(\carry[30] ) );
  NAND2_X1 U774 ( .A1(net57069), .A2(B[45]), .ZN(n324) );
  XOR2_X1 U775 ( .A(net57100), .B(net56887), .Z(SUM[18]) );
  NAND3_X1 U776 ( .A1(net58292), .A2(n309), .A3(net56140), .ZN(n325) );
  NAND2_X1 U777 ( .A1(n341), .A2(B[59]), .ZN(n326) );
  NAND2_X1 U778 ( .A1(n341), .A2(B[59]), .ZN(n358) );
  NAND3_X1 U779 ( .A1(n358), .A2(n357), .A3(n356), .ZN(n327) );
  NAND3_X1 U780 ( .A1(net69188), .A2(net55836), .A3(net55837), .ZN(\carry[15] ) );
  NAND2_X1 U781 ( .A1(\carry[58] ), .A2(A[58]), .ZN(n328) );
  NAND2_X1 U782 ( .A1(\carry[58] ), .A2(A[58]), .ZN(n353) );
  XOR2_X1 U783 ( .A(A[5]), .B(B[5]), .Z(n329) );
  XOR2_X1 U784 ( .A(n329), .B(n323), .Z(SUM[5]) );
  NAND2_X1 U785 ( .A1(A[5]), .A2(B[5]), .ZN(n330) );
  NAND2_X1 U786 ( .A1(\carry[5] ), .A2(A[5]), .ZN(n331) );
  NAND2_X1 U787 ( .A1(n322), .A2(B[5]), .ZN(n332) );
  XOR2_X1 U788 ( .A(net56753), .B(n261), .Z(SUM[6]) );
  NAND2_X1 U789 ( .A1(n258), .A2(A[6]), .ZN(net56755) );
  NAND3_X1 U790 ( .A1(n249), .A2(net55682), .A3(n324), .ZN(n334) );
  NAND3_X1 U791 ( .A1(n315), .A2(net55682), .A3(net56880), .ZN(n333) );
  XOR2_X1 U792 ( .A(B[38]), .B(A[38]), .Z(n335) );
  XOR2_X1 U793 ( .A(net64059), .B(n335), .Z(SUM[38]) );
  NAND2_X1 U794 ( .A1(B[38]), .A2(A[38]), .ZN(net56739) );
  BUF_X1 U795 ( .A(n389), .Z(n336) );
  XOR2_X1 U796 ( .A(net79866), .B(net56639), .Z(SUM[39]) );
  NAND2_X1 U797 ( .A1(net56651), .A2(net56650), .ZN(SUM[63]) );
  INV_X1 U798 ( .A(net56540), .ZN(net56649) );
  INV_X1 U799 ( .A(net55816), .ZN(net56540) );
  BUF_X1 U800 ( .A(n337), .Z(n338) );
  NAND3_X1 U801 ( .A1(n369), .A2(net57091), .A3(n368), .ZN(\carry[20] ) );
  INV_X32 U802 ( .A(net56477), .ZN(net56598) );
  XOR2_X1 U803 ( .A(net56744), .B(net56562), .Z(SUM[40]) );
  XOR2_X1 U804 ( .A(net57006), .B(net56571), .Z(SUM[51]) );
  NAND2_X1 U805 ( .A1(net77806), .A2(net57059), .ZN(net56561) );
  NAND3_X1 U806 ( .A1(net56931), .A2(n376), .A3(n314), .ZN(n339) );
  NAND3_X1 U807 ( .A1(net73524), .A2(n376), .A3(n316), .ZN(n373) );
  NAND2_X1 U808 ( .A1(\carry[48] ), .A2(A[48]), .ZN(net56152) );
  BUF_X1 U809 ( .A(n326), .Z(n340) );
  BUF_X1 U810 ( .A(net62212), .Z(net56467) );
  NAND3_X1 U811 ( .A1(net56549), .A2(n328), .A3(n354), .ZN(n341) );
  XOR2_X1 U812 ( .A(net56468), .B(net56433), .Z(SUM[30]) );
  XOR2_X1 U813 ( .A(net56471), .B(net56437), .Z(SUM[23]) );
  BUF_X1 U814 ( .A(n328), .Z(n342) );
  BUF_X1 U815 ( .A(net56549), .Z(net56363) );
  XOR2_X1 U816 ( .A(net79893), .B(net56368), .Z(SUM[41]) );
  XOR2_X1 U817 ( .A(net56332), .B(net56427), .Z(SUM[42]) );
  XOR2_X1 U818 ( .A(net56336), .B(net56933), .Z(SUM[43]) );
  XOR2_X1 U819 ( .A(net56309), .B(net73634), .Z(SUM[7]) );
  XOR2_X1 U820 ( .A(net56313), .B(net56366), .Z(SUM[8]) );
  BUF_X1 U821 ( .A(n254), .Z(n344) );
  NAND3_X1 U822 ( .A1(net69168), .A2(n239), .A3(n346), .ZN(\carry[4] ) );
  XOR2_X1 U823 ( .A(A[3]), .B(B[3]), .Z(n345) );
  XOR2_X1 U824 ( .A(n345), .B(net56405), .Z(SUM[3]) );
  NAND2_X1 U825 ( .A1(A[3]), .A2(B[3]), .ZN(n346) );
  XOR2_X1 U826 ( .A(A[4]), .B(B[4]), .Z(n347) );
  XOR2_X1 U827 ( .A(n347), .B(n344), .Z(SUM[4]) );
  NAND2_X1 U828 ( .A1(A[4]), .A2(B[4]), .ZN(n348) );
  NAND3_X1 U829 ( .A1(net56363), .A2(n354), .A3(n342), .ZN(n349) );
  NAND3_X1 U830 ( .A1(n13), .A2(n340), .A3(n356), .ZN(n350) );
  BUF_X1 U831 ( .A(B[0]), .Z(n351) );
  XOR2_X1 U832 ( .A(B[58]), .B(A[58]), .Z(n352) );
  XOR2_X1 U833 ( .A(net56400), .B(n352), .Z(SUM[58]) );
  NAND2_X1 U834 ( .A1(B[58]), .A2(A[58]), .ZN(n354) );
  NAND3_X1 U835 ( .A1(n326), .A2(n357), .A3(n356), .ZN(\carry[60] ) );
  XOR2_X1 U836 ( .A(A[59]), .B(B[59]), .Z(n355) );
  XOR2_X1 U837 ( .A(n355), .B(n349), .Z(SUM[59]) );
  NAND2_X1 U838 ( .A1(A[59]), .A2(B[59]), .ZN(n356) );
  XOR2_X1 U839 ( .A(A[60]), .B(B[60]), .Z(n359) );
  NAND2_X1 U840 ( .A1(A[60]), .A2(B[60]), .ZN(net56225) );
  NAND2_X1 U841 ( .A1(\carry[60] ), .A2(A[60]), .ZN(net56226) );
  NAND2_X1 U842 ( .A1(n327), .A2(B[60]), .ZN(net56227) );
  BUF_X1 U843 ( .A(A[0]), .Z(n360) );
  XOR2_X1 U844 ( .A(A[52]), .B(B[52]), .Z(n361) );
  XOR2_X1 U845 ( .A(net58121), .B(n361), .Z(SUM[52]) );
  NAND2_X1 U846 ( .A1(A[52]), .A2(B[52]), .ZN(net56140) );
  XOR2_X1 U847 ( .A(A[53]), .B(B[53]), .Z(n362) );
  XOR2_X1 U848 ( .A(n325), .B(n362), .Z(SUM[53]) );
  XOR2_X1 U849 ( .A(net56883), .B(net56150), .Z(SUM[48]) );
  XOR2_X1 U850 ( .A(net56628), .B(net56154), .Z(SUM[31]) );
  XOR2_X1 U851 ( .A(net58323), .B(net56036), .Z(SUM[49]) );
  XOR2_X1 U852 ( .A(net56040), .B(net58351), .Z(SUM[50]) );
  XOR2_X1 U853 ( .A(net56044), .B(net56210), .Z(SUM[32]) );
  XOR2_X1 U854 ( .A(net56048), .B(n252), .Z(SUM[33]) );
  XOR2_X1 U855 ( .A(net56052), .B(net56428), .Z(SUM[21]) );
  XOR2_X1 U856 ( .A(net56056), .B(net60835), .Z(SUM[22]) );
  XOR2_X1 U857 ( .A(net56060), .B(net56467), .Z(SUM[28]) );
  XOR2_X1 U858 ( .A(A[29]), .B(B[29]), .Z(n363) );
  XOR2_X1 U859 ( .A(n363), .B(net56209), .Z(SUM[29]) );
  NAND2_X1 U860 ( .A1(A[29]), .A2(B[29]), .ZN(n364) );
  NAND2_X1 U861 ( .A1(\carry[29] ), .A2(A[29]), .ZN(n365) );
  BUF_X1 U862 ( .A(net77826), .Z(net56069) );
  NAND2_X1 U863 ( .A1(n339), .A2(B[55]), .ZN(n366) );
  XOR2_X1 U864 ( .A(n256), .B(net56022), .Z(SUM[9]) );
  XOR2_X1 U865 ( .A(A[19]), .B(B[19]), .Z(n367) );
  XOR2_X1 U866 ( .A(n367), .B(net57025), .Z(SUM[19]) );
  NAND2_X1 U867 ( .A1(A[19]), .A2(B[19]), .ZN(n368) );
  NAND2_X1 U868 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n369) );
  XOR2_X1 U869 ( .A(A[20]), .B(B[20]), .Z(n370) );
  XOR2_X1 U870 ( .A(n370), .B(n338), .Z(SUM[20]) );
  NAND2_X1 U871 ( .A1(A[20]), .A2(B[20]), .ZN(net55964) );
  NAND2_X1 U872 ( .A1(\carry[20] ), .A2(A[20]), .ZN(net55965) );
  NAND2_X1 U873 ( .A1(n337), .A2(B[20]), .ZN(net55966) );
  XOR2_X1 U874 ( .A(net55967), .B(net56069), .Z(SUM[10]) );
  BUF_X1 U875 ( .A(n302), .Z(n371) );
  XOR2_X1 U876 ( .A(net55923), .B(net56481), .Z(SUM[12]) );
  XOR2_X1 U877 ( .A(net55927), .B(net56020), .Z(SUM[13]) );
  NAND3_X1 U878 ( .A1(n287), .A2(n382), .A3(n366), .ZN(n372) );
  BUF_X1 U879 ( .A(net60880), .Z(net55936) );
  NAND3_X1 U880 ( .A1(n57), .A2(n307), .A3(n382), .ZN(\carry[56] ) );
  XOR2_X1 U881 ( .A(net55808), .B(net57059), .Z(SUM[1]) );
  XOR2_X1 U882 ( .A(net55812), .B(net56545), .Z(SUM[2]) );
  XOR2_X1 U883 ( .A(B[63]), .B(A[63]), .Z(net55816) );
  XOR2_X1 U884 ( .A(B[54]), .B(A[54]), .Z(n374) );
  XOR2_X1 U885 ( .A(net57004), .B(n374), .Z(SUM[54]) );
  NAND2_X1 U886 ( .A1(B[54]), .A2(A[54]), .ZN(n376) );
  XOR2_X1 U887 ( .A(net56476), .B(net55822), .Z(SUM[44]) );
  XOR2_X1 U888 ( .A(net56158), .B(net55826), .Z(SUM[34]) );
  XOR2_X1 U889 ( .A(net56470), .B(net55830), .Z(SUM[24]) );
  XOR2_X1 U890 ( .A(B[14]), .B(A[14]), .Z(n377) );
  XOR2_X1 U891 ( .A(net56808), .B(n377), .Z(SUM[14]) );
  NAND2_X1 U892 ( .A1(B[14]), .A2(A[14]), .ZN(net55837) );
  NAND3_X1 U893 ( .A1(n336), .A2(n388), .A3(n319), .ZN(n378) );
  NAND3_X1 U894 ( .A1(n318), .A2(n320), .A3(n392), .ZN(n379) );
  XOR2_X1 U895 ( .A(B[55]), .B(A[55]), .Z(n380) );
  XOR2_X1 U896 ( .A(n339), .B(n380), .Z(SUM[55]) );
  NAND2_X1 U897 ( .A1(B[55]), .A2(A[55]), .ZN(n382) );
  XOR2_X1 U898 ( .A(B[45]), .B(A[45]), .Z(n383) );
  XOR2_X1 U899 ( .A(net57069), .B(n383), .Z(SUM[45]) );
  NAND2_X1 U900 ( .A1(B[45]), .A2(A[45]), .ZN(net55682) );
  XOR2_X1 U901 ( .A(net62200), .B(net55683), .Z(SUM[35]) );
  XOR2_X1 U902 ( .A(B[25]), .B(A[25]), .Z(n384) );
  XOR2_X1 U903 ( .A(net55936), .B(n384), .Z(SUM[25]) );
  NAND2_X1 U904 ( .A1(net82511), .A2(B[25]), .ZN(n385) );
  NAND2_X1 U905 ( .A1(B[25]), .A2(A[25]), .ZN(n386) );
  XOR2_X1 U906 ( .A(net67457), .B(net55691), .Z(SUM[15]) );
  NAND3_X1 U907 ( .A1(n390), .A2(n389), .A3(n388), .ZN(\carry[57] ) );
  NAND3_X1 U908 ( .A1(n394), .A2(n393), .A3(n392), .ZN(\carry[47] ) );
  AND2_X2 U909 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
  XOR2_X1 U910 ( .A(A[56]), .B(B[56]), .Z(n387) );
  XOR2_X1 U911 ( .A(n387), .B(n372), .Z(SUM[56]) );
  NAND2_X1 U912 ( .A1(A[56]), .A2(B[56]), .ZN(n388) );
  NAND2_X1 U913 ( .A1(\carry[56] ), .A2(B[56]), .ZN(n390) );
  XOR2_X1 U914 ( .A(net55571), .B(n378), .Z(SUM[57]) );
  XOR2_X1 U915 ( .A(A[46]), .B(B[46]), .Z(n391) );
  XOR2_X1 U916 ( .A(n334), .B(n391), .Z(SUM[46]) );
  NAND2_X1 U917 ( .A1(A[46]), .A2(B[46]), .ZN(n392) );
  NAND2_X1 U918 ( .A1(\carry[46] ), .A2(B[46]), .ZN(n394) );
  XOR2_X1 U919 ( .A(net55579), .B(n379), .Z(SUM[47]) );
  XOR2_X1 U920 ( .A(net55583), .B(net55817), .Z(SUM[36]) );
  XOR2_X1 U921 ( .A(net55587), .B(net55672), .Z(SUM[37]) );
  XOR2_X1 U922 ( .A(A[26]), .B(B[26]), .Z(n395) );
  XOR2_X1 U923 ( .A(n395), .B(n371), .Z(SUM[26]) );
  NAND2_X1 U924 ( .A1(A[26]), .A2(B[26]), .ZN(net55592) );
  XOR2_X1 U925 ( .A(net55595), .B(net55673), .Z(SUM[27]) );
  XOR2_X1 U926 ( .A(net55599), .B(net55976), .Z(SUM[16]) );
  XOR2_X1 U927 ( .A(net55603), .B(net55674), .Z(SUM[17]) );
  XOR2_X1 U928 ( .A(n351), .B(n360), .Z(SUM[0]) );
endmodule


module up_island ( CLK, reset, BUS_NREADY, BUS_BUSY, BUS_MR, BUS_MW, 
        BUS_ADDR_OUTBUS, BUS_DATA_INBUS, BUS_DATA_OUTBUS );
  output [31:0] BUS_ADDR_OUTBUS;
  input [31:0] BUS_DATA_INBUS;
  output [31:0] BUS_DATA_OUTBUS;
  input CLK, reset, BUS_NREADY;
  output BUS_BUSY, BUS_MR, BUS_MW;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, I_BUSY,
         dmem_read, dmem_write, dmem_isbyte, dmem_ishalf, dram_mr, dram_mw,
         iram_rd, N19, N20, N21, N22, N24, N25, N26, N27, N29, N30, N31, N33,
         N34, N35, N37, N38, N40, N41, N42, N43, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, \UUT/N77 ,
         \UUT/N76 , \UUT/m_mem_command[SIGN] , \UUT/m_mem_command[MR] ,
         \UUT/m_we , \UUT/x_we , \UUT/Alu_command[OP][0] ,
         \UUT/Alu_command[OP][1] , \UUT/Alu_command[OP][2] ,
         \UUT/Alu_command[OP][3] , \UUT/Alu_command[OP][4] ,
         \UUT/Alu_command[OP][5] , \UUT/byp_controlB[0] ,
         \UUT/byp_controlB[2] , \UUT/byp_controlA[0] , \UUT/byp_controlA[2] ,
         \UUT/break_code[0] , \UUT/break_code[1] , \UUT/break_code[2] ,
         \UUT/break_code[3] , \UUT/break_code[4] , \UUT/break_code[5] ,
         \UUT/break_code[6] , \UUT/break_code[7] , \UUT/break_code[8] ,
         \UUT/break_code[9] , \UUT/break_code[10] , \UUT/break_code[11] ,
         \UUT/break_code[12] , \UUT/break_code[13] , \UUT/break_code[14] ,
         \UUT/break_code[15] , \UUT/break_code[16] , \UUT/break_code[17] ,
         \UUT/break_code[18] , \UUT/break_code[19] , \UUT/break_code[20] ,
         \UUT/break_code[21] , \UUT/break_code[22] , \UUT/break_code[23] ,
         \UUT/N3 , \UUT/regfile/N457 , \UUT/regfile/N456 , \UUT/regfile/N455 ,
         \UUT/regfile/N451 , \UUT/regfile/N450 , \UUT/regfile/N445 ,
         \UUT/regfile/N444 , \UUT/regfile/N439 , \UUT/regfile/N438 ,
         \UUT/regfile/N433 , \UUT/regfile/N432 , \UUT/regfile/N427 ,
         \UUT/regfile/N426 , \UUT/regfile/N421 , \UUT/regfile/N420 ,
         \UUT/regfile/N415 , \UUT/regfile/N414 , \UUT/regfile/N409 ,
         \UUT/regfile/N408 , \UUT/regfile/N403 , \UUT/regfile/N402 ,
         \UUT/regfile/N397 , \UUT/regfile/N396 , \UUT/regfile/N391 ,
         \UUT/regfile/N390 , \UUT/regfile/N385 , \UUT/regfile/N384 ,
         \UUT/regfile/N379 , \UUT/regfile/N378 , \UUT/regfile/N373 ,
         \UUT/regfile/N372 , \UUT/regfile/N367 , \UUT/regfile/N366 ,
         \UUT/regfile/N360 , \UUT/regfile/N359 , \UUT/regfile/N358 ,
         \UUT/regfile/N354 , \UUT/regfile/N353 , \UUT/regfile/N348 ,
         \UUT/regfile/N347 , \UUT/regfile/N342 , \UUT/regfile/N341 ,
         \UUT/regfile/N336 , \UUT/regfile/N335 , \UUT/regfile/N330 ,
         \UUT/regfile/N329 , \UUT/regfile/N324 , \UUT/regfile/N323 ,
         \UUT/regfile/N318 , \UUT/regfile/N317 , \UUT/regfile/N315 ,
         \UUT/regfile/N311 , \UUT/regfile/N310 , \UUT/regfile/N305 ,
         \UUT/regfile/N304 , \UUT/regfile/N299 , \UUT/regfile/N298 ,
         \UUT/regfile/N293 , \UUT/regfile/N292 , \UUT/regfile/N290 ,
         \UUT/regfile/N286 , \UUT/regfile/N285 , \UUT/regfile/N280 ,
         \UUT/regfile/N279 , \UUT/regfile/N273 , \UUT/regfile/N272 ,
         \UUT/regfile/N269 , \UUT/regfile/N267 , \UUT/regfile/N266 ,
         \UUT/regfile/N265 , \UUT/regfile/N262 , \UUT/regfile/N261 ,
         \UUT/regfile/N260 , \UUT/regfile/reg_out[18][0] ,
         \UUT/regfile/reg_out[18][1] , \UUT/regfile/reg_out[18][2] ,
         \UUT/regfile/reg_out[18][3] , \UUT/regfile/reg_out[18][4] ,
         \UUT/regfile/reg_out[18][5] , \UUT/regfile/reg_out[18][6] ,
         \UUT/regfile/reg_out[18][7] , \UUT/regfile/reg_out[18][8] ,
         \UUT/regfile/reg_out[18][9] , \UUT/regfile/reg_out[18][10] ,
         \UUT/regfile/reg_out[18][11] , \UUT/regfile/reg_out[18][12] ,
         \UUT/regfile/reg_out[18][13] , \UUT/regfile/reg_out[18][14] ,
         \UUT/regfile/reg_out[18][15] , \UUT/regfile/reg_out[18][16] ,
         \UUT/regfile/reg_out[18][17] , \UUT/regfile/reg_out[18][18] ,
         \UUT/regfile/reg_out[18][19] , \UUT/regfile/reg_out[18][20] ,
         \UUT/regfile/reg_out[18][21] , \UUT/regfile/reg_out[18][22] ,
         \UUT/regfile/reg_out[18][23] , \UUT/regfile/reg_out[18][24] ,
         \UUT/regfile/reg_out[18][25] , \UUT/regfile/reg_out[18][26] ,
         \UUT/regfile/reg_out[18][27] , \UUT/regfile/reg_out[18][28] ,
         \UUT/regfile/reg_out[18][29] , \UUT/regfile/reg_out[18][30] ,
         \UUT/regfile/reg_out[18][31] , \UUT/regfile/reg_out[19][0] ,
         \UUT/regfile/reg_out[19][1] , \UUT/regfile/reg_out[19][2] ,
         \UUT/regfile/reg_out[19][3] , \UUT/regfile/reg_out[19][4] ,
         \UUT/regfile/reg_out[19][5] , \UUT/regfile/reg_out[19][6] ,
         \UUT/regfile/reg_out[19][7] , \UUT/regfile/reg_out[19][8] ,
         \UUT/regfile/reg_out[19][9] , \UUT/regfile/reg_out[19][10] ,
         \UUT/regfile/reg_out[19][11] , \UUT/regfile/reg_out[19][12] ,
         \UUT/regfile/reg_out[19][13] , \UUT/regfile/reg_out[19][14] ,
         \UUT/regfile/reg_out[19][15] , \UUT/regfile/reg_out[19][16] ,
         \UUT/regfile/reg_out[19][17] , \UUT/regfile/reg_out[19][18] ,
         \UUT/regfile/reg_out[19][19] , \UUT/regfile/reg_out[19][20] ,
         \UUT/regfile/reg_out[19][21] , \UUT/regfile/reg_out[19][22] ,
         \UUT/regfile/reg_out[19][23] , \UUT/regfile/reg_out[19][24] ,
         \UUT/regfile/reg_out[19][25] , \UUT/regfile/reg_out[19][26] ,
         \UUT/regfile/reg_out[19][27] , \UUT/regfile/reg_out[19][28] ,
         \UUT/regfile/reg_out[19][29] , \UUT/regfile/reg_out[19][30] ,
         \UUT/regfile/reg_out[19][31] , \UUT/regfile/reg_out[20][0] ,
         \UUT/regfile/reg_out[20][1] , \UUT/regfile/reg_out[20][2] ,
         \UUT/regfile/reg_out[20][3] , \UUT/regfile/reg_out[20][4] ,
         \UUT/regfile/reg_out[20][5] , \UUT/regfile/reg_out[20][6] ,
         \UUT/regfile/reg_out[20][7] , \UUT/regfile/reg_out[20][8] ,
         \UUT/regfile/reg_out[20][9] , \UUT/regfile/reg_out[20][10] ,
         \UUT/regfile/reg_out[20][11] , \UUT/regfile/reg_out[20][12] ,
         \UUT/regfile/reg_out[20][13] , \UUT/regfile/reg_out[20][14] ,
         \UUT/regfile/reg_out[20][15] , \UUT/regfile/reg_out[20][16] ,
         \UUT/regfile/reg_out[20][17] , \UUT/regfile/reg_out[20][18] ,
         \UUT/regfile/reg_out[20][19] , \UUT/regfile/reg_out[20][20] ,
         \UUT/regfile/reg_out[20][21] , \UUT/regfile/reg_out[20][22] ,
         \UUT/regfile/reg_out[20][23] , \UUT/regfile/reg_out[20][24] ,
         \UUT/regfile/reg_out[20][25] , \UUT/regfile/reg_out[20][26] ,
         \UUT/regfile/reg_out[20][27] , \UUT/regfile/reg_out[20][28] ,
         \UUT/regfile/reg_out[20][29] , \UUT/regfile/reg_out[20][30] ,
         \UUT/regfile/reg_out[20][31] , \UUT/regfile/reg_out[21][0] ,
         \UUT/regfile/reg_out[21][1] , \UUT/regfile/reg_out[21][2] ,
         \UUT/regfile/reg_out[21][3] , \UUT/regfile/reg_out[21][4] ,
         \UUT/regfile/reg_out[21][5] , \UUT/regfile/reg_out[21][6] ,
         \UUT/regfile/reg_out[21][7] , \UUT/regfile/reg_out[21][8] ,
         \UUT/regfile/reg_out[21][9] , \UUT/regfile/reg_out[21][10] ,
         \UUT/regfile/reg_out[21][11] , \UUT/regfile/reg_out[21][12] ,
         \UUT/regfile/reg_out[21][13] , \UUT/regfile/reg_out[21][14] ,
         \UUT/regfile/reg_out[21][15] , \UUT/regfile/reg_out[21][16] ,
         \UUT/regfile/reg_out[21][17] , \UUT/regfile/reg_out[21][18] ,
         \UUT/regfile/reg_out[21][19] , \UUT/regfile/reg_out[21][20] ,
         \UUT/regfile/reg_out[21][21] , \UUT/regfile/reg_out[21][22] ,
         \UUT/regfile/reg_out[21][23] , \UUT/regfile/reg_out[21][24] ,
         \UUT/regfile/reg_out[21][25] , \UUT/regfile/reg_out[21][26] ,
         \UUT/regfile/reg_out[21][27] , \UUT/regfile/reg_out[21][28] ,
         \UUT/regfile/reg_out[21][29] , \UUT/regfile/reg_out[21][30] ,
         \UUT/regfile/reg_out[21][31] , \UUT/regfile/reg_out[24][0] ,
         \UUT/regfile/reg_out[24][1] , \UUT/regfile/reg_out[24][2] ,
         \UUT/regfile/reg_out[24][3] , \UUT/regfile/reg_out[24][4] ,
         \UUT/regfile/reg_out[24][5] , \UUT/regfile/reg_out[24][6] ,
         \UUT/regfile/reg_out[24][7] , \UUT/regfile/reg_out[24][8] ,
         \UUT/regfile/reg_out[24][9] , \UUT/regfile/reg_out[24][10] ,
         \UUT/regfile/reg_out[24][11] , \UUT/regfile/reg_out[24][12] ,
         \UUT/regfile/reg_out[24][13] , \UUT/regfile/reg_out[24][14] ,
         \UUT/regfile/reg_out[24][15] , \UUT/regfile/reg_out[24][16] ,
         \UUT/regfile/reg_out[24][17] , \UUT/regfile/reg_out[24][18] ,
         \UUT/regfile/reg_out[24][19] , \UUT/regfile/reg_out[24][20] ,
         \UUT/regfile/reg_out[24][21] , \UUT/regfile/reg_out[24][22] ,
         \UUT/regfile/reg_out[24][23] , \UUT/regfile/reg_out[24][24] ,
         \UUT/regfile/reg_out[24][25] , \UUT/regfile/reg_out[24][26] ,
         \UUT/regfile/reg_out[24][27] , \UUT/regfile/reg_out[24][28] ,
         \UUT/regfile/reg_out[24][29] , \UUT/regfile/reg_out[24][30] ,
         \UUT/regfile/reg_out[24][31] , \UUT/regfile/reg_out[25][0] ,
         \UUT/regfile/reg_out[25][1] , \UUT/regfile/reg_out[25][2] ,
         \UUT/regfile/reg_out[25][3] , \UUT/regfile/reg_out[25][4] ,
         \UUT/regfile/reg_out[25][5] , \UUT/regfile/reg_out[25][6] ,
         \UUT/regfile/reg_out[25][7] , \UUT/regfile/reg_out[25][8] ,
         \UUT/regfile/reg_out[25][9] , \UUT/regfile/reg_out[25][10] ,
         \UUT/regfile/reg_out[25][11] , \UUT/regfile/reg_out[25][12] ,
         \UUT/regfile/reg_out[25][13] , \UUT/regfile/reg_out[25][14] ,
         \UUT/regfile/reg_out[25][15] , \UUT/regfile/reg_out[25][16] ,
         \UUT/regfile/reg_out[25][17] , \UUT/regfile/reg_out[25][18] ,
         \UUT/regfile/reg_out[25][19] , \UUT/regfile/reg_out[25][20] ,
         \UUT/regfile/reg_out[25][21] , \UUT/regfile/reg_out[25][22] ,
         \UUT/regfile/reg_out[25][23] , \UUT/regfile/reg_out[25][24] ,
         \UUT/regfile/reg_out[25][25] , \UUT/regfile/reg_out[25][26] ,
         \UUT/regfile/reg_out[25][27] , \UUT/regfile/reg_out[25][28] ,
         \UUT/regfile/reg_out[25][29] , \UUT/regfile/reg_out[25][30] ,
         \UUT/regfile/reg_out[25][31] , \UUT/regfile/reg_out[28][0] ,
         \UUT/regfile/reg_out[28][1] , \UUT/regfile/reg_out[28][2] ,
         \UUT/regfile/reg_out[28][3] , \UUT/regfile/reg_out[28][4] ,
         \UUT/regfile/reg_out[28][5] , \UUT/regfile/reg_out[28][6] ,
         \UUT/regfile/reg_out[28][7] , \UUT/regfile/reg_out[28][8] ,
         \UUT/regfile/reg_out[28][9] , \UUT/regfile/reg_out[28][10] ,
         \UUT/regfile/reg_out[28][11] , \UUT/regfile/reg_out[28][12] ,
         \UUT/regfile/reg_out[28][13] , \UUT/regfile/reg_out[28][14] ,
         \UUT/regfile/reg_out[28][15] , \UUT/regfile/reg_out[28][16] ,
         \UUT/regfile/reg_out[28][17] , \UUT/regfile/reg_out[28][18] ,
         \UUT/regfile/reg_out[28][19] , \UUT/regfile/reg_out[28][20] ,
         \UUT/regfile/reg_out[28][21] , \UUT/regfile/reg_out[28][22] ,
         \UUT/regfile/reg_out[28][23] , \UUT/regfile/reg_out[28][24] ,
         \UUT/regfile/reg_out[28][25] , \UUT/regfile/reg_out[28][26] ,
         \UUT/regfile/reg_out[28][27] , \UUT/regfile/reg_out[28][28] ,
         \UUT/regfile/reg_out[28][29] , \UUT/regfile/reg_out[28][30] ,
         \UUT/regfile/reg_out[28][31] , \UUT/regfile/reg_out[29][0] ,
         \UUT/regfile/reg_out[29][1] , \UUT/regfile/reg_out[29][2] ,
         \UUT/regfile/reg_out[29][3] , \UUT/regfile/reg_out[29][4] ,
         \UUT/regfile/reg_out[29][5] , \UUT/regfile/reg_out[29][6] ,
         \UUT/regfile/reg_out[29][7] , \UUT/regfile/reg_out[29][8] ,
         \UUT/regfile/reg_out[29][9] , \UUT/regfile/reg_out[29][10] ,
         \UUT/regfile/reg_out[29][11] , \UUT/regfile/reg_out[29][12] ,
         \UUT/regfile/reg_out[29][13] , \UUT/regfile/reg_out[29][14] ,
         \UUT/regfile/reg_out[29][15] , \UUT/regfile/reg_out[29][16] ,
         \UUT/regfile/reg_out[29][17] , \UUT/regfile/reg_out[29][18] ,
         \UUT/regfile/reg_out[29][19] , \UUT/regfile/reg_out[29][20] ,
         \UUT/regfile/reg_out[29][21] , \UUT/regfile/reg_out[29][22] ,
         \UUT/regfile/reg_out[29][23] , \UUT/regfile/reg_out[29][24] ,
         \UUT/regfile/reg_out[29][25] , \UUT/regfile/reg_out[29][26] ,
         \UUT/regfile/reg_out[29][27] , \UUT/regfile/reg_out[29][28] ,
         \UUT/regfile/reg_out[29][29] , \UUT/regfile/reg_out[29][30] ,
         \UUT/regfile/reg_out[29][31] , \UUT/regfile/reg_out[4][0] ,
         \UUT/regfile/reg_out[4][1] , \UUT/regfile/reg_out[4][2] ,
         \UUT/regfile/reg_out[4][3] , \UUT/regfile/reg_out[4][4] ,
         \UUT/regfile/reg_out[4][5] , \UUT/regfile/reg_out[4][6] ,
         \UUT/regfile/reg_out[4][7] , \UUT/regfile/reg_out[4][8] ,
         \UUT/regfile/reg_out[4][9] , \UUT/regfile/reg_out[4][10] ,
         \UUT/regfile/reg_out[4][11] , \UUT/regfile/reg_out[4][12] ,
         \UUT/regfile/reg_out[4][13] , \UUT/regfile/reg_out[4][14] ,
         \UUT/regfile/reg_out[4][15] , \UUT/regfile/reg_out[4][16] ,
         \UUT/regfile/reg_out[4][17] , \UUT/regfile/reg_out[4][18] ,
         \UUT/regfile/reg_out[4][19] , \UUT/regfile/reg_out[4][20] ,
         \UUT/regfile/reg_out[4][21] , \UUT/regfile/reg_out[4][22] ,
         \UUT/regfile/reg_out[4][23] , \UUT/regfile/reg_out[4][24] ,
         \UUT/regfile/reg_out[4][25] , \UUT/regfile/reg_out[4][26] ,
         \UUT/regfile/reg_out[4][27] , \UUT/regfile/reg_out[4][28] ,
         \UUT/regfile/reg_out[4][29] , \UUT/regfile/reg_out[4][30] ,
         \UUT/regfile/reg_out[4][31] , \UUT/regfile/reg_out[5][0] ,
         \UUT/regfile/reg_out[5][1] , \UUT/regfile/reg_out[5][2] ,
         \UUT/regfile/reg_out[5][3] , \UUT/regfile/reg_out[5][4] ,
         \UUT/regfile/reg_out[5][5] , \UUT/regfile/reg_out[5][6] ,
         \UUT/regfile/reg_out[5][7] , \UUT/regfile/reg_out[5][8] ,
         \UUT/regfile/reg_out[5][9] , \UUT/regfile/reg_out[5][10] ,
         \UUT/regfile/reg_out[5][11] , \UUT/regfile/reg_out[5][12] ,
         \UUT/regfile/reg_out[5][13] , \UUT/regfile/reg_out[5][14] ,
         \UUT/regfile/reg_out[5][15] , \UUT/regfile/reg_out[5][16] ,
         \UUT/regfile/reg_out[5][17] , \UUT/regfile/reg_out[5][18] ,
         \UUT/regfile/reg_out[5][19] , \UUT/regfile/reg_out[5][20] ,
         \UUT/regfile/reg_out[5][21] , \UUT/regfile/reg_out[5][22] ,
         \UUT/regfile/reg_out[5][23] , \UUT/regfile/reg_out[5][24] ,
         \UUT/regfile/reg_out[5][25] , \UUT/regfile/reg_out[5][26] ,
         \UUT/regfile/reg_out[5][27] , \UUT/regfile/reg_out[5][28] ,
         \UUT/regfile/reg_out[5][29] , \UUT/regfile/reg_out[5][30] ,
         \UUT/regfile/reg_out[5][31] , \UUT/BYP_BRANCH_MUXB/N39 ,
         \UUT/BYP_BRANCH_MUXB/N4 , \UUT/Mcontrol/N19 ,
         \UUT/Mcontrol/x_sampled_dmem_command[SIGN] ,
         \UUT/Mcontrol/x_sampled_dmem_command[MW] ,
         \UUT/Mcontrol/x_sampled_dmem_command[MR] ,
         \UUT/Mcontrol/x_sampled_dmem_command[MH] ,
         \UUT/Mcontrol/x_sampled_dmem_command[MB] ,
         \UUT/Mcontrol/m_sampled_xrd[0] , \UUT/Mcontrol/m_sampled_xrd[1] ,
         \UUT/Mcontrol/m_sampled_xrd[2] , \UUT/Mcontrol/m_sampled_xrd[3] ,
         \UUT/Mcontrol/m_sampled_xrd[4] , \UUT/Mcontrol/x_rd[0] ,
         \UUT/Mcontrol/x_rd[1] , \UUT/Mcontrol/x_rd[2] ,
         \UUT/Mcontrol/x_rd[3] , \UUT/Mcontrol/x_rd[4] ,
         \UUT/Mcontrol/d_jump_type[0] , \UUT/Mcontrol/d_jump_type[1] ,
         \UUT/Mcontrol/d_jump_type[2] , \UUT/Mcontrol/d_jump_type[3] ,
         \UUT/Mcontrol/int_reset , \UUT/Mcontrol/Program_counter/N24 ,
         \UUT/Mcontrol/Program_counter/N22 ,
         \UUT/Mcontrol/Program_counter/N20 , \UUT/Mcontrol/Program_counter/N8 ,
         \UUT/Mcontrol/Operation_decoding32/N2089 ,
         \UUT/Mcontrol/Operation_decoding32/N2088 ,
         \UUT/Mcontrol/Operation_decoding32/N2087 ,
         \UUT/Mcontrol/Operation_decoding32/N2086 ,
         \UUT/Mcontrol/Operation_decoding32/N2085 ,
         \UUT/Mcontrol/Operation_decoding32/N2084 ,
         \UUT/Mcontrol/Operation_decoding32/N2083 ,
         \UUT/Mcontrol/Operation_decoding32/N2082 ,
         \UUT/Mcontrol/Operation_decoding32/N2081 ,
         \UUT/Mcontrol/Operation_decoding32/N2080 ,
         \UUT/Mcontrol/Operation_decoding32/N2079 ,
         \UUT/Mcontrol/Operation_decoding32/N2077 ,
         \UUT/Mcontrol/Operation_decoding32/N2076 ,
         \UUT/Mcontrol/Operation_decoding32/N2075 ,
         \UUT/Mcontrol/Operation_decoding32/N2074 ,
         \UUT/Mcontrol/Operation_decoding32/N2071 ,
         \UUT/Mcontrol/Operation_decoding32/N2070 ,
         \UUT/Mcontrol/Operation_decoding32/N2069 ,
         \UUT/Mcontrol/Operation_decoding32/N2068 ,
         \UUT/Mcontrol/Operation_decoding32/N2066 ,
         \UUT/Mcontrol/Operation_decoding32/N2065 ,
         \UUT/Mcontrol/Operation_decoding32/N2064 ,
         \UUT/Mcontrol/Operation_decoding32/N2063 ,
         \UUT/Mcontrol/Operation_decoding32/N2062 ,
         \UUT/Mcontrol/Operation_decoding32/N2061 ,
         \UUT/Mcontrol/Operation_decoding32/N2060 ,
         \UUT/Mcontrol/Operation_decoding32/N2059 ,
         \UUT/Mcontrol/Operation_decoding32/N2058 ,
         \UUT/Mcontrol/Operation_decoding32/N2057 ,
         \UUT/Mcontrol/Operation_decoding32/N2056 ,
         \UUT/Mcontrol/Operation_decoding32/N2054 ,
         \UUT/Mcontrol/Operation_decoding32/N2053 ,
         \UUT/Mcontrol/Operation_decoding32/N2052 ,
         \UUT/Mcontrol/Operation_decoding32/N2051 ,
         \UUT/Mcontrol/Operation_decoding32/N2050 ,
         \UUT/Mcontrol/Operation_decoding32/N2047 ,
         \UUT/Mcontrol/Operation_decoding32/N2046 ,
         \UUT/Mcontrol/Operation_decoding32/N2045 ,
         \UUT/Mcontrol/Operation_decoding32/N2044 ,
         \UUT/Mcontrol/Operation_decoding32/N2043 ,
         \UUT/Mcontrol/Operation_decoding32/N2041 ,
         \UUT/Mcontrol/Operation_decoding32/N2040 ,
         \UUT/Mcontrol/Operation_decoding32/N2039 ,
         \UUT/Mcontrol/Operation_decoding32/N2038 ,
         \UUT/Mcontrol/Operation_decoding32/N2037 ,
         \UUT/Mcontrol/Operation_decoding32/N2036 ,
         \UUT/Mcontrol/Operation_decoding32/N2035 ,
         \UUT/Mcontrol/Operation_decoding32/N2034 ,
         \UUT/Mcontrol/Operation_decoding32/N2033 ,
         \UUT/Mcontrol/Operation_decoding32/N2032 ,
         \UUT/Mcontrol/Operation_decoding32/N2030 ,
         \UUT/Mcontrol/Operation_decoding32/N2029 ,
         \UUT/Mcontrol/Operation_decoding32/N2028 ,
         \UUT/Mcontrol/Operation_decoding32/N2027 ,
         \UUT/Mcontrol/Operation_decoding32/N2026 ,
         \UUT/Mcontrol/Operation_decoding32/N2025 ,
         \UUT/Mcontrol/Operation_decoding32/N2023 ,
         \UUT/Mcontrol/Operation_decoding32/N2022 ,
         \UUT/Mcontrol/Operation_decoding32/N2021 ,
         \UUT/Mcontrol/Operation_decoding32/N2020 ,
         \UUT/Mcontrol/Operation_decoding32/N2019 ,
         \UUT/Mcontrol/Operation_decoding32/N2017 ,
         \UUT/Mcontrol/Operation_decoding32/N2016 ,
         \UUT/Mcontrol/Operation_decoding32/N2015 ,
         \UUT/Mcontrol/Operation_decoding32/N2014 ,
         \UUT/Mcontrol/Operation_decoding32/N2010 ,
         \UUT/Mcontrol/Operation_decoding32/N2009 ,
         \UUT/Mcontrol/Operation_decoding32/N2008 ,
         \UUT/Mcontrol/Operation_decoding32/N2007 ,
         \UUT/Mcontrol/Operation_decoding32/N2005 ,
         \UUT/Mcontrol/Operation_decoding32/N2004 ,
         \UUT/Mcontrol/Operation_decoding32/N2003 ,
         \UUT/Mcontrol/Operation_decoding32/N2002 ,
         \UUT/Mcontrol/Operation_decoding32/N2001 ,
         \UUT/Mcontrol/Operation_decoding32/N1999 ,
         \UUT/Mcontrol/Operation_decoding32/N1998 ,
         \UUT/Mcontrol/Operation_decoding32/N1997 ,
         \UUT/Mcontrol/Operation_decoding32/N1996 ,
         \UUT/Mcontrol/Operation_decoding32/N1995 ,
         \UUT/Mcontrol/Operation_decoding32/N1994 ,
         \UUT/Mcontrol/Operation_decoding32/N1993 ,
         \UUT/Mcontrol/Operation_decoding32/N1992 ,
         \UUT/Mcontrol/Operation_decoding32/N1991 ,
         \UUT/Mcontrol/Operation_decoding32/N1990 ,
         \UUT/Mcontrol/Operation_decoding32/N1989 ,
         \UUT/Mcontrol/Operation_decoding32/N1987 ,
         \UUT/Mcontrol/Operation_decoding32/N1986 ,
         \UUT/Mcontrol/Operation_decoding32/N1985 ,
         \UUT/Mcontrol/Operation_decoding32/N1984 ,
         \UUT/Mcontrol/Operation_decoding32/N1983 ,
         \UUT/Mcontrol/Operation_decoding32/N1981 ,
         \UUT/Mcontrol/Operation_decoding32/N1980 ,
         \UUT/Mcontrol/Operation_decoding32/N1979 ,
         \UUT/Mcontrol/Operation_decoding32/N1978 ,
         \UUT/Mcontrol/Operation_decoding32/N1977 ,
         \UUT/Mcontrol/Operation_decoding32/N1976 ,
         \UUT/Mcontrol/Operation_decoding32/N1975 ,
         \UUT/Mcontrol/Operation_decoding32/N1974 ,
         \UUT/Mcontrol/Operation_decoding32/N1973 ,
         \UUT/Mcontrol/Operation_decoding32/N1972 ,
         \UUT/Mcontrol/Operation_decoding32/N1971 ,
         \UUT/Mcontrol/Operation_decoding32/N1970 ,
         \UUT/Mcontrol/Operation_decoding32/N1969 ,
         \UUT/Mcontrol/Operation_decoding32/N1968 ,
         \UUT/Mcontrol/Operation_decoding32/N1967 ,
         \UUT/Mcontrol/Operation_decoding32/N1966 ,
         \UUT/Mcontrol/Operation_decoding32/N1965 ,
         \UUT/Mcontrol/Operation_decoding32/N1964 ,
         \UUT/Mcontrol/Operation_decoding32/N1963 ,
         \UUT/Mcontrol/Operation_decoding32/N1962 ,
         \UUT/Mcontrol/Operation_decoding32/N1961 ,
         \UUT/Mcontrol/Operation_decoding32/N1960 ,
         \UUT/Mcontrol/Operation_decoding32/N1959 ,
         \UUT/Mcontrol/Operation_decoding32/N1958 ,
         \UUT/Mcontrol/Operation_decoding32/N1957 ,
         \UUT/Mcontrol/Operation_decoding32/N1956 ,
         \UUT/Mcontrol/Operation_decoding32/N1955 ,
         \UUT/Mcontrol/Operation_decoding32/N1954 ,
         \UUT/Mcontrol/Operation_decoding32/N1953 ,
         \UUT/Mcontrol/Operation_decoding32/N1952 ,
         \UUT/Mcontrol/Operation_decoding32/N1951 ,
         \UUT/Mcontrol/Operation_decoding32/N1950 ,
         \UUT/Mcontrol/Operation_decoding32/N1949 ,
         \UUT/Mcontrol/Operation_decoding32/N1948 ,
         \UUT/Mcontrol/Operation_decoding32/N1947 ,
         \UUT/Mcontrol/Operation_decoding32/N1946 ,
         \UUT/Mcontrol/Operation_decoding32/N1945 ,
         \UUT/Mcontrol/Operation_decoding32/N1944 ,
         \UUT/Mcontrol/Operation_decoding32/N1943 ,
         \UUT/Mcontrol/Operation_decoding32/N1942 ,
         \UUT/Mcontrol/Operation_decoding32/N1941 ,
         \UUT/Mcontrol/Operation_decoding32/N1940 ,
         \UUT/Mcontrol/Operation_decoding32/N1939 ,
         \UUT/Mcontrol/Operation_decoding32/N1938 ,
         \UUT/Mcontrol/Operation_decoding32/N1937 ,
         \UUT/Mcontrol/Operation_decoding32/N1936 ,
         \UUT/Mcontrol/Operation_decoding32/N1935 ,
         \UUT/Mcontrol/Operation_decoding32/N1934 ,
         \UUT/Mcontrol/Operation_decoding32/N1933 ,
         \UUT/Mcontrol/Operation_decoding32/N1932 ,
         \UUT/Mcontrol/Operation_decoding32/N1931 ,
         \UUT/Mcontrol/Operation_decoding32/N1930 ,
         \UUT/Mcontrol/Operation_decoding32/N1929 ,
         \UUT/Mcontrol/Operation_decoding32/N1928 ,
         \UUT/Mcontrol/Operation_decoding32/N1927 ,
         \UUT/Mcontrol/Operation_decoding32/N1926 ,
         \UUT/Mcontrol/Operation_decoding32/N1925 ,
         \UUT/Mcontrol/Operation_decoding32/N1924 ,
         \UUT/Mcontrol/Operation_decoding32/N1923 ,
         \UUT/Mcontrol/Operation_decoding32/N1922 ,
         \UUT/Mcontrol/Operation_decoding32/N1921 ,
         \UUT/Mcontrol/Operation_decoding32/N1920 ,
         \UUT/Mcontrol/Operation_decoding32/N1919 ,
         \UUT/Mcontrol/Operation_decoding32/N1918 ,
         \UUT/Mcontrol/Operation_decoding32/N1917 ,
         \UUT/Mcontrol/Operation_decoding32/N1916 ,
         \UUT/Mcontrol/Operation_decoding32/N1915 ,
         \UUT/Mcontrol/Operation_decoding32/N1914 ,
         \UUT/Mcontrol/Operation_decoding32/N1913 ,
         \UUT/Mcontrol/Operation_decoding32/N1912 ,
         \UUT/Mcontrol/Operation_decoding32/N1911 ,
         \UUT/Mcontrol/Operation_decoding32/N1910 ,
         \UUT/Mcontrol/Operation_decoding32/N1909 ,
         \UUT/Mcontrol/Operation_decoding32/N1908 ,
         \UUT/Mcontrol/Operation_decoding32/N1907 ,
         \UUT/Mcontrol/Operation_decoding32/N1906 ,
         \UUT/Mcontrol/Operation_decoding32/N1905 ,
         \UUT/Mcontrol/Operation_decoding32/N1904 ,
         \UUT/Mcontrol/Operation_decoding32/N1903 ,
         \UUT/Mcontrol/Operation_decoding32/N1902 ,
         \UUT/Mcontrol/Operation_decoding32/N1901 ,
         \UUT/Mcontrol/Operation_decoding32/N1900 ,
         \UUT/Mcontrol/Operation_decoding32/N1899 ,
         \UUT/Mcontrol/Operation_decoding32/N1898 ,
         \UUT/Mcontrol/Operation_decoding32/N1897 ,
         \UUT/Mcontrol/Operation_decoding32/N1896 ,
         \UUT/Mcontrol/Operation_decoding32/N1895 ,
         \UUT/Mcontrol/Operation_decoding32/N1894 ,
         \UUT/Mcontrol/Operation_decoding32/N1893 ,
         \UUT/Mcontrol/Operation_decoding32/N1892 ,
         \UUT/Mcontrol/Operation_decoding32/N1891 ,
         \UUT/Mcontrol/Operation_decoding32/N1890 ,
         \UUT/Mcontrol/Operation_decoding32/N1889 ,
         \UUT/Mcontrol/Operation_decoding32/N1888 ,
         \UUT/Mcontrol/Operation_decoding32/N1887 ,
         \UUT/Mcontrol/Operation_decoding32/N1886 ,
         \UUT/Mcontrol/Operation_decoding32/N1885 ,
         \UUT/Mcontrol/Operation_decoding32/N1884 ,
         \UUT/Mcontrol/Operation_decoding32/N1883 ,
         \UUT/Mcontrol/Operation_decoding32/N1882 ,
         \UUT/Mcontrol/Operation_decoding32/N1881 ,
         \UUT/Mcontrol/Operation_decoding32/N1880 ,
         \UUT/Mcontrol/Operation_decoding32/N1879 ,
         \UUT/Mcontrol/Operation_decoding32/N1878 ,
         \UUT/Mcontrol/Operation_decoding32/N1877 ,
         \UUT/Mcontrol/Operation_decoding32/N1876 ,
         \UUT/Mcontrol/Operation_decoding32/N1875 ,
         \UUT/Mcontrol/Operation_decoding32/N1873 ,
         \UUT/Mcontrol/Operation_decoding32/N1871 ,
         \UUT/Mcontrol/Operation_decoding32/N89 ,
         \UUT/Mcontrol/Operation_decoding32/N62 ,
         \UUT/Mcontrol/Nextpc_decoding/N266 ,
         \UUT/Mcontrol/Nextpc_decoding/N265 ,
         \UUT/Mcontrol/Nextpc_decoding/N264 ,
         \UUT/Mcontrol/Nextpc_decoding/N263 ,
         \UUT/Mcontrol/Nextpc_decoding/N262 ,
         \UUT/Mcontrol/Nextpc_decoding/N260 ,
         \UUT/Mcontrol/Nextpc_decoding/N259 ,
         \UUT/Mcontrol/Nextpc_decoding/N258 ,
         \UUT/Mcontrol/Nextpc_decoding/N257 ,
         \UUT/Mcontrol/Nextpc_decoding/N256 ,
         \UUT/Mcontrol/Nextpc_decoding/N255 ,
         \UUT/Mcontrol/Nextpc_decoding/N254 ,
         \UUT/Mcontrol/Nextpc_decoding/N253 ,
         \UUT/Mcontrol/Nextpc_decoding/N252 ,
         \UUT/Mcontrol/Nextpc_decoding/N251 ,
         \UUT/Mcontrol/Nextpc_decoding/N250 ,
         \UUT/Mcontrol/Nextpc_decoding/N248 ,
         \UUT/Mcontrol/Nextpc_decoding/N247 ,
         \UUT/Mcontrol/Nextpc_decoding/N246 ,
         \UUT/Mcontrol/Nextpc_decoding/N245 ,
         \UUT/Mcontrol/Nextpc_decoding/N244 ,
         \UUT/Mcontrol/Nextpc_decoding/N242 ,
         \UUT/Mcontrol/Nextpc_decoding/N241 ,
         \UUT/Mcontrol/Nextpc_decoding/N240 ,
         \UUT/Mcontrol/Nextpc_decoding/N239 ,
         \UUT/Mcontrol/Nextpc_decoding/N238 ,
         \UUT/Mcontrol/Nextpc_decoding/N236 ,
         \UUT/Mcontrol/Nextpc_decoding/N235 ,
         \UUT/Mcontrol/Nextpc_decoding/N234 ,
         \UUT/Mcontrol/Nextpc_decoding/N233 ,
         \UUT/Mcontrol/Nextpc_decoding/N232 ,
         \UUT/Mcontrol/Nextpc_decoding/N230 ,
         \UUT/Mcontrol/Nextpc_decoding/N229 ,
         \UUT/Mcontrol/Nextpc_decoding/N228 ,
         \UUT/Mcontrol/Nextpc_decoding/N227 ,
         \UUT/Mcontrol/Nextpc_decoding/N226 ,
         \UUT/Mcontrol/Nextpc_decoding/N224 ,
         \UUT/Mcontrol/Nextpc_decoding/N223 ,
         \UUT/Mcontrol/Nextpc_decoding/N222 ,
         \UUT/Mcontrol/Nextpc_decoding/N191 ,
         \UUT/Mcontrol/Nextpc_decoding/N160 ,
         \UUT/Mcontrol/Nextpc_decoding/N159 ,
         \UUT/Mcontrol/Nextpc_decoding/N125 ,
         \UUT/Mcontrol/Nextpc_decoding/N124 ,
         \UUT/Mcontrol/Nextpc_decoding/N123 ,
         \UUT/Mcontrol/Nextpc_decoding/N122 ,
         \UUT/Mcontrol/Nextpc_decoding/N120 ,
         \UUT/Mcontrol/Nextpc_decoding/N116 ,
         \UUT/Mcontrol/Nextpc_decoding/N115 ,
         \UUT/Mcontrol/Nextpc_decoding/N114 ,
         \UUT/Mcontrol/Nextpc_decoding/N32 ,
         \UUT/Mcontrol/Nextpc_decoding/N27 ,
         \UUT/Mcontrol/Nextpc_decoding/N25 ,
         \UUT/Mcontrol/Nextpc_decoding/condition ,
         \UUT/Mcontrol/Nextpc_decoding/N22 , \UUT/Mcontrol/bp_logicA/N16 ,
         \UUT/Mcontrol/bp_logicA/N15 , \UUT/Mcontrol/bp_logicA/N14 ,
         \UUT/Mcontrol/bp_logicA/N13 , \UUT/Mcontrol/bp_logicA/N12 ,
         \UUT/Mcontrol/bp_logicA/N11 , \UUT/Mcontrol/bp_logicA/N10 ,
         \UUT/Mcontrol/bp_logicA/N9 , \UUT/Mcontrol/bp_logicA/N8 ,
         \UUT/Mcontrol/bp_logicA/N7 , \UUT/Mcontrol/bp_logicA/N6 ,
         \UUT/Mcontrol/bp_logicA/N5 , \UUT/Mcontrol/bp_logicA/memory_main ,
         \UUT/Mcontrol/bp_logicA/N3 , \UUT/Mcontrol/bp_logicA/exec_main ,
         \UUT/Mcontrol/bp_logicA/N2 , \UUT/Mcontrol/bp_logicB/N16 ,
         \UUT/Mcontrol/bp_logicB/N15 , \UUT/Mcontrol/bp_logicB/N14 ,
         \UUT/Mcontrol/bp_logicB/N13 , \UUT/Mcontrol/bp_logicB/N12 ,
         \UUT/Mcontrol/bp_logicB/N11 , \UUT/Mcontrol/bp_logicB/N10 ,
         \UUT/Mcontrol/bp_logicB/N9 , \UUT/Mcontrol/bp_logicB/N8 ,
         \UUT/Mcontrol/bp_logicB/N7 , \UUT/Mcontrol/bp_logicB/N6 ,
         \UUT/Mcontrol/bp_logicB/N5 , \UUT/Mcontrol/bp_logicB/memory_main ,
         \UUT/Mcontrol/bp_logicB/N3 , \UUT/Mcontrol/bp_logicB/exec_main ,
         \UUT/Mcontrol/bp_logicB/N2 , \UUT/Mcontrol/st_logic/N120 ,
         \UUT/Mcontrol/st_logic/N119 , \UUT/Mcontrol/st_logic/N118 ,
         \UUT/Mcontrol/st_logic/N117 , \UUT/Mcontrol/st_logic/N116 ,
         \UUT/Mcontrol/st_logic/N115 , \UUT/Mcontrol/st_logic/N114 ,
         \UUT/Mcontrol/st_logic/N113 , \UUT/Mcontrol/st_logic/N112 ,
         \UUT/Mcontrol/st_logic/N111 , \UUT/Mcontrol/st_logic/N110 ,
         \UUT/Mcontrol/st_logic/N109 , \UUT/Mcontrol/st_logic/N108 ,
         \UUT/Mcontrol/st_logic/N107 , \UUT/Mcontrol/st_logic/N106 ,
         \UUT/Mcontrol/st_logic/N105 , \UUT/Mcontrol/st_logic/N103 ,
         \UUT/Mcontrol/st_logic/N102 , \UUT/Mcontrol/st_logic/N101 ,
         \UUT/Mcontrol/st_logic/N100 , \UUT/Mcontrol/st_logic/N99 ,
         \UUT/Mcontrol/st_logic/N98 , \UUT/Mcontrol/st_logic/N96 ,
         \UUT/Mcontrol/st_logic/N95 , \UUT/Mcontrol/st_logic/N94 ,
         \UUT/Mcontrol/st_logic/N93 , \UUT/Mcontrol/st_logic/N92 ,
         \UUT/Mcontrol/st_logic/N90 , \UUT/Mcontrol/st_logic/N89 ,
         \UUT/Mcontrol/st_logic/N88 , \UUT/Mcontrol/st_logic/N87 ,
         \UUT/Mcontrol/st_logic/N86 , \UUT/Mcontrol/st_logic/N85 ,
         \UUT/Mcontrol/st_logic/N83 , \UUT/Mcontrol/st_logic/N82 ,
         \UUT/Mcontrol/st_logic/N81 , \UUT/Mcontrol/st_logic/N80 ,
         \UUT/Mcontrol/st_logic/N79 , \UUT/Mcontrol/st_logic/N77 ,
         \UUT/Mcontrol/st_logic/N76 , \UUT/Mcontrol/st_logic/N75 ,
         \UUT/Mcontrol/st_logic/N74 , \UUT/Mcontrol/st_logic/N73 ,
         \UUT/Mcontrol/st_logic/N71 , \UUT/Mcontrol/st_logic/N70 ,
         \UUT/Mcontrol/st_logic/N69 , \UUT/Mcontrol/st_logic/N68 ,
         \UUT/Mcontrol/st_logic/N67 , \UUT/Mcontrol/st_logic/N65 ,
         \UUT/Mcontrol/st_logic/N64 , \UUT/Mcontrol/st_logic/N63 ,
         \UUT/Mcontrol/st_logic/N62 , \UUT/Mcontrol/st_logic/N61 ,
         \UUT/Mcontrol/st_logic/N60 , \UUT/Mcontrol/st_logic/N58 ,
         \UUT/Mcontrol/st_logic/N57 , \UUT/Mcontrol/st_logic/N56 ,
         \UUT/Mcontrol/st_logic/N55 , \UUT/Mcontrol/st_logic/N54 ,
         \UUT/Mcontrol/st_logic/N53 , \UUT/Mcontrol/st_logic/N52 ,
         \UUT/Mcontrol/st_logic/N51 , \UUT/Mcontrol/st_logic/N50 ,
         \UUT/Mcontrol/st_logic/N49 , \UUT/Mcontrol/st_logic/N47 ,
         \UUT/Mcontrol/st_logic/N46 , \UUT/Mcontrol/st_logic/N45 ,
         \UUT/Mcontrol/st_logic/N44 , \UUT/Mcontrol/st_logic/N42 ,
         \UUT/Mcontrol/st_logic/N41 , \UUT/Mcontrol/st_logic/N40 ,
         \UUT/Mcontrol/st_logic/N39 , \UUT/Mcontrol/st_logic/N38 ,
         \UUT/Mcontrol/st_logic/N37 , \UUT/Mcontrol/st_logic/N36 ,
         \UUT/Mcontrol/st_logic/N35 , \UUT/Mcontrol/st_logic/N34 ,
         \UUT/Mcontrol/st_logic/N33 , \UUT/Mcontrol/st_logic/N32 ,
         \UUT/Mcontrol/st_logic/N31 , \UUT/Mcontrol/st_logic/N30 ,
         \UUT/Mcontrol/st_logic/N29 , \UUT/Mcontrol/st_logic/N28 ,
         \UUT/Mcontrol/st_logic/N27 , \UUT/Mcontrol/st_logic/N26 ,
         \UUT/Mcontrol/st_logic/N25 , \UUT/Mcontrol/st_logic/N24 ,
         \UUT/Mcontrol/st_logic/N23 , \UUT/Mcontrol/st_logic/N22 ,
         \UUT/Mcontrol/st_logic/N19 , \UUT/Mcontrol/st_logic/N18 ,
         \UUT/Mcontrol/st_logic/N15 , \UUT/Mcontrol/st_logic/N14 ,
         \UUT/Mcontrol/st_logic/N13 , \UUT/Mcontrol/st_logic/N12 ,
         \UUT/Mcontrol/st_logic/N10 , \UUT/Mcontrol/st_logic/branchmul_stall ,
         \UUT/Mcontrol/st_logic/N8 ,
         \UUT/Mcontrol/st_logic/branch_uses_main_exe_result ,
         \UUT/Mcontrol/st_logic/N7 , \UUT/Mcontrol/st_logic/branchlw_stall ,
         \UUT/Mcontrol/st_logic/N6 ,
         \UUT/Mcontrol/st_logic/branch_uses_main_mem_result ,
         \UUT/Mcontrol/st_logic/N5 , \UUT/Mcontrol/st_logic/branch_uses_regb ,
         \UUT/Mcontrol/st_logic/N4 , \UUT/Mcontrol/st_logic/branch_uses_rega ,
         \UUT/Mcontrol/st_logic/N3 , \UUT/Mcontrol/st_logic/load_stall ,
         \UUT/Mcontrol/st_logic/N2 , \UUT/Mpath/N128 , \UUT/Mpath/N127 ,
         \UUT/Mpath/N125 , \UUT/Mpath/N124 , \UUT/Mpath/N121 ,
         \UUT/Mpath/N119 , \UUT/Mpath/N118 , \UUT/Mpath/N117 ,
         \UUT/Mpath/N116 , \UUT/Mpath/N115 , \UUT/Mpath/N114 ,
         \UUT/Mpath/N113 , \UUT/Mpath/N112 , \UUT/Mpath/N111 ,
         \UUT/Mpath/out_jar[0] , \UUT/Mpath/out_jar[1] ,
         \UUT/Mpath/out_jar[2] , \UUT/Mpath/out_jar[3] ,
         \UUT/Mpath/out_jar[4] , \UUT/Mpath/out_jar[5] ,
         \UUT/Mpath/out_jar[6] , \UUT/Mpath/out_jar[7] ,
         \UUT/Mpath/out_jar[8] , \UUT/Mpath/out_jar[9] ,
         \UUT/Mpath/out_jar[10] , \UUT/Mpath/out_jar[11] ,
         \UUT/Mpath/out_jar[12] , \UUT/Mpath/out_jar[13] ,
         \UUT/Mpath/out_jar[14] , \UUT/Mpath/out_jar[15] ,
         \UUT/Mpath/out_jar[16] , \UUT/Mpath/out_jar[17] ,
         \UUT/Mpath/out_jar[18] , \UUT/Mpath/out_jar[19] ,
         \UUT/Mpath/out_jar[20] , \UUT/Mpath/out_jar[21] ,
         \UUT/Mpath/out_jar[22] , \UUT/Mpath/out_jar[23] ,
         \UUT/Mpath/out_regB[0] , \UUT/Mpath/out_regB[1] ,
         \UUT/Mpath/out_regB[2] , \UUT/Mpath/out_regB[3] ,
         \UUT/Mpath/out_regB[4] , \UUT/Mpath/out_regB[5] ,
         \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[7] ,
         \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[9] ,
         \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[11] ,
         \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[13] ,
         \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[15] ,
         \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[17] ,
         \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[19] ,
         \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[21] ,
         \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[23] ,
         \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[25] ,
         \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[27] ,
         \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[29] ,
         \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[31] ,
         \UUT/Mpath/out_regA[0] , \UUT/Mpath/out_regA[1] ,
         \UUT/Mpath/out_regA[2] , \UUT/Mpath/out_regA[3] ,
         \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[5] ,
         \UUT/Mpath/out_regA[6] , \UUT/Mpath/out_regA[7] ,
         \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[9] ,
         \UUT/Mpath/out_regA[10] , \UUT/Mpath/out_regA[11] ,
         \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[13] ,
         \UUT/Mpath/out_regA[14] , \UUT/Mpath/out_regA[15] ,
         \UUT/Mpath/out_regA[16] , \UUT/Mpath/out_regA[17] ,
         \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[19] ,
         \UUT/Mpath/out_regA[20] , \UUT/Mpath/out_regA[21] ,
         \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[23] ,
         \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[25] ,
         \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[27] ,
         \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[29] ,
         \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[31] ,
         \UUT/Mpath/the_alu/N526 , \UUT/Mpath/the_alu/N525 ,
         \UUT/Mpath/the_alu/N524 , \UUT/Mpath/the_alu/N523 ,
         \UUT/Mpath/the_alu/N520 , \UUT/Mpath/the_alu/N519 ,
         \UUT/Mpath/the_alu/N518 , \UUT/Mpath/the_alu/N517 ,
         \UUT/Mpath/the_alu/N515 , \UUT/Mpath/the_alu/N514 ,
         \UUT/Mpath/the_alu/N513 , \UUT/Mpath/the_alu/N512 ,
         \UUT/Mpath/the_alu/N511 , \UUT/Mpath/the_alu/N509 ,
         \UUT/Mpath/the_alu/N508 , \UUT/Mpath/the_alu/N507 ,
         \UUT/Mpath/the_alu/N506 , \UUT/Mpath/the_alu/N505 ,
         \UUT/Mpath/the_alu/N503 , \UUT/Mpath/the_alu/N502 ,
         \UUT/Mpath/the_alu/N501 , \UUT/Mpath/the_alu/N500 ,
         \UUT/Mpath/the_alu/N499 , \UUT/Mpath/the_alu/N498 ,
         \UUT/Mpath/the_alu/N497 , \UUT/Mpath/the_alu/N496 ,
         \UUT/Mpath/the_alu/N495 , \UUT/Mpath/the_alu/N494 ,
         \UUT/Mpath/the_alu/N493 , \UUT/Mpath/the_alu/N492 ,
         \UUT/Mpath/the_alu/N491 , \UUT/Mpath/the_alu/N490 ,
         \UUT/Mpath/the_alu/N489 , \UUT/Mpath/the_alu/N488 ,
         \UUT/Mpath/the_alu/N487 , \UUT/Mpath/the_alu/N486 ,
         \UUT/Mpath/the_alu/N485 , \UUT/Mpath/the_alu/N484 ,
         \UUT/Mpath/the_alu/N483 , \UUT/Mpath/the_alu/N482 ,
         \UUT/Mpath/the_alu/N481 , \UUT/Mpath/the_alu/N480 ,
         \UUT/Mpath/the_alu/N479 , \UUT/Mpath/the_alu/N478 ,
         \UUT/Mpath/the_alu/N477 , \UUT/Mpath/the_alu/N476 ,
         \UUT/Mpath/the_alu/N475 , \UUT/Mpath/the_alu/N474 ,
         \UUT/Mpath/the_alu/N473 , \UUT/Mpath/the_alu/N472 ,
         \UUT/Mpath/the_alu/N471 , \UUT/Mpath/the_alu/N470 ,
         \UUT/Mpath/the_alu/N469 , \UUT/Mpath/the_alu/N468 ,
         \UUT/Mpath/the_alu/N467 , \UUT/Mpath/the_alu/N466 ,
         \UUT/Mpath/the_alu/N453 , \UUT/Mpath/the_alu/N221 ,
         \UUT/Mpath/the_alu/N219 , \UUT/Mpath/the_alu/N218 ,
         \UUT/Mpath/the_alu/N217 , \UUT/Mpath/the_alu/N216 ,
         \UUT/Mpath/the_alu/N215 , \UUT/Mpath/the_alu/N214 ,
         \UUT/Mpath/the_alu/N213 , \UUT/Mpath/the_alu/N212 ,
         \UUT/Mpath/the_alu/N211 , \UUT/Mpath/the_alu/N210 ,
         \UUT/Mpath/the_alu/N209 , \UUT/Mpath/the_alu/N208 ,
         \UUT/Mpath/the_alu/N207 , \UUT/Mpath/the_alu/N206 ,
         \UUT/Mpath/the_alu/N205 , \UUT/Mpath/the_alu/N204 ,
         \UUT/Mpath/the_alu/N203 , \UUT/Mpath/the_alu/N202 ,
         \UUT/Mpath/the_alu/N201 , \UUT/Mpath/the_alu/N200 ,
         \UUT/Mpath/the_alu/N199 , \UUT/Mpath/the_alu/N198 ,
         \UUT/Mpath/the_alu/N197 , \UUT/Mpath/the_alu/N196 ,
         \UUT/Mpath/the_alu/N195 , \UUT/Mpath/the_alu/N194 ,
         \UUT/Mpath/the_alu/N193 , \UUT/Mpath/the_alu/N192 ,
         \UUT/Mpath/the_alu/N191 , \UUT/Mpath/the_alu/N190 ,
         \UUT/Mpath/the_alu/N189 , \UUT/Mpath/the_alu/N187 ,
         \UUT/Mpath/the_alu/N186 , \UUT/Mpath/the_alu/N185 ,
         \UUT/Mpath/the_alu/N184 , \UUT/Mpath/the_alu/N183 ,
         \UUT/Mpath/the_alu/N182 , \UUT/Mpath/the_alu/N181 ,
         \UUT/Mpath/the_alu/N180 , \UUT/Mpath/the_alu/N179 ,
         \UUT/Mpath/the_alu/N178 , \UUT/Mpath/the_alu/N177 ,
         \UUT/Mpath/the_alu/N176 , \UUT/Mpath/the_alu/N175 ,
         \UUT/Mpath/the_alu/N174 , \UUT/Mpath/the_alu/N173 ,
         \UUT/Mpath/the_alu/N172 , \UUT/Mpath/the_alu/N171 ,
         \UUT/Mpath/the_alu/N170 , \UUT/Mpath/the_alu/N169 ,
         \UUT/Mpath/the_alu/N168 , \UUT/Mpath/the_alu/N167 ,
         \UUT/Mpath/the_alu/N166 , \UUT/Mpath/the_alu/N165 ,
         \UUT/Mpath/the_alu/N164 , \UUT/Mpath/the_alu/N163 ,
         \UUT/Mpath/the_alu/N162 , \UUT/Mpath/the_alu/N161 ,
         \UUT/Mpath/the_alu/N160 , \UUT/Mpath/the_alu/N159 ,
         \UUT/Mpath/the_alu/N158 , \UUT/Mpath/the_alu/N157 ,
         \UUT/Mpath/the_alu/N155 , \UUT/Mpath/the_alu/N154 ,
         \UUT/Mpath/the_alu/N153 , \UUT/Mpath/the_alu/N152 ,
         \UUT/Mpath/the_alu/N151 , \UUT/Mpath/the_alu/N150 ,
         \UUT/Mpath/the_alu/N149 , \UUT/Mpath/the_alu/N148 ,
         \UUT/Mpath/the_alu/N147 , \UUT/Mpath/the_alu/N146 ,
         \UUT/Mpath/the_alu/N145 , \UUT/Mpath/the_alu/N144 ,
         \UUT/Mpath/the_alu/N143 , \UUT/Mpath/the_alu/N142 ,
         \UUT/Mpath/the_alu/N141 , \UUT/Mpath/the_alu/N140 ,
         \UUT/Mpath/the_alu/N139 , \UUT/Mpath/the_alu/N138 ,
         \UUT/Mpath/the_alu/N137 , \UUT/Mpath/the_alu/N136 ,
         \UUT/Mpath/the_alu/N135 , \UUT/Mpath/the_alu/N134 ,
         \UUT/Mpath/the_alu/N133 , \UUT/Mpath/the_alu/N132 ,
         \UUT/Mpath/the_alu/N131 , \UUT/Mpath/the_alu/N130 ,
         \UUT/Mpath/the_alu/N129 , \UUT/Mpath/the_alu/N128 ,
         \UUT/Mpath/the_alu/N127 , \UUT/Mpath/the_alu/N126 ,
         \UUT/Mpath/the_alu/N125 , \UUT/Mpath/the_alu/N123 ,
         \UUT/Mpath/the_alu/N122 , \UUT/Mpath/the_alu/N121 ,
         \UUT/Mpath/the_alu/N120 , \UUT/Mpath/the_alu/N119 ,
         \UUT/Mpath/the_alu/N118 , \UUT/Mpath/the_alu/N117 ,
         \UUT/Mpath/the_alu/N116 , \UUT/Mpath/the_alu/N115 ,
         \UUT/Mpath/the_alu/N114 , \UUT/Mpath/the_alu/N113 ,
         \UUT/Mpath/the_alu/N112 , \UUT/Mpath/the_alu/N111 ,
         \UUT/Mpath/the_alu/N110 , \UUT/Mpath/the_alu/N109 ,
         \UUT/Mpath/the_alu/N108 , \UUT/Mpath/the_alu/N107 ,
         \UUT/Mpath/the_alu/N106 , \UUT/Mpath/the_alu/N105 ,
         \UUT/Mpath/the_alu/N104 , \UUT/Mpath/the_alu/N103 ,
         \UUT/Mpath/the_alu/N102 , \UUT/Mpath/the_alu/N101 ,
         \UUT/Mpath/the_alu/N100 , \UUT/Mpath/the_alu/N99 ,
         \UUT/Mpath/the_alu/N98 , \UUT/Mpath/the_alu/N97 ,
         \UUT/Mpath/the_alu/N96 , \UUT/Mpath/the_alu/N95 ,
         \UUT/Mpath/the_alu/N94 , \UUT/Mpath/the_alu/N93 ,
         \UUT/Mpath/the_alu/N91 , \UUT/Mpath/the_alu/diff[0] ,
         \UUT/Mpath/the_alu/diff[1] , \UUT/Mpath/the_alu/diff[2] ,
         \UUT/Mpath/the_alu/diff[3] , \UUT/Mpath/the_alu/diff[4] ,
         \UUT/Mpath/the_alu/diff[5] , \UUT/Mpath/the_alu/diff[6] ,
         \UUT/Mpath/the_alu/diff[7] , \UUT/Mpath/the_alu/diff[8] ,
         \UUT/Mpath/the_alu/diff[9] , \UUT/Mpath/the_alu/diff[10] ,
         \UUT/Mpath/the_alu/diff[11] , \UUT/Mpath/the_alu/diff[12] ,
         \UUT/Mpath/the_alu/diff[13] , \UUT/Mpath/the_alu/diff[14] ,
         \UUT/Mpath/the_alu/diff[15] , \UUT/Mpath/the_alu/diff[16] ,
         \UUT/Mpath/the_alu/diff[17] , \UUT/Mpath/the_alu/diff[18] ,
         \UUT/Mpath/the_alu/diff[19] , \UUT/Mpath/the_alu/diff[20] ,
         \UUT/Mpath/the_alu/diff[21] , \UUT/Mpath/the_alu/diff[22] ,
         \UUT/Mpath/the_alu/diff[23] , \UUT/Mpath/the_alu/diff[24] ,
         \UUT/Mpath/the_alu/diff[25] , \UUT/Mpath/the_alu/diff[26] ,
         \UUT/Mpath/the_alu/diff[27] , \UUT/Mpath/the_alu/diff[28] ,
         \UUT/Mpath/the_alu/diff[29] , \UUT/Mpath/the_alu/diff[30] ,
         \UUT/Mpath/the_alu/diff[31] , \UUT/Mpath/the_alu/sum[0] ,
         \UUT/Mpath/the_alu/sum[1] , \UUT/Mpath/the_alu/sum[2] ,
         \UUT/Mpath/the_alu/sum[3] , \UUT/Mpath/the_alu/sum[4] ,
         \UUT/Mpath/the_alu/sum[5] , \UUT/Mpath/the_alu/sum[6] ,
         \UUT/Mpath/the_alu/sum[7] , \UUT/Mpath/the_alu/sum[8] ,
         \UUT/Mpath/the_alu/sum[9] , \UUT/Mpath/the_alu/sum[10] ,
         \UUT/Mpath/the_alu/sum[11] , \UUT/Mpath/the_alu/sum[12] ,
         \UUT/Mpath/the_alu/sum[13] , \UUT/Mpath/the_alu/sum[14] ,
         \UUT/Mpath/the_alu/sum[15] , \UUT/Mpath/the_alu/sum[16] ,
         \UUT/Mpath/the_alu/sum[17] , \UUT/Mpath/the_alu/sum[18] ,
         \UUT/Mpath/the_alu/sum[19] , \UUT/Mpath/the_alu/sum[20] ,
         \UUT/Mpath/the_alu/sum[21] , \UUT/Mpath/the_alu/sum[22] ,
         \UUT/Mpath/the_alu/sum[23] , \UUT/Mpath/the_alu/sum[24] ,
         \UUT/Mpath/the_alu/sum[25] , \UUT/Mpath/the_alu/sum[26] ,
         \UUT/Mpath/the_alu/sum[27] , \UUT/Mpath/the_alu/sum[28] ,
         \UUT/Mpath/the_alu/sum[29] , \UUT/Mpath/the_alu/sum[30] ,
         \UUT/Mpath/the_alu/sum[31] , \UUT/Mpath/the_alu/N84 ,
         \UUT/Mpath/the_alu/N83 , \UUT/Mpath/the_alu/N82 ,
         \UUT/Mpath/the_alu/N81 , \UUT/Mpath/the_alu/N80 ,
         \UUT/Mpath/the_alu/N79 , \UUT/Mpath/the_alu/N78 ,
         \UUT/Mpath/the_alu/N77 , \UUT/Mpath/the_alu/N76 ,
         \UUT/Mpath/the_alu/N75 , \UUT/Mpath/the_alu/N74 ,
         \UUT/Mpath/the_alu/N73 , \UUT/Mpath/the_alu/N72 ,
         \UUT/Mpath/the_alu/N71 , \UUT/Mpath/the_alu/N70 ,
         \UUT/Mpath/the_alu/N69 , \UUT/Mpath/the_alu/N68 ,
         \UUT/Mpath/the_alu/N67 , \UUT/Mpath/the_alu/N66 ,
         \UUT/Mpath/the_alu/N65 , \UUT/Mpath/the_alu/N64 ,
         \UUT/Mpath/the_alu/N63 , \UUT/Mpath/the_alu/N62 ,
         \UUT/Mpath/the_alu/N61 , \UUT/Mpath/the_alu/N60 ,
         \UUT/Mpath/the_alu/N59 , \UUT/Mpath/the_alu/N58 ,
         \UUT/Mpath/the_alu/N57 , \UUT/Mpath/the_alu/N56 ,
         \UUT/Mpath/the_alu/N55 , \UUT/Mpath/the_alu/N54 ,
         \UUT/Mpath/the_alu/N53 , \UUT/Mpath/the_alu/N52 ,
         \UUT/Mpath/the_alu/N51 , \UUT/Mpath/the_alu/N50 ,
         \UUT/Mpath/the_alu/N49 , \UUT/Mpath/the_alu/N48 ,
         \UUT/Mpath/the_alu/N47 , \UUT/Mpath/the_alu/N46 ,
         \UUT/Mpath/the_alu/N45 , \UUT/Mpath/the_alu/N44 ,
         \UUT/Mpath/the_alu/N43 , \UUT/Mpath/the_alu/N42 ,
         \UUT/Mpath/the_alu/N41 , \UUT/Mpath/the_alu/N40 ,
         \UUT/Mpath/the_alu/N39 , \UUT/Mpath/the_alu/N38 ,
         \UUT/Mpath/the_alu/N37 , \UUT/Mpath/the_alu/N36 ,
         \UUT/Mpath/the_alu/N35 , \UUT/Mpath/the_alu/N34 ,
         \UUT/Mpath/the_alu/N33 , \UUT/Mpath/the_alu/N32 ,
         \UUT/Mpath/the_alu/N31 , \UUT/Mpath/the_alu/N30 ,
         \UUT/Mpath/the_alu/N29 , \UUT/Mpath/the_alu/N28 ,
         \UUT/Mpath/the_alu/N27 , \UUT/Mpath/the_alu/N26 ,
         \UUT/Mpath/the_alu/N25 , \UUT/Mpath/the_alu/N24 ,
         \UUT/Mpath/the_alu/N23 , \UUT/Mpath/the_alu/N22 ,
         \UUT/Mpath/the_alu/N21 , \UUT/Mpath/the_shift/N118 ,
         \UUT/Mpath/the_shift/N117 , \UUT/Mpath/the_shift/N116 ,
         \UUT/Mpath/the_shift/N115 , \UUT/Mpath/the_shift/N114 ,
         \UUT/Mpath/the_shift/N113 , \UUT/Mpath/the_shift/N112 ,
         \UUT/Mpath/the_shift/N111 , \UUT/Mpath/the_shift/N110 ,
         \UUT/Mpath/the_shift/N109 , \UUT/Mpath/the_shift/N108 ,
         \UUT/Mpath/the_shift/N107 , \UUT/Mpath/the_shift/N106 ,
         \UUT/Mpath/the_shift/N105 , \UUT/Mpath/the_shift/N104 ,
         \UUT/Mpath/the_mult/N313 , \UUT/Mpath/the_mult/N312 ,
         \UUT/Mpath/the_mult/N311 , \UUT/Mpath/the_mult/N298 ,
         \UUT/Mpath/the_mult/N297 , \UUT/Mpath/the_mult/N296 ,
         \UUT/Mpath/the_mult/N295 , \UUT/Mpath/the_mult/N294 ,
         \UUT/Mpath/the_mult/N293 , \UUT/Mpath/the_mult/N292 ,
         \UUT/Mpath/the_mult/N291 , \UUT/Mpath/the_mult/N290 ,
         \UUT/Mpath/the_mult/N289 , \UUT/Mpath/the_mult/N288 ,
         \UUT/Mpath/the_mult/N287 , \UUT/Mpath/the_mult/N285 ,
         \UUT/Mpath/the_mult/N284 , \UUT/Mpath/the_mult/N283 ,
         \UUT/Mpath/the_mult/N282 , \UUT/Mpath/the_mult/N281 ,
         \UUT/Mpath/the_mult/N280 , \UUT/Mpath/the_mult/N279 ,
         \UUT/Mpath/the_mult/N278 , \UUT/Mpath/the_mult/N277 ,
         \UUT/Mpath/the_mult/N276 , \UUT/Mpath/the_mult/N275 ,
         \UUT/Mpath/the_mult/N274 , \UUT/Mpath/the_mult/N273 ,
         \UUT/Mpath/the_mult/N272 , \UUT/Mpath/the_mult/N271 ,
         \UUT/Mpath/the_mult/N270 , \UUT/Mpath/the_mult/N269 ,
         \UUT/Mpath/the_mult/N268 , \UUT/Mpath/the_mult/N267 ,
         \UUT/Mpath/the_mult/N266 , \UUT/Mpath/the_mult/N265 ,
         \UUT/Mpath/the_mult/N264 , \UUT/Mpath/the_mult/N263 ,
         \UUT/Mpath/the_mult/N262 , \UUT/Mpath/the_mult/N261 ,
         \UUT/Mpath/the_mult/N260 , \UUT/Mpath/the_mult/N259 ,
         \UUT/Mpath/the_mult/N258 , \UUT/Mpath/the_mult/N257 ,
         \UUT/Mpath/the_mult/N255 , \UUT/Mpath/the_mult/N254 ,
         \UUT/Mpath/the_mult/N253 , \UUT/Mpath/the_mult/N252 ,
         \UUT/Mpath/the_mult/N251 , \UUT/Mpath/the_mult/N244 ,
         \UUT/Mpath/the_mult/N231 , \UUT/Mpath/the_mult/N230 ,
         \UUT/Mpath/the_mult/N229 , \UUT/Mpath/the_mult/N227 ,
         \UUT/Mpath/the_mult/N226 , \UUT/Mpath/the_mult/N225 ,
         \UUT/Mpath/the_mult/N224 , \UUT/Mpath/the_mult/N223 ,
         \UUT/Mpath/the_mult/N222 , \UUT/Mpath/the_mult/N221 ,
         \UUT/Mpath/the_mult/N220 , \UUT/Mpath/the_mult/N216 ,
         \UUT/Mpath/the_mult/N215 , \UUT/Mpath/the_mult/N214 ,
         \UUT/Mpath/the_mult/N213 , \UUT/Mpath/the_mult/N212 ,
         \UUT/Mpath/the_mult/N198 , \UUT/Mpath/the_mult/N197 ,
         \UUT/Mpath/the_mult/N196 , \UUT/Mpath/the_mult/N195 ,
         \UUT/Mpath/the_mult/N194 , \UUT/Mpath/the_mult/N193 ,
         \UUT/Mpath/the_mult/N192 , \UUT/Mpath/the_mult/acc_out[0] ,
         \UUT/Mpath/the_mult/acc_out[1] , \UUT/Mpath/the_mult/acc_out[2] ,
         \UUT/Mpath/the_mult/acc_out[3] , \UUT/Mpath/the_mult/acc_out[4] ,
         \UUT/Mpath/the_mult/acc_out[5] , \UUT/Mpath/the_mult/acc_out[6] ,
         \UUT/Mpath/the_mult/acc_out[7] , \UUT/Mpath/the_mult/acc_out[8] ,
         \UUT/Mpath/the_mult/acc_out[9] , \UUT/Mpath/the_mult/acc_out[10] ,
         \UUT/Mpath/the_mult/acc_out[11] , \UUT/Mpath/the_mult/acc_out[12] ,
         \UUT/Mpath/the_mult/acc_out[13] , \UUT/Mpath/the_mult/acc_out[14] ,
         \UUT/Mpath/the_mult/acc_out[15] , \UUT/Mpath/the_mult/acc_out[16] ,
         \UUT/Mpath/the_mult/acc_out[17] , \UUT/Mpath/the_mult/acc_out[18] ,
         \UUT/Mpath/the_mult/acc_out[19] , \UUT/Mpath/the_mult/acc_out[20] ,
         \UUT/Mpath/the_mult/acc_out[21] , \UUT/Mpath/the_mult/acc_out[22] ,
         \UUT/Mpath/the_mult/acc_out[23] , \UUT/Mpath/the_mult/acc_out[24] ,
         \UUT/Mpath/the_mult/acc_out[25] , \UUT/Mpath/the_mult/acc_out[26] ,
         \UUT/Mpath/the_mult/acc_out[27] , \UUT/Mpath/the_mult/acc_out[28] ,
         \UUT/Mpath/the_mult/acc_out[29] , \UUT/Mpath/the_mult/acc_out[30] ,
         \UUT/Mpath/the_mult/acc_out[31] , \UUT/Mpath/the_mult/acc_out[32] ,
         \UUT/Mpath/the_mult/acc_out[33] , \UUT/Mpath/the_mult/acc_out[34] ,
         \UUT/Mpath/the_mult/acc_out[35] , \UUT/Mpath/the_mult/acc_out[36] ,
         \UUT/Mpath/the_mult/acc_out[37] , \UUT/Mpath/the_mult/acc_out[38] ,
         \UUT/Mpath/the_mult/acc_out[39] , \UUT/Mpath/the_mult/acc_out[40] ,
         \UUT/Mpath/the_mult/acc_out[41] , \UUT/Mpath/the_mult/acc_out[42] ,
         \UUT/Mpath/the_mult/acc_out[43] , \UUT/Mpath/the_mult/acc_out[44] ,
         \UUT/Mpath/the_mult/acc_out[45] , \UUT/Mpath/the_mult/acc_out[46] ,
         \UUT/Mpath/the_mult/acc_out[47] , \UUT/Mpath/the_mult/acc_out[48] ,
         \UUT/Mpath/the_mult/acc_out[49] , \UUT/Mpath/the_mult/acc_out[50] ,
         \UUT/Mpath/the_mult/acc_out[51] , \UUT/Mpath/the_mult/acc_out[52] ,
         \UUT/Mpath/the_mult/acc_out[53] , \UUT/Mpath/the_mult/acc_out[54] ,
         \UUT/Mpath/the_mult/acc_out[55] , \UUT/Mpath/the_mult/acc_out[56] ,
         \UUT/Mpath/the_mult/acc_out[57] , \UUT/Mpath/the_mult/acc_out[58] ,
         \UUT/Mpath/the_mult/acc_out[59] , \UUT/Mpath/the_mult/acc_out[60] ,
         \UUT/Mpath/the_mult/acc_out[61] , \UUT/Mpath/the_mult/acc_out[62] ,
         \UUT/Mpath/the_mult/acc_out[63] , \UUT/Mpath/the_mult/Mult_out[0] ,
         \UUT/Mpath/the_mult/Mult_out[1] , \UUT/Mpath/the_mult/Mult_out[2] ,
         \UUT/Mpath/the_mult/Mult_out[3] , \UUT/Mpath/the_mult/Mult_out[4] ,
         \UUT/Mpath/the_mult/Mult_out[5] , \UUT/Mpath/the_mult/Mult_out[6] ,
         \UUT/Mpath/the_mult/Mult_out[7] , \UUT/Mpath/the_mult/Mult_out[8] ,
         \UUT/Mpath/the_mult/Mult_out[9] , \UUT/Mpath/the_mult/Mult_out[10] ,
         \UUT/Mpath/the_mult/Mult_out[11] , \UUT/Mpath/the_mult/Mult_out[12] ,
         \UUT/Mpath/the_mult/Mult_out[13] , \UUT/Mpath/the_mult/Mult_out[14] ,
         \UUT/Mpath/the_mult/Mult_out[15] , \UUT/Mpath/the_mult/Mult_out[16] ,
         \UUT/Mpath/the_mult/Mult_out[17] , \UUT/Mpath/the_mult/Mult_out[18] ,
         \UUT/Mpath/the_mult/Mult_out[19] , \UUT/Mpath/the_mult/Mult_out[20] ,
         \UUT/Mpath/the_mult/Mult_out[21] , \UUT/Mpath/the_mult/Mult_out[22] ,
         \UUT/Mpath/the_mult/Mult_out[23] , \UUT/Mpath/the_mult/Mult_out[24] ,
         \UUT/Mpath/the_mult/Mult_out[25] , \UUT/Mpath/the_mult/Mult_out[26] ,
         \UUT/Mpath/the_mult/Mult_out[27] , \UUT/Mpath/the_mult/Mult_out[28] ,
         \UUT/Mpath/the_mult/Mult_out[29] , \UUT/Mpath/the_mult/Mult_out[30] ,
         \UUT/Mpath/the_mult/Mult_out[31] , \UUT/Mpath/the_mult/Mult_out[32] ,
         \UUT/Mpath/the_mult/Mult_out[33] , \UUT/Mpath/the_mult/Mult_out[34] ,
         \UUT/Mpath/the_mult/Mult_out[35] , \UUT/Mpath/the_mult/Mult_out[36] ,
         \UUT/Mpath/the_mult/Mult_out[37] , \UUT/Mpath/the_mult/Mult_out[38] ,
         \UUT/Mpath/the_mult/Mult_out[39] , \UUT/Mpath/the_mult/Mult_out[40] ,
         \UUT/Mpath/the_mult/Mult_out[41] , \UUT/Mpath/the_mult/Mult_out[42] ,
         \UUT/Mpath/the_mult/Mult_out[43] , \UUT/Mpath/the_mult/Mult_out[44] ,
         \UUT/Mpath/the_mult/Mult_out[45] , \UUT/Mpath/the_mult/Mult_out[46] ,
         \UUT/Mpath/the_mult/Mult_out[47] , \UUT/Mpath/the_mult/Mult_out[48] ,
         \UUT/Mpath/the_mult/Mult_out[49] , \UUT/Mpath/the_mult/Mult_out[50] ,
         \UUT/Mpath/the_mult/Mult_out[51] , \UUT/Mpath/the_mult/Mult_out[52] ,
         \UUT/Mpath/the_mult/Mult_out[53] , \UUT/Mpath/the_mult/Mult_out[54] ,
         \UUT/Mpath/the_mult/Mult_out[55] , \UUT/Mpath/the_mult/Mult_out[56] ,
         \UUT/Mpath/the_mult/Mult_out[57] , \UUT/Mpath/the_mult/Mult_out[58] ,
         \UUT/Mpath/the_mult/Mult_out[59] , \UUT/Mpath/the_mult/Mult_out[60] ,
         \UUT/Mpath/the_mult/Mult_out[61] , \UUT/Mpath/the_mult/Mult_out[62] ,
         \UUT/Mpath/the_mult/Mult_out[63] ,
         \UUT/Mpath/the_mult/m_mul_command[0] ,
         \UUT/Mpath/the_mult/m_mul_command[1] ,
         \UUT/Mpath/the_mult/m_mul_command[2] ,
         \UUT/Mpath/the_mult/m_mul_command[3] ,
         \UUT/Mpath/the_mult/m_mul_command[4] ,
         \UUT/Mpath/the_mult/m_mul_command[5] ,
         \UUT/Mpath/the_mult/x_mult_out[0] ,
         \UUT/Mpath/the_mult/x_mult_out[1] ,
         \UUT/Mpath/the_mult/x_mult_out[2] ,
         \UUT/Mpath/the_mult/x_mult_out[3] ,
         \UUT/Mpath/the_mult/x_mult_out[4] ,
         \UUT/Mpath/the_mult/x_mult_out[5] ,
         \UUT/Mpath/the_mult/x_mult_out[6] ,
         \UUT/Mpath/the_mult/x_mult_out[7] ,
         \UUT/Mpath/the_mult/x_mult_out[8] ,
         \UUT/Mpath/the_mult/x_mult_out[9] ,
         \UUT/Mpath/the_mult/x_mult_out[10] ,
         \UUT/Mpath/the_mult/x_mult_out[11] ,
         \UUT/Mpath/the_mult/x_mult_out[12] ,
         \UUT/Mpath/the_mult/x_mult_out[13] ,
         \UUT/Mpath/the_mult/x_mult_out[14] ,
         \UUT/Mpath/the_mult/x_mult_out[15] ,
         \UUT/Mpath/the_mult/x_mult_out[16] ,
         \UUT/Mpath/the_mult/x_mult_out[17] ,
         \UUT/Mpath/the_mult/x_mult_out[18] ,
         \UUT/Mpath/the_mult/x_mult_out[19] ,
         \UUT/Mpath/the_mult/x_mult_out[20] ,
         \UUT/Mpath/the_mult/x_mult_out[21] ,
         \UUT/Mpath/the_mult/x_mult_out[22] ,
         \UUT/Mpath/the_mult/x_mult_out[23] ,
         \UUT/Mpath/the_mult/x_mult_out[24] ,
         \UUT/Mpath/the_mult/x_mult_out[25] ,
         \UUT/Mpath/the_mult/x_mult_out[26] ,
         \UUT/Mpath/the_mult/x_mult_out[27] ,
         \UUT/Mpath/the_mult/x_mult_out[28] ,
         \UUT/Mpath/the_mult/x_mult_out[29] ,
         \UUT/Mpath/the_mult/x_mult_out[30] ,
         \UUT/Mpath/the_mult/x_mult_out[31] ,
         \UUT/Mpath/the_mult/x_mult_out[32] ,
         \UUT/Mpath/the_mult/x_mult_out[33] ,
         \UUT/Mpath/the_mult/x_mult_out[34] ,
         \UUT/Mpath/the_mult/x_mult_out[35] ,
         \UUT/Mpath/the_mult/x_mult_out[36] ,
         \UUT/Mpath/the_mult/x_mult_out[37] ,
         \UUT/Mpath/the_mult/x_mult_out[38] ,
         \UUT/Mpath/the_mult/x_mult_out[39] ,
         \UUT/Mpath/the_mult/x_mult_out[40] ,
         \UUT/Mpath/the_mult/x_mult_out[41] ,
         \UUT/Mpath/the_mult/x_mult_out[42] ,
         \UUT/Mpath/the_mult/x_mult_out[43] ,
         \UUT/Mpath/the_mult/x_mult_out[44] ,
         \UUT/Mpath/the_mult/x_mult_out[45] ,
         \UUT/Mpath/the_mult/x_mult_out[46] ,
         \UUT/Mpath/the_mult/x_mult_out[47] ,
         \UUT/Mpath/the_mult/x_mult_out[48] ,
         \UUT/Mpath/the_mult/x_mult_out[49] ,
         \UUT/Mpath/the_mult/x_mult_out[50] ,
         \UUT/Mpath/the_mult/x_mult_out[51] ,
         \UUT/Mpath/the_mult/x_mult_out[52] ,
         \UUT/Mpath/the_mult/x_mult_out[53] ,
         \UUT/Mpath/the_mult/x_mult_out[54] ,
         \UUT/Mpath/the_mult/x_mult_out[55] ,
         \UUT/Mpath/the_mult/x_mult_out[56] ,
         \UUT/Mpath/the_mult/x_mult_out[57] ,
         \UUT/Mpath/the_mult/x_mult_out[58] ,
         \UUT/Mpath/the_mult/x_mult_out[59] ,
         \UUT/Mpath/the_mult/x_mult_out[60] ,
         \UUT/Mpath/the_mult/x_mult_out[61] ,
         \UUT/Mpath/the_mult/x_mult_out[62] ,
         \UUT/Mpath/the_mult/x_mult_out[63] ,
         \UUT/Mpath/the_mult/x_mul_command[0] ,
         \UUT/Mpath/the_mult/x_mul_command[1] ,
         \UUT/Mpath/the_mult/x_mul_command[2] ,
         \UUT/Mpath/the_mult/x_mul_command[3] ,
         \UUT/Mpath/the_mult/x_mul_command[4] ,
         \UUT/Mpath/the_mult/x_mul_command[5] ,
         \UUT/Mpath/the_mult/x_operand1[0] ,
         \UUT/Mpath/the_mult/x_operand1[1] ,
         \UUT/Mpath/the_mult/x_operand1[2] ,
         \UUT/Mpath/the_mult/x_operand1[3] ,
         \UUT/Mpath/the_mult/x_operand1[4] ,
         \UUT/Mpath/the_mult/x_operand1[5] ,
         \UUT/Mpath/the_mult/x_operand1[6] ,
         \UUT/Mpath/the_mult/x_operand1[7] ,
         \UUT/Mpath/the_mult/x_operand1[8] ,
         \UUT/Mpath/the_mult/x_operand1[9] ,
         \UUT/Mpath/the_mult/x_operand1[10] ,
         \UUT/Mpath/the_mult/x_operand1[11] ,
         \UUT/Mpath/the_mult/x_operand1[12] ,
         \UUT/Mpath/the_mult/x_operand1[13] ,
         \UUT/Mpath/the_mult/x_operand1[14] ,
         \UUT/Mpath/the_mult/x_operand1[15] ,
         \UUT/Mpath/the_mult/x_operand1[16] ,
         \UUT/Mpath/the_mult/x_operand1[17] ,
         \UUT/Mpath/the_mult/x_operand1[18] ,
         \UUT/Mpath/the_mult/x_operand1[19] ,
         \UUT/Mpath/the_mult/x_operand1[20] ,
         \UUT/Mpath/the_mult/x_operand1[21] ,
         \UUT/Mpath/the_mult/x_operand1[22] ,
         \UUT/Mpath/the_mult/x_operand1[23] ,
         \UUT/Mpath/the_mult/x_operand1[24] ,
         \UUT/Mpath/the_mult/x_operand1[25] ,
         \UUT/Mpath/the_mult/x_operand1[26] ,
         \UUT/Mpath/the_mult/x_operand1[27] ,
         \UUT/Mpath/the_mult/x_operand1[28] ,
         \UUT/Mpath/the_mult/x_operand1[29] ,
         \UUT/Mpath/the_mult/x_operand1[30] ,
         \UUT/Mpath/the_mult/x_operand1[31] , \UUT/Mpath/the_memhandle/N244 ,
         \UUT/Mpath/the_memhandle/N243 , \UUT/Mpath/the_memhandle/N242 ,
         \UUT/Mpath/the_memhandle/N241 , \UUT/Mpath/the_memhandle/N240 ,
         \UUT/Mpath/the_memhandle/N239 , \UUT/Mpath/the_memhandle/N238 ,
         \UUT/Mpath/the_memhandle/N237 , \UUT/Mpath/the_memhandle/N236 ,
         \UUT/Mpath/the_memhandle/N235 , \UUT/Mpath/the_memhandle/N234 ,
         \UUT/Mpath/the_memhandle/N120 , \UUT/Mpath/the_memhandle/N86 ,
         \UUT/Mpath/the_memhandle/N77 , \UUT/Mpath/the_memhandle/N76 ,
         \UUT/Mpath/the_memhandle/N74 , \UUT/Mpath/the_memhandle/N72 ,
         \UUT/Mpath/the_memhandle/N39 , \UUT/Mpath/the_memhandle/N38 ,
         \UUT/Mpath/the_memhandle/N37 , \UUT/Mpath/the_memhandle/N36 ,
         \UUT/Mpath/the_memhandle/N34 , \UUT/Mpath/the_memhandle/smdr_out[8] ,
         \UUT/Mpath/the_memhandle/smdr_out[9] ,
         \UUT/Mpath/the_memhandle/smdr_out[10] ,
         \UUT/Mpath/the_memhandle/smdr_out[11] ,
         \UUT/Mpath/the_memhandle/smdr_out[12] ,
         \UUT/Mpath/the_memhandle/smdr_out[13] ,
         \UUT/Mpath/the_memhandle/smdr_out[14] ,
         \UUT/Mpath/the_memhandle/smdr_out[15] ,
         \UUT/Mpath/the_memhandle/smdr_out[16] ,
         \UUT/Mpath/the_memhandle/smdr_out[17] ,
         \UUT/Mpath/the_memhandle/smdr_out[18] ,
         \UUT/Mpath/the_memhandle/smdr_out[19] ,
         \UUT/Mpath/the_memhandle/smdr_out[20] ,
         \UUT/Mpath/the_memhandle/smdr_out[21] ,
         \UUT/Mpath/the_memhandle/smdr_out[22] ,
         \UUT/Mpath/the_memhandle/smdr_out[23] ,
         \UUT/Mpath/the_memhandle/smdr_out[24] ,
         \UUT/Mpath/the_memhandle/smdr_out[25] ,
         \UUT/Mpath/the_memhandle/smdr_out[26] ,
         \UUT/Mpath/the_memhandle/smdr_out[27] ,
         \UUT/Mpath/the_memhandle/smdr_out[28] ,
         \UUT/Mpath/the_memhandle/smdr_out[29] ,
         \UUT/Mpath/the_memhandle/smdr_out[30] ,
         \UUT/Mpath/the_memhandle/smdr_out[31] , \localbus/N338 ,
         \localbus/N337 , \localbus/N336 , \localbus/N335 , \localbus/N334 ,
         \localbus/N333 , \localbus/N331 , \localbus/N329 , \localbus/N328 ,
         \localbus/N327 , \localbus/N326 , \localbus/N325 , \localbus/N324 ,
         \localbus/N323 , \localbus/N322 , \localbus/N321 , \localbus/N320 ,
         \localbus/N319 , \localbus/N318 , \localbus/N297 , \localbus/N296 ,
         \localbus/N293 , \localbus/N271 , \localbus/N270 , \localbus/N268 ,
         \localbus/N267 , \localbus/N266 , \localbus/N265 , \localbus/N263 ,
         \localbus/N262 , \localbus/N261 , \localbus/N260 , \localbus/N258 ,
         \localbus/N257 , \localbus/N256 , \localbus/N255 , \localbus/N254 ,
         \localbus/N252 , \localbus/N251 , \localbus/N250 , \localbus/N229 ,
         \localbus/N228 , \localbus/N227 , \localbus/N226 , \localbus/N225 ,
         \localbus/N219 , \localbus/N218 , \localbus/N217 , \localbus/N215 ,
         \localbus/N214 , \localbus/N199 , \localbus/N95 , \localbus/N93 ,
         \localbus/c2_op[OP][1] , \localbus/c2_op[SLAVE][0] ,
         \localbus/c2_op[SLAVE][1] , \localbus/c2_op[SLAVE][2] ,
         \localbus/c2_op[MASTER] , \localbus/N90 , \localbus/N89 ,
         \localbus/N86 , \localbus/N85 , \localbus/N62 , \localbus/N61 ,
         \localbus/N60 , \localbus/N57 , \localbus/N56 , \localbus/N55 ,
         \localbus/N51 , \localbus/c1_addr_outbus[13] ,
         \localbus/c1_addr_outbus[14] , \localbus/c1_addr_outbus[15] ,
         \localbus/c1_addr_outbus[16] , \localbus/c1_addr_outbus[17] ,
         \localbus/c1_addr_outbus[18] , \localbus/c1_addr_outbus[19] ,
         \localbus/c1_addr_outbus[20] , \localbus/c1_addr_outbus[21] ,
         \localbus/c1_addr_outbus[22] , \localbus/c1_addr_outbus[23] ,
         \localbus/c1_addr_outbus[24] , \localbus/c1_addr_outbus[25] ,
         \localbus/c1_addr_outbus[26] , \localbus/c1_addr_outbus[27] ,
         \localbus/c1_addr_outbus[28] , \localbus/c1_addr_outbus[29] ,
         \localbus/c1_addr_outbus[30] , \localbus/N50 , \localbus/N46 ,
         \localbus/c1_op[OP][0] , \localbus/c1_op[OP][1] ,
         \localbus/c1_op[SLAVE][0] , \localbus/c1_op[MASTER] , n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1178, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2639, n2642, n2645, n2648, n2651,
         n2654, n2657, n2660, n2663, n2666, n2668, n2671, n2677, n2679, n2682,
         n2685, n2688, n2691, n2694, n2698, n2725, n2727, n2728, n2729, n2730,
         n2732, n2735, n2737, n2739, n2741, n2748, n2750, n2752, n2754, n2756,
         n2781, n2783, n2784, n2785, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4324, n4325, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4337, n4339, n4340, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5551, n5552, n5553, n5554, n5555, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6048, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         net54953, net54949, net54947, net54945, net54943, net54941, net54939,
         net54937, net54935, net54933, net54931, net54929, net54927, net54925,
         net54923, net54921, net54919, net54917, net54915, net54913, net54911,
         net54909, net54907, net54905, net54903, net54895, net54893, net54891,
         net54889, net54887, net54885, net54883, net54881, net54879, net54877,
         net54875, net54873, net54871, net54869, net54867, net54865, net54863,
         net54861, net54859, net54857, net54855, net54853, net54851, net54849,
         net54847, net54845, net54843, net56414, net87679, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939;
  wire   [31:0] I_DATA_INBUS;
  wire   [31:0] D_ADDR_OUTBUS;
  wire   [31:0] D_DATA_OUTBUS;
  wire   [12:2] dram_addr_outbus;
  wire   [31:0] dram_data_inbus;
  wire   [31:0] dram_data_outbus;
  wire   [31:0] d_select;
  wire   [5:0] \UUT/d_mul_command ;
  wire   [2:0] \UUT/exe_outsel ;
  wire   [2:0] \UUT/shift_op ;
  wire   [23:0] \UUT/jar_in ;
  wire   [31:0] \UUT/branch_regb ;
  wire   [31:0] \UUT/branch_rega ;
  wire   [4:0] \UUT/rd_addr ;
  wire   [4:0] \UUT/rs2_addr ;
  wire   [4:0] \UUT/rs1_addr ;
  wire   [31:0] \UUT/daddr_out ;
  wire   [5:0] \UUT/Mcontrol/x_mul_command ;
  wire   [31:0] \UUT/Mcontrol/d_instr ;
  wire   [31:0] \UUT/Mcontrol/d_sampled_finstr ;
  wire   [23:0] \UUT/Mcontrol/f_currpc ;
  wire   [23:0] \UUT/Mcontrol/Nextpc_decoding/Bta ;
  wire   [1:0] \UUT/Mpath/mem_baddr ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_sll ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_srl ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_sra ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_ror ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_rol ;
  wire   [63:0] \UUT/Mpath/the_mult/Mad_out ;
  wire   [31:0] \UUT/Mpath/the_mult/x_operand2 ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;
  assign BUS_BUSY = 1'b1;
  assign \UUT/Mcontrol/int_reset  = reset;

  SRAM DMem ( .address(dram_addr_outbus), .bit_wen(dram_data_outbus), 
        .data_in({d_select[31], d_select[31], d_select[31], d_select[31], 
        d_select[31], d_select[31], d_select[31], d_select[31], d_select[23], 
        d_select[23], d_select[23], d_select[23], d_select[23], d_select[23], 
        d_select[23], d_select[23], d_select[9], d_select[9], d_select[9], 
        d_select[9], d_select[9], d_select[9], d_select[9], d_select[9], 
        d_select[7], d_select[7], d_select[7], d_select[7], d_select[7], 
        d_select[7], d_select[7], d_select[7]}), .data_out(dram_data_inbus), 
        .clk(CLK), .rdn(dram_mr), .wrn(dram_mw) );
  SRAM IMem ( .address({n6686, n6487, \UUT/Mcontrol/Program_counter/N24 , 
        \UUT/Mcontrol/Program_counter/N22 , \UUT/Mcontrol/Program_counter/N20 , 
        n6649, n6654, n6848, n6855, n6647, \UUT/Mcontrol/Program_counter/N8 }), 
        .bit_wen({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .data_out(I_DATA_INBUS), .clk(CLK), .rdn(iram_rd), .wrn(1'b1) );
  OR2_X2 \localbus/C745  ( .A1(\localbus/c1_op[SLAVE][0] ), .A2(
        \localbus/N227 ), .ZN(\localbus/N214 ) );
  INV_X2 \localbus/I_1  ( .A(\localbus/N214 ), .ZN(\localbus/N215 ) );
  OR2_X2 \localbus/C748  ( .A1(\localbus/c1_op[SLAVE][0] ), .A2(
        \localbus/N227 ), .ZN(\localbus/N217 ) );
  INV_X2 \localbus/I_2  ( .A(\localbus/N217 ), .ZN(\localbus/N218 ) );
  OR2_X2 \localbus/C756  ( .A1(n6637), .A2(\localbus/N227 ), .ZN(
        \localbus/N225 ) );
  INV_X2 \localbus/I_6  ( .A(\localbus/N225 ), .ZN(\localbus/N226 ) );
  OR2_X2 \localbus/C760  ( .A1(n6637), .A2(\localbus/N227 ), .ZN(
        \localbus/N228 ) );
  INV_X2 \localbus/I_7  ( .A(\localbus/N228 ), .ZN(\localbus/N229 ) );
  INV_X2 \localbus/I_16  ( .A(\localbus/c1_op[OP][0] ), .ZN(\localbus/N250 )
         );
  OR2_X2 \localbus/C790  ( .A1(\localbus/N250 ), .A2(\localbus/c1_op[OP][1] ), 
        .ZN(\localbus/N251 ) );
  INV_X2 \localbus/I_17  ( .A(\localbus/N251 ), .ZN(\localbus/N252 ) );
  OR2_X2 \localbus/C793  ( .A1(\localbus/c1_op[SLAVE][0] ), .A2(
        \localbus/N227 ), .ZN(\localbus/N254 ) );
  INV_X2 \localbus/I_18  ( .A(\localbus/N254 ), .ZN(\localbus/N255 ) );
  INV_X2 \localbus/I_19  ( .A(\localbus/c1_op[OP][1] ), .ZN(\localbus/N256 )
         );
  OR2_X2 \localbus/C796  ( .A1(\localbus/c1_op[OP][0] ), .A2(\localbus/N256 ), 
        .ZN(\localbus/N257 ) );
  INV_X2 \localbus/I_20  ( .A(\localbus/N257 ), .ZN(\localbus/N258 ) );
  OR2_X2 \localbus/C799  ( .A1(\localbus/c1_op[SLAVE][0] ), .A2(
        \localbus/N227 ), .ZN(\localbus/N260 ) );
  INV_X2 \localbus/I_21  ( .A(\localbus/N260 ), .ZN(\localbus/N261 ) );
  OR2_X2 \localbus/C802  ( .A1(\localbus/N250 ), .A2(\localbus/c1_op[OP][1] ), 
        .ZN(\localbus/N262 ) );
  INV_X2 \localbus/I_22  ( .A(\localbus/N262 ), .ZN(\localbus/N263 ) );
  OR2_X2 \localbus/C806  ( .A1(n6637), .A2(\localbus/N227 ), .ZN(
        \localbus/N265 ) );
  INV_X2 \localbus/I_23  ( .A(\localbus/N265 ), .ZN(\localbus/N266 ) );
  OR2_X2 \localbus/C809  ( .A1(\localbus/c1_op[OP][0] ), .A2(\localbus/N256 ), 
        .ZN(\localbus/N267 ) );
  INV_X2 \localbus/I_24  ( .A(\localbus/N267 ), .ZN(\localbus/N268 ) );
  OR2_X2 \localbus/C813  ( .A1(n6637), .A2(\localbus/N227 ), .ZN(
        \localbus/N270 ) );
  INV_X2 \localbus/I_25  ( .A(\localbus/N270 ), .ZN(\localbus/N271 ) );
  OR2_X2 \localbus/C850  ( .A1(\localbus/c1_op[OP][0] ), .A2(\localbus/N256 ), 
        .ZN(\localbus/N296 ) );
  INV_X2 \localbus/I_37  ( .A(\localbus/N296 ), .ZN(\localbus/N297 ) );
  OR2_X2 \localbus/C881  ( .A1(\localbus/c2_op[SLAVE][1] ), .A2(
        \localbus/c2_op[SLAVE][2] ), .ZN(\localbus/N318 ) );
  OR2_X2 \localbus/C882  ( .A1(\localbus/N219 ), .A2(\localbus/N318 ), .ZN(
        \localbus/N319 ) );
  INV_X2 \localbus/I_46  ( .A(\localbus/N319 ), .ZN(\localbus/N320 ) );
  OR2_X2 \localbus/C885  ( .A1(\localbus/N293 ), .A2(\localbus/c2_op[OP][1] ), 
        .ZN(\localbus/N321 ) );
  INV_X2 \localbus/I_47  ( .A(\localbus/N321 ), .ZN(\localbus/N322 ) );
  OR2_X2 \localbus/C888  ( .A1(\localbus/c2_op[SLAVE][1] ), .A2(
        \localbus/c2_op[SLAVE][2] ), .ZN(\localbus/N323 ) );
  OR2_X2 \localbus/C889  ( .A1(\localbus/N219 ), .A2(\localbus/N323 ), .ZN(
        \localbus/N324 ) );
  INV_X2 \localbus/I_48  ( .A(\localbus/N324 ), .ZN(\localbus/N325 ) );
  OR2_X2 \localbus/C892  ( .A1(\localbus/N293 ), .A2(\localbus/c2_op[OP][1] ), 
        .ZN(\localbus/N326 ) );
  INV_X2 \localbus/I_49  ( .A(\localbus/N326 ), .ZN(\localbus/N327 ) );
  OR2_X2 \localbus/C894  ( .A1(\localbus/c2_op[SLAVE][1] ), .A2(
        \localbus/c2_op[SLAVE][2] ), .ZN(\localbus/N328 ) );
  OR2_X2 \localbus/C895  ( .A1(\localbus/c2_op[SLAVE][0] ), .A2(
        \localbus/N328 ), .ZN(\localbus/N329 ) );
  OR2_X2 \localbus/C898  ( .A1(\localbus/N293 ), .A2(\localbus/c2_op[OP][1] ), 
        .ZN(\localbus/N331 ) );
  OR2_X2 \localbus/C900  ( .A1(\localbus/c2_op[SLAVE][1] ), .A2(
        \localbus/c2_op[SLAVE][2] ), .ZN(\localbus/N333 ) );
  OR2_X2 \localbus/C901  ( .A1(\localbus/c2_op[SLAVE][0] ), .A2(
        \localbus/N333 ), .ZN(\localbus/N334 ) );
  INV_X2 \localbus/I_52  ( .A(\localbus/N334 ), .ZN(\localbus/N335 ) );
  OR2_X2 \localbus/C904  ( .A1(\localbus/N293 ), .A2(\localbus/c2_op[OP][1] ), 
        .ZN(\localbus/N336 ) );
  INV_X2 \localbus/I_53  ( .A(\localbus/N336 ), .ZN(\localbus/N337 ) );
  OR2_X2 \localbus/C906  ( .A1(\localbus/c1_op[OP][0] ), .A2(
        \localbus/c1_op[OP][1] ), .ZN(\localbus/N338 ) );
  INV_X2 \localbus/I_55  ( .A(dmem_read), .ZN(\localbus/c1_op[OP][0] ) );
  INV_X2 \localbus/I_56  ( .A(dmem_write), .ZN(\localbus/N46 ) );
  AND2_X2 \localbus/C959  ( .A1(\localbus/N50 ), .A2(\localbus/N297 ), .ZN(
        \localbus/N51 ) );
  AND2_X2 \localbus/C964  ( .A1(\localbus/N55 ), .A2(\localbus/N56 ), .ZN(
        \localbus/N57 ) );
  AND2_X2 \localbus/C967  ( .A1(\localbus/N60 ), .A2(\localbus/N61 ), .ZN(
        \localbus/N62 ) );
  AND2_X2 \localbus/C983  ( .A1(\localbus/N252 ), .A2(\localbus/N255 ), .ZN(
        \localbus/N85 ) );
  AND2_X2 \localbus/C984  ( .A1(\localbus/N263 ), .A2(\localbus/N266 ), .ZN(
        \localbus/N86 ) );
  AND2_X2 \localbus/C987  ( .A1(\localbus/N258 ), .A2(\localbus/N261 ), .ZN(
        \localbus/N89 ) );
  AND2_X2 \localbus/C988  ( .A1(\localbus/N268 ), .A2(\localbus/N271 ), .ZN(
        \localbus/N90 ) );
  AND2_X2 \localbus/C993  ( .A1(\localbus/N325 ), .A2(\localbus/N327 ), .ZN(
        \localbus/N95 ) );
  AND2_X2 \localbus/C1001  ( .A1(\localbus/N320 ), .A2(\localbus/N322 ), .ZN(
        \localbus/N199 ) );
  INV_X2 \UUT/Mpath/the_memhandle/I_0  ( .A(dmem_isbyte), .ZN(
        \UUT/Mpath/the_memhandle/N234 ) );
  INV_X2 \UUT/Mpath/the_memhandle/I_3  ( .A(dmem_ishalf), .ZN(
        \UUT/Mpath/the_memhandle/N237 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C342  ( .A1(\UUT/Mpath/the_memhandle/N235 ), 
        .A2(\UUT/Mpath/the_memhandle/N236 ), .ZN(\UUT/Mpath/the_memhandle/N34 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C344  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N36 ) );
  INV_X2 \UUT/Mpath/the_memhandle/I_8  ( .A(\UUT/Mpath/the_memhandle/N241 ), 
        .ZN(\UUT/Mpath/the_memhandle/N37 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C348  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N241 )
         );
  INV_X2 \UUT/Mpath/the_memhandle/I_9  ( .A(\UUT/Mpath/the_memhandle/N242 ), 
        .ZN(\UUT/Mpath/the_memhandle/N38 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C351  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N242 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C353  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N39 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C354  ( .A1(\UUT/m_mem_command[SIGN] ), 
        .A2(\UUT/Mpath/the_memhandle/N236 ), .ZN(\UUT/Mpath/the_memhandle/N72 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C356  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N74 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C360  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N243 )
         );
  INV_X2 \UUT/Mpath/the_memhandle/I_12  ( .A(\UUT/Mpath/the_memhandle/N244 ), 
        .ZN(\UUT/Mpath/the_memhandle/N76 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C363  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N244 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C365  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N77 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C366  ( .A1(\UUT/Mpath/the_memhandle/N235 ), 
        .A2(\UUT/Mpath/the_memhandle/N238 ), .ZN(\UUT/Mpath/the_memhandle/N86 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C369  ( .A1(\UUT/m_mem_command[SIGN] ), 
        .A2(\UUT/Mpath/the_memhandle/N238 ), .ZN(
        \UUT/Mpath/the_memhandle/N120 ) );
  OR2_X2 \UUT/Mpath/the_mult/C331  ( .A1(\UUT/Mpath/the_mult/x_mul_command[4] ), .A2(\UUT/Mpath/the_mult/x_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N194 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C332  ( .A1(\UUT/Mpath/the_mult/N192 ), .A2(
        \UUT/Mpath/the_mult/N194 ), .ZN(\UUT/Mpath/the_mult/N195 ) );
  OR2_X2 \UUT/Mpath/the_mult/C333  ( .A1(\UUT/Mpath/the_mult/x_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N195 ), .ZN(\UUT/Mpath/the_mult/N196 ) );
  OR2_X2 \UUT/Mpath/the_mult/C334  ( .A1(\UUT/Mpath/the_mult/x_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N196 ), .ZN(\UUT/Mpath/the_mult/N197 ) );
  OR2_X2 \UUT/Mpath/the_mult/C335  ( .A1(\UUT/Mpath/the_mult/N193 ), .A2(
        \UUT/Mpath/the_mult/N197 ), .ZN(\UUT/Mpath/the_mult/N198 ) );
  OR2_X2 \UUT/Mpath/the_mult/C353  ( .A1(\UUT/Mpath/the_mult/x_mul_command[4] ), .A2(\UUT/Mpath/the_mult/x_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N212 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C354  ( .A1(\UUT/Mpath/the_mult/N192 ), .A2(
        \UUT/Mpath/the_mult/N212 ), .ZN(\UUT/Mpath/the_mult/N213 ) );
  OR2_X2 \UUT/Mpath/the_mult/C355  ( .A1(\UUT/Mpath/the_mult/x_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N213 ), .ZN(\UUT/Mpath/the_mult/N214 ) );
  OR2_X2 \UUT/Mpath/the_mult/C356  ( .A1(\UUT/Mpath/the_mult/x_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N214 ), .ZN(\UUT/Mpath/the_mult/N215 ) );
  INV_X2 \UUT/Mpath/the_mult/I_8  ( .A(\UUT/d_mul_command [3]), .ZN(
        \UUT/Mpath/the_mult/N220 ) );
  INV_X2 \UUT/Mpath/the_mult/I_9  ( .A(\UUT/d_mul_command [2]), .ZN(
        \UUT/Mpath/the_mult/N221 ) );
  INV_X2 \UUT/Mpath/the_mult/I_10  ( .A(\UUT/d_mul_command [1]), .ZN(
        \UUT/Mpath/the_mult/N222 ) );
  INV_X2 \UUT/Mpath/the_mult/I_11  ( .A(\UUT/d_mul_command [0]), .ZN(
        \UUT/Mpath/the_mult/N223 ) );
  OR2_X2 \UUT/Mpath/the_mult/C370  ( .A1(\UUT/d_mul_command [4]), .A2(
        \UUT/d_mul_command [5]), .ZN(\UUT/Mpath/the_mult/N224 ) );
  OR2_X2 \UUT/Mpath/the_mult/C371  ( .A1(\UUT/Mpath/the_mult/N220 ), .A2(
        \UUT/Mpath/the_mult/N224 ), .ZN(\UUT/Mpath/the_mult/N225 ) );
  OR2_X2 \UUT/Mpath/the_mult/C372  ( .A1(\UUT/Mpath/the_mult/N221 ), .A2(
        \UUT/Mpath/the_mult/N225 ), .ZN(\UUT/Mpath/the_mult/N226 ) );
  OR2_X2 \UUT/Mpath/the_mult/C373  ( .A1(\UUT/Mpath/the_mult/N222 ), .A2(
        \UUT/Mpath/the_mult/N226 ), .ZN(\UUT/Mpath/the_mult/N227 ) );
  OR2_X2 \UUT/Mpath/the_mult/C404  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N251 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C405  ( .A1(\UUT/Mpath/the_mult/N229 ), .A2(
        \UUT/Mpath/the_mult/N251 ), .ZN(\UUT/Mpath/the_mult/N252 ) );
  OR2_X2 \UUT/Mpath/the_mult/C406  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N252 ), .ZN(\UUT/Mpath/the_mult/N253 ) );
  OR2_X2 \UUT/Mpath/the_mult/C407  ( .A1(\UUT/Mpath/the_mult/N230 ), .A2(
        \UUT/Mpath/the_mult/N253 ), .ZN(\UUT/Mpath/the_mult/N254 ) );
  OR2_X2 \UUT/Mpath/the_mult/C408  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N254 ), .ZN(\UUT/Mpath/the_mult/N255 ) );
  OR2_X2 \UUT/Mpath/the_mult/C410  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N257 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C411  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N257 ), .ZN(\UUT/Mpath/the_mult/N258 ) );
  OR2_X2 \UUT/Mpath/the_mult/C412  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N258 ), .ZN(\UUT/Mpath/the_mult/N259 ) );
  OR2_X2 \UUT/Mpath/the_mult/C413  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N259 ), .ZN(\UUT/Mpath/the_mult/N260 ) );
  OR2_X2 \UUT/Mpath/the_mult/C414  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N260 ), .ZN(\UUT/Mpath/the_mult/N261 ) );
  INV_X2 \UUT/Mpath/the_mult/I_21  ( .A(\UUT/Mpath/the_mult/N261 ), .ZN(
        \UUT/Mpath/the_mult/N262 ) );
  OR2_X2 \UUT/Mpath/the_mult/C417  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N263 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C418  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N263 ), .ZN(\UUT/Mpath/the_mult/N264 ) );
  OR2_X2 \UUT/Mpath/the_mult/C419  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N264 ), .ZN(\UUT/Mpath/the_mult/N265 ) );
  OR2_X2 \UUT/Mpath/the_mult/C420  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N265 ), .ZN(\UUT/Mpath/the_mult/N266 ) );
  OR2_X2 \UUT/Mpath/the_mult/C421  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N266 ), .ZN(\UUT/Mpath/the_mult/N267 ) );
  INV_X2 \UUT/Mpath/the_mult/I_22  ( .A(\UUT/Mpath/the_mult/N267 ), .ZN(
        \UUT/Mpath/the_mult/N268 ) );
  OR2_X2 \UUT/Mpath/the_mult/C424  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N269 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C425  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N269 ), .ZN(\UUT/Mpath/the_mult/N270 ) );
  OR2_X2 \UUT/Mpath/the_mult/C426  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N270 ), .ZN(\UUT/Mpath/the_mult/N271 ) );
  OR2_X2 \UUT/Mpath/the_mult/C427  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N271 ), .ZN(\UUT/Mpath/the_mult/N272 ) );
  OR2_X2 \UUT/Mpath/the_mult/C428  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N272 ), .ZN(\UUT/Mpath/the_mult/N273 ) );
  INV_X2 \UUT/Mpath/the_mult/I_23  ( .A(\UUT/Mpath/the_mult/N273 ), .ZN(
        \UUT/Mpath/the_mult/N274 ) );
  OR2_X2 \UUT/Mpath/the_mult/C432  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N275 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C433  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N275 ), .ZN(\UUT/Mpath/the_mult/N276 ) );
  OR2_X2 \UUT/Mpath/the_mult/C434  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N276 ), .ZN(\UUT/Mpath/the_mult/N277 ) );
  OR2_X2 \UUT/Mpath/the_mult/C435  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N277 ), .ZN(\UUT/Mpath/the_mult/N278 ) );
  OR2_X2 \UUT/Mpath/the_mult/C436  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N278 ), .ZN(\UUT/Mpath/the_mult/N279 ) );
  INV_X2 \UUT/Mpath/the_mult/I_24  ( .A(\UUT/Mpath/the_mult/N279 ), .ZN(
        \UUT/Mpath/the_mult/N280 ) );
  OR2_X2 \UUT/Mpath/the_mult/C440  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N281 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C441  ( .A1(\UUT/Mpath/the_mult/N229 ), .A2(
        \UUT/Mpath/the_mult/N281 ), .ZN(\UUT/Mpath/the_mult/N282 ) );
  OR2_X2 \UUT/Mpath/the_mult/C442  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N282 ), .ZN(\UUT/Mpath/the_mult/N283 ) );
  OR2_X2 \UUT/Mpath/the_mult/C443  ( .A1(\UUT/Mpath/the_mult/N230 ), .A2(
        \UUT/Mpath/the_mult/N283 ), .ZN(\UUT/Mpath/the_mult/N284 ) );
  OR2_X2 \UUT/Mpath/the_mult/C444  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N284 ), .ZN(\UUT/Mpath/the_mult/N285 ) );
  OR2_X2 \UUT/Mpath/the_mult/C446  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N287 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C447  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N287 ), .ZN(\UUT/Mpath/the_mult/N288 ) );
  OR2_X2 \UUT/Mpath/the_mult/C448  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N288 ), .ZN(\UUT/Mpath/the_mult/N289 ) );
  OR2_X2 \UUT/Mpath/the_mult/C449  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N289 ), .ZN(\UUT/Mpath/the_mult/N290 ) );
  OR2_X2 \UUT/Mpath/the_mult/C450  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N290 ), .ZN(\UUT/Mpath/the_mult/N291 ) );
  INV_X2 \UUT/Mpath/the_mult/I_26  ( .A(\UUT/Mpath/the_mult/N291 ), .ZN(
        \UUT/Mpath/the_mult/N292 ) );
  OR2_X2 \UUT/Mpath/the_mult/C453  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N293 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C454  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N293 ), .ZN(\UUT/Mpath/the_mult/N294 ) );
  OR2_X2 \UUT/Mpath/the_mult/C455  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N294 ), .ZN(\UUT/Mpath/the_mult/N295 ) );
  OR2_X2 \UUT/Mpath/the_mult/C456  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N295 ), .ZN(\UUT/Mpath/the_mult/N296 ) );
  OR2_X2 \UUT/Mpath/the_mult/C457  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N296 ), .ZN(\UUT/Mpath/the_mult/N297 ) );
  INV_X2 \UUT/Mpath/the_mult/I_27  ( .A(\UUT/Mpath/the_mult/N297 ), .ZN(
        \UUT/Mpath/the_mult/N298 ) );
  OR2_X2 \UUT/Mpath/the_mult/C496  ( .A1(\UUT/Mpath/the_mult/N262 ), .A2(
        \UUT/Mpath/the_mult/N268 ), .ZN(\UUT/Mpath/the_mult/N311 ) );
  OR2_X2 \UUT/Mpath/the_mult/C499  ( .A1(\UUT/Mpath/the_mult/N274 ), .A2(
        \UUT/Mpath/the_mult/N280 ), .ZN(\UUT/Mpath/the_mult/N312 ) );
  OR2_X2 \UUT/Mpath/the_mult/C504  ( .A1(\UUT/Mpath/the_mult/N292 ), .A2(
        \UUT/Mpath/the_mult/N298 ), .ZN(\UUT/Mpath/the_mult/N313 ) );
  OR2_X2 \UUT/Mpath/the_shift/C151  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/Mpath/the_shift/N104 ), .ZN(\UUT/Mpath/the_shift/N106 ) );
  OR2_X2 \UUT/Mpath/the_shift/C152  ( .A1(\UUT/Mpath/the_shift/N105 ), .A2(
        \UUT/Mpath/the_shift/N106 ), .ZN(\UUT/Mpath/the_shift/N107 ) );
  INV_X2 \UUT/Mpath/the_shift/I_2  ( .A(\UUT/Mpath/the_shift/N107 ), .ZN(
        \UUT/Mpath/the_shift/N108 ) );
  OR2_X2 \UUT/Mpath/the_shift/C155  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/Mpath/the_shift/N104 ), .ZN(\UUT/Mpath/the_shift/N109 ) );
  OR2_X2 \UUT/Mpath/the_shift/C156  ( .A1(\UUT/shift_op [0]), .A2(
        \UUT/Mpath/the_shift/N109 ), .ZN(\UUT/Mpath/the_shift/N110 ) );
  INV_X2 \UUT/Mpath/the_shift/I_3  ( .A(\UUT/Mpath/the_shift/N110 ), .ZN(
        \UUT/Mpath/the_shift/N111 ) );
  OR2_X2 \UUT/Mpath/the_shift/C159  ( .A1(\UUT/Mpath/the_shift/N112 ), .A2(
        \UUT/shift_op [2]), .ZN(\UUT/Mpath/the_shift/N113 ) );
  OR2_X2 \UUT/Mpath/the_shift/C160  ( .A1(\UUT/shift_op [0]), .A2(
        \UUT/Mpath/the_shift/N113 ), .ZN(\UUT/Mpath/the_shift/N114 ) );
  INV_X2 \UUT/Mpath/the_shift/I_5  ( .A(\UUT/Mpath/the_shift/N114 ), .ZN(
        \UUT/Mpath/the_shift/N115 ) );
  OR2_X2 \UUT/Mpath/the_shift/C163  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/shift_op [2]), .ZN(\UUT/Mpath/the_shift/N116 ) );
  OR2_X2 \UUT/Mpath/the_shift/C164  ( .A1(\UUT/Mpath/the_shift/N105 ), .A2(
        \UUT/Mpath/the_shift/N116 ), .ZN(\UUT/Mpath/the_shift/N117 ) );
  INV_X2 \UUT/Mpath/the_shift/I_6  ( .A(\UUT/Mpath/the_shift/N117 ), .ZN(
        \UUT/Mpath/the_shift/N118 ) );
  OR2_X2 \UUT/Mpath/the_alu/C476  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N469 ) );
  OR2_X2 \UUT/Mpath/the_alu/C477  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N469 ), .ZN(\UUT/Mpath/the_alu/N470 ) );
  OR2_X2 \UUT/Mpath/the_alu/C478  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N470 ), .ZN(\UUT/Mpath/the_alu/N471 ) );
  OR2_X2 \UUT/Mpath/the_alu/C479  ( .A1(\UUT/Mpath/the_alu/N467 ), .A2(
        \UUT/Mpath/the_alu/N471 ), .ZN(\UUT/Mpath/the_alu/N472 ) );
  OR2_X2 \UUT/Mpath/the_alu/C480  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N472 ), .ZN(\UUT/Mpath/the_alu/N473 ) );
  INV_X2 \UUT/Mpath/the_alu/I_9  ( .A(\UUT/Mpath/the_alu/N473 ), .ZN(
        \UUT/Mpath/the_alu/N474 ) );
  OR2_X2 \UUT/Mpath/the_alu/C485  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N475 ) );
  OR2_X2 \UUT/Mpath/the_alu/C486  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N475 ), .ZN(\UUT/Mpath/the_alu/N476 ) );
  OR2_X2 \UUT/Mpath/the_alu/C487  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N476 ), .ZN(\UUT/Mpath/the_alu/N477 ) );
  OR2_X2 \UUT/Mpath/the_alu/C488  ( .A1(\UUT/Mpath/the_alu/N467 ), .A2(
        \UUT/Mpath/the_alu/N477 ), .ZN(\UUT/Mpath/the_alu/N478 ) );
  OR2_X2 \UUT/Mpath/the_alu/C489  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N478 ), .ZN(\UUT/Mpath/the_alu/N479 ) );
  INV_X2 \UUT/Mpath/the_alu/I_10  ( .A(\UUT/Mpath/the_alu/N479 ), .ZN(
        \UUT/Mpath/the_alu/N480 ) );
  OR2_X2 \UUT/Mpath/the_alu/C494  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N481 ) );
  OR2_X2 \UUT/Mpath/the_alu/C495  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N481 ), .ZN(\UUT/Mpath/the_alu/N482 ) );
  OR2_X2 \UUT/Mpath/the_alu/C496  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N482 ), .ZN(\UUT/Mpath/the_alu/N483 ) );
  OR2_X2 \UUT/Mpath/the_alu/C497  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N483 ), .ZN(\UUT/Mpath/the_alu/N484 ) );
  OR2_X2 \UUT/Mpath/the_alu/C498  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N484 ), .ZN(\UUT/Mpath/the_alu/N485 ) );
  INV_X2 \UUT/Mpath/the_alu/I_11  ( .A(\UUT/Mpath/the_alu/N485 ), .ZN(
        \UUT/Mpath/the_alu/N486 ) );
  OR2_X2 \UUT/Mpath/the_alu/C502  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N487 ) );
  OR2_X2 \UUT/Mpath/the_alu/C503  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N487 ), .ZN(\UUT/Mpath/the_alu/N488 ) );
  OR2_X2 \UUT/Mpath/the_alu/C504  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N488 ), .ZN(\UUT/Mpath/the_alu/N489 ) );
  OR2_X2 \UUT/Mpath/the_alu/C505  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N489 ), .ZN(\UUT/Mpath/the_alu/N490 ) );
  OR2_X2 \UUT/Mpath/the_alu/C506  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N490 ), .ZN(\UUT/Mpath/the_alu/N491 ) );
  OR2_X2 \UUT/Mpath/the_alu/C510  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N493 ) );
  OR2_X2 \UUT/Mpath/the_alu/C511  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N493 ), .ZN(\UUT/Mpath/the_alu/N494 ) );
  OR2_X2 \UUT/Mpath/the_alu/C512  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N494 ), .ZN(\UUT/Mpath/the_alu/N495 ) );
  OR2_X2 \UUT/Mpath/the_alu/C513  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N495 ), .ZN(\UUT/Mpath/the_alu/N496 ) );
  OR2_X2 \UUT/Mpath/the_alu/C514  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N496 ), .ZN(\UUT/Mpath/the_alu/N497 ) );
  INV_X2 \UUT/Mpath/the_alu/I_13  ( .A(\UUT/Mpath/the_alu/N497 ), .ZN(
        \UUT/Mpath/the_alu/N498 ) );
  OR2_X2 \UUT/Mpath/the_alu/C517  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N499 ) );
  OR2_X2 \UUT/Mpath/the_alu/C518  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N499 ), .ZN(\UUT/Mpath/the_alu/N500 ) );
  OR2_X2 \UUT/Mpath/the_alu/C519  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N500 ), .ZN(\UUT/Mpath/the_alu/N501 ) );
  OR2_X2 \UUT/Mpath/the_alu/C520  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N501 ), .ZN(\UUT/Mpath/the_alu/N502 ) );
  OR2_X2 \UUT/Mpath/the_alu/C521  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N502 ), .ZN(\UUT/Mpath/the_alu/N503 ) );
  OR2_X2 \UUT/Mpath/the_alu/C524  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Alu_command[OP][5] ), .ZN(\UUT/Mpath/the_alu/N505 ) );
  OR2_X2 \UUT/Mpath/the_alu/C525  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N505 ), .ZN(\UUT/Mpath/the_alu/N506 ) );
  OR2_X2 \UUT/Mpath/the_alu/C526  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N506 ), .ZN(\UUT/Mpath/the_alu/N507 ) );
  OR2_X2 \UUT/Mpath/the_alu/C527  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N507 ), .ZN(\UUT/Mpath/the_alu/N508 ) );
  OR2_X2 \UUT/Mpath/the_alu/C528  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N508 ), .ZN(\UUT/Mpath/the_alu/N509 ) );
  OR2_X2 \UUT/Mpath/the_alu/C532  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Alu_command[OP][5] ), .ZN(\UUT/Mpath/the_alu/N511 ) );
  OR2_X2 \UUT/Mpath/the_alu/C533  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N511 ), .ZN(\UUT/Mpath/the_alu/N512 ) );
  OR2_X2 \UUT/Mpath/the_alu/C534  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N512 ), .ZN(\UUT/Mpath/the_alu/N513 ) );
  OR2_X2 \UUT/Mpath/the_alu/C535  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N513 ), .ZN(\UUT/Mpath/the_alu/N514 ) );
  OR2_X2 \UUT/Mpath/the_alu/C536  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N514 ), .ZN(\UUT/Mpath/the_alu/N515 ) );
  OR2_X2 \UUT/Mpath/the_alu/C538  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Alu_command[OP][5] ), .ZN(\UUT/Mpath/the_alu/N517 ) );
  OR2_X2 \UUT/Mpath/the_alu/C539  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N517 ), .ZN(\UUT/Mpath/the_alu/N518 ) );
  OR2_X2 \UUT/Mpath/the_alu/C540  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N518 ), .ZN(\UUT/Mpath/the_alu/N519 ) );
  OR2_X2 \UUT/Mpath/the_alu/C541  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N519 ), .ZN(\UUT/Mpath/the_alu/N520 ) );
  OR2_X2 \UUT/Mpath/the_alu/C545  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Alu_command[OP][5] ), .ZN(\UUT/Mpath/the_alu/N523 ) );
  OR2_X2 \UUT/Mpath/the_alu/C546  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N523 ), .ZN(\UUT/Mpath/the_alu/N524 ) );
  OR2_X2 \UUT/Mpath/the_alu/C547  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N524 ), .ZN(\UUT/Mpath/the_alu/N525 ) );
  OR2_X2 \UUT/Mpath/the_alu/C548  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N525 ), .ZN(\UUT/Mpath/the_alu/N526 ) );
  AND2_X2 \UUT/Mpath/the_alu/C575  ( .A1(\UUT/Mpath/out_regA[31] ), .A2(
        \UUT/Mpath/out_regB[31] ), .ZN(\UUT/Mpath/the_alu/N94 ) );
  OR2_X2 \UUT/Mpath/the_alu/C608  ( .A1(\UUT/Mpath/out_regA[31] ), .A2(
        \UUT/Mpath/out_regB[31] ), .ZN(\UUT/Mpath/the_alu/N126 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C641  ( .A(\UUT/Mpath/out_regA[31] ), .B(
        \UUT/Mpath/out_regB[31] ), .Z(\UUT/Mpath/the_alu/N158 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C642  ( .A(\UUT/Mpath/out_regA[30] ), .B(
        \UUT/Mpath/out_regB[30] ), .Z(\UUT/Mpath/the_alu/N159 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C643  ( .A(\UUT/Mpath/out_regA[29] ), .B(
        \UUT/Mpath/out_regB[29] ), .Z(\UUT/Mpath/the_alu/N160 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C644  ( .A(\UUT/Mpath/out_regA[28] ), .B(
        \UUT/Mpath/out_regB[28] ), .Z(\UUT/Mpath/the_alu/N161 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C645  ( .A(\UUT/Mpath/out_regA[27] ), .B(
        \UUT/Mpath/out_regB[27] ), .Z(\UUT/Mpath/the_alu/N162 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C646  ( .A(\UUT/Mpath/out_regA[26] ), .B(
        \UUT/Mpath/out_regB[26] ), .Z(\UUT/Mpath/the_alu/N163 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C647  ( .A(\UUT/Mpath/out_regA[25] ), .B(
        \UUT/Mpath/out_regB[25] ), .Z(\UUT/Mpath/the_alu/N164 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C648  ( .A(\UUT/Mpath/out_regA[24] ), .B(
        \UUT/Mpath/out_regB[24] ), .Z(\UUT/Mpath/the_alu/N165 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C649  ( .A(\UUT/Mpath/out_regA[23] ), .B(
        \UUT/Mpath/out_regB[23] ), .Z(\UUT/Mpath/the_alu/N166 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C650  ( .A(\UUT/Mpath/out_regA[22] ), .B(
        \UUT/Mpath/out_regB[22] ), .Z(\UUT/Mpath/the_alu/N167 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C651  ( .A(\UUT/Mpath/out_regA[21] ), .B(
        \UUT/Mpath/out_regB[21] ), .Z(\UUT/Mpath/the_alu/N168 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C652  ( .A(\UUT/Mpath/out_regA[20] ), .B(
        \UUT/Mpath/out_regB[20] ), .Z(\UUT/Mpath/the_alu/N169 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C653  ( .A(\UUT/Mpath/out_regA[19] ), .B(
        \UUT/Mpath/out_regB[19] ), .Z(\UUT/Mpath/the_alu/N170 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C654  ( .A(\UUT/Mpath/out_regA[18] ), .B(
        \UUT/Mpath/out_regB[18] ), .Z(\UUT/Mpath/the_alu/N171 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C655  ( .A(\UUT/Mpath/out_regA[17] ), .B(
        \UUT/Mpath/out_regB[17] ), .Z(\UUT/Mpath/the_alu/N172 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C656  ( .A(\UUT/Mpath/out_regA[16] ), .B(
        \UUT/Mpath/out_regB[16] ), .Z(\UUT/Mpath/the_alu/N173 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C657  ( .A(\UUT/Mpath/out_regA[15] ), .B(
        \UUT/Mpath/out_regB[15] ), .Z(\UUT/Mpath/the_alu/N174 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C658  ( .A(\UUT/Mpath/out_regA[14] ), .B(
        \UUT/Mpath/out_regB[14] ), .Z(\UUT/Mpath/the_alu/N175 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C659  ( .A(\UUT/Mpath/out_regA[13] ), .B(
        \UUT/Mpath/out_regB[13] ), .Z(\UUT/Mpath/the_alu/N176 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C660  ( .A(\UUT/Mpath/out_regA[12] ), .B(
        \UUT/Mpath/out_regB[12] ), .Z(\UUT/Mpath/the_alu/N177 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C661  ( .A(\UUT/Mpath/out_regA[11] ), .B(
        \UUT/Mpath/out_regB[11] ), .Z(\UUT/Mpath/the_alu/N178 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C662  ( .A(\UUT/Mpath/out_regA[10] ), .B(
        \UUT/Mpath/out_regB[10] ), .Z(\UUT/Mpath/the_alu/N179 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C663  ( .A(\UUT/Mpath/out_regA[9] ), .B(
        \UUT/Mpath/out_regB[9] ), .Z(\UUT/Mpath/the_alu/N180 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C664  ( .A(\UUT/Mpath/out_regA[8] ), .B(
        \UUT/Mpath/out_regB[8] ), .Z(\UUT/Mpath/the_alu/N181 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C665  ( .A(\UUT/Mpath/out_regA[7] ), .B(
        \UUT/Mpath/out_regB[7] ), .Z(\UUT/Mpath/the_alu/N182 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C666  ( .A(\UUT/Mpath/out_regA[6] ), .B(
        \UUT/Mpath/out_regB[6] ), .Z(\UUT/Mpath/the_alu/N183 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C667  ( .A(\UUT/Mpath/out_regA[5] ), .B(
        \UUT/Mpath/out_regB[5] ), .Z(\UUT/Mpath/the_alu/N184 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C668  ( .A(\UUT/Mpath/out_regA[4] ), .B(n6897), 
        .Z(\UUT/Mpath/the_alu/N185 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C669  ( .A(\UUT/Mpath/out_regA[3] ), .B(n6898), 
        .Z(\UUT/Mpath/the_alu/N186 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C670  ( .A(\UUT/Mpath/out_regA[2] ), .B(n6899), 
        .Z(\UUT/Mpath/the_alu/N187 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C672  ( .A(n6525), .B(n6675), .Z(
        \UUT/Mpath/the_alu/N189 ) );
  AND2_X2 \UUT/Mpath/the_alu/C674  ( .A1(\UUT/Mpath/the_alu/N21 ), .A2(
        \UUT/Mpath/the_alu/N22 ), .ZN(\UUT/Mpath/the_alu/N190 ) );
  AND2_X2 \UUT/Mpath/the_alu/C675  ( .A1(\UUT/Mpath/the_alu/N23 ), .A2(
        \UUT/Mpath/the_alu/N24 ), .ZN(\UUT/Mpath/the_alu/N191 ) );
  AND2_X2 \UUT/Mpath/the_alu/C676  ( .A1(\UUT/Mpath/the_alu/N25 ), .A2(
        \UUT/Mpath/the_alu/N26 ), .ZN(\UUT/Mpath/the_alu/N192 ) );
  AND2_X2 \UUT/Mpath/the_alu/C677  ( .A1(\UUT/Mpath/the_alu/N27 ), .A2(
        \UUT/Mpath/the_alu/N28 ), .ZN(\UUT/Mpath/the_alu/N193 ) );
  AND2_X2 \UUT/Mpath/the_alu/C678  ( .A1(\UUT/Mpath/the_alu/N29 ), .A2(
        \UUT/Mpath/the_alu/N30 ), .ZN(\UUT/Mpath/the_alu/N194 ) );
  AND2_X2 \UUT/Mpath/the_alu/C679  ( .A1(\UUT/Mpath/the_alu/N31 ), .A2(
        \UUT/Mpath/the_alu/N32 ), .ZN(\UUT/Mpath/the_alu/N195 ) );
  AND2_X2 \UUT/Mpath/the_alu/C680  ( .A1(\UUT/Mpath/the_alu/N33 ), .A2(
        \UUT/Mpath/the_alu/N34 ), .ZN(\UUT/Mpath/the_alu/N196 ) );
  AND2_X2 \UUT/Mpath/the_alu/C681  ( .A1(\UUT/Mpath/the_alu/N35 ), .A2(
        \UUT/Mpath/the_alu/N36 ), .ZN(\UUT/Mpath/the_alu/N197 ) );
  AND2_X2 \UUT/Mpath/the_alu/C682  ( .A1(\UUT/Mpath/the_alu/N37 ), .A2(
        \UUT/Mpath/the_alu/N38 ), .ZN(\UUT/Mpath/the_alu/N198 ) );
  AND2_X2 \UUT/Mpath/the_alu/C683  ( .A1(\UUT/Mpath/the_alu/N39 ), .A2(
        \UUT/Mpath/the_alu/N40 ), .ZN(\UUT/Mpath/the_alu/N199 ) );
  AND2_X2 \UUT/Mpath/the_alu/C684  ( .A1(\UUT/Mpath/the_alu/N41 ), .A2(
        \UUT/Mpath/the_alu/N42 ), .ZN(\UUT/Mpath/the_alu/N200 ) );
  AND2_X2 \UUT/Mpath/the_alu/C685  ( .A1(\UUT/Mpath/the_alu/N43 ), .A2(
        \UUT/Mpath/the_alu/N44 ), .ZN(\UUT/Mpath/the_alu/N201 ) );
  AND2_X2 \UUT/Mpath/the_alu/C686  ( .A1(\UUT/Mpath/the_alu/N45 ), .A2(
        \UUT/Mpath/the_alu/N46 ), .ZN(\UUT/Mpath/the_alu/N202 ) );
  AND2_X2 \UUT/Mpath/the_alu/C687  ( .A1(\UUT/Mpath/the_alu/N47 ), .A2(
        \UUT/Mpath/the_alu/N48 ), .ZN(\UUT/Mpath/the_alu/N203 ) );
  AND2_X2 \UUT/Mpath/the_alu/C688  ( .A1(\UUT/Mpath/the_alu/N49 ), .A2(
        \UUT/Mpath/the_alu/N50 ), .ZN(\UUT/Mpath/the_alu/N204 ) );
  AND2_X2 \UUT/Mpath/the_alu/C689  ( .A1(\UUT/Mpath/the_alu/N51 ), .A2(
        \UUT/Mpath/the_alu/N52 ), .ZN(\UUT/Mpath/the_alu/N205 ) );
  AND2_X2 \UUT/Mpath/the_alu/C690  ( .A1(\UUT/Mpath/the_alu/N53 ), .A2(
        \UUT/Mpath/the_alu/N54 ), .ZN(\UUT/Mpath/the_alu/N206 ) );
  AND2_X2 \UUT/Mpath/the_alu/C691  ( .A1(\UUT/Mpath/the_alu/N55 ), .A2(
        \UUT/Mpath/the_alu/N56 ), .ZN(\UUT/Mpath/the_alu/N207 ) );
  AND2_X2 \UUT/Mpath/the_alu/C692  ( .A1(\UUT/Mpath/the_alu/N57 ), .A2(
        \UUT/Mpath/the_alu/N58 ), .ZN(\UUT/Mpath/the_alu/N208 ) );
  AND2_X2 \UUT/Mpath/the_alu/C693  ( .A1(\UUT/Mpath/the_alu/N59 ), .A2(
        \UUT/Mpath/the_alu/N60 ), .ZN(\UUT/Mpath/the_alu/N209 ) );
  AND2_X2 \UUT/Mpath/the_alu/C694  ( .A1(\UUT/Mpath/the_alu/N61 ), .A2(
        \UUT/Mpath/the_alu/N62 ), .ZN(\UUT/Mpath/the_alu/N210 ) );
  AND2_X2 \UUT/Mpath/the_alu/C695  ( .A1(\UUT/Mpath/the_alu/N63 ), .A2(
        \UUT/Mpath/the_alu/N64 ), .ZN(\UUT/Mpath/the_alu/N211 ) );
  AND2_X2 \UUT/Mpath/the_alu/C696  ( .A1(\UUT/Mpath/the_alu/N65 ), .A2(
        \UUT/Mpath/the_alu/N66 ), .ZN(\UUT/Mpath/the_alu/N212 ) );
  AND2_X2 \UUT/Mpath/the_alu/C697  ( .A1(\UUT/Mpath/the_alu/N67 ), .A2(
        \UUT/Mpath/the_alu/N68 ), .ZN(\UUT/Mpath/the_alu/N213 ) );
  AND2_X2 \UUT/Mpath/the_alu/C698  ( .A1(\UUT/Mpath/the_alu/N69 ), .A2(
        \UUT/Mpath/the_alu/N70 ), .ZN(\UUT/Mpath/the_alu/N214 ) );
  AND2_X2 \UUT/Mpath/the_alu/C699  ( .A1(\UUT/Mpath/the_alu/N71 ), .A2(
        \UUT/Mpath/the_alu/N72 ), .ZN(\UUT/Mpath/the_alu/N215 ) );
  AND2_X2 \UUT/Mpath/the_alu/C700  ( .A1(\UUT/Mpath/the_alu/N73 ), .A2(
        \UUT/Mpath/the_alu/N74 ), .ZN(\UUT/Mpath/the_alu/N216 ) );
  AND2_X2 \UUT/Mpath/the_alu/C701  ( .A1(\UUT/Mpath/the_alu/N75 ), .A2(
        \UUT/Mpath/the_alu/N76 ), .ZN(\UUT/Mpath/the_alu/N217 ) );
  AND2_X2 \UUT/Mpath/the_alu/C702  ( .A1(\UUT/Mpath/the_alu/N77 ), .A2(
        \UUT/Mpath/the_alu/N78 ), .ZN(\UUT/Mpath/the_alu/N218 ) );
  AND2_X2 \UUT/Mpath/the_alu/C703  ( .A1(\UUT/Mpath/the_alu/N79 ), .A2(
        \UUT/Mpath/the_alu/N80 ), .ZN(\UUT/Mpath/the_alu/N219 ) );
  AND2_X2 \UUT/Mpath/the_alu/C705  ( .A1(\UUT/Mpath/the_alu/N83 ), .A2(
        \UUT/Mpath/the_alu/N84 ), .ZN(\UUT/Mpath/the_alu/N221 ) );
  OR2_X2 \UUT/Mpath/C262  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/Mpath/N111 ), 
        .ZN(\UUT/Mpath/N113 ) );
  OR2_X2 \UUT/Mpath/C263  ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N113 ), .ZN(
        \UUT/Mpath/N114 ) );
  INV_X2 \UUT/Mpath/I_3  ( .A(\UUT/Mpath/N114 ), .ZN(\UUT/Mpath/N115 ) );
  OR2_X2 \UUT/Mpath/C266  ( .A1(\UUT/Mpath/N116 ), .A2(\UUT/exe_outsel [2]), 
        .ZN(\UUT/Mpath/N117 ) );
  OR2_X2 \UUT/Mpath/C267  ( .A1(\UUT/exe_outsel [0]), .A2(\UUT/Mpath/N117 ), 
        .ZN(\UUT/Mpath/N118 ) );
  INV_X2 \UUT/Mpath/I_5  ( .A(\UUT/Mpath/N118 ), .ZN(\UUT/Mpath/N119 ) );
  OR2_X2 \UUT/Mpath/C275  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/exe_outsel [2]), 
        .ZN(\UUT/Mpath/N124 ) );
  OR2_X2 \UUT/Mpath/C276  ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N124 ), .ZN(
        \UUT/Mpath/N125 ) );
  OR2_X2 \UUT/Mpath/C280  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/Mpath/N111 ), 
        .ZN(\UUT/Mpath/N127 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_0  ( .A(\UUT/Mcontrol/st_logic/load_stall ), 
        .ZN(\UUT/Mcontrol/st_logic/N12 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_1  ( .A(
        \UUT/Mcontrol/st_logic/branchlw_stall ), .ZN(
        \UUT/Mcontrol/st_logic/N13 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_2  ( .A(
        \UUT/Mcontrol/st_logic/branchmul_stall ), .ZN(
        \UUT/Mcontrol/st_logic/N14 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_3  ( .A(dmem_read), .ZN(
        \UUT/Mcontrol/st_logic/N15 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_4  ( .A(\UUT/byp_controlA[2] ), .ZN(
        \UUT/Mcontrol/st_logic/N55 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C75  ( .A1(\UUT/byp_controlA[0] ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N18 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_5  ( .A(\UUT/Mcontrol/st_logic/N18 ), .ZN(
        \UUT/Mcontrol/st_logic/N19 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_6  ( .A(\UUT/byp_controlB[2] ), .ZN(
        \UUT/Mcontrol/st_logic/N52 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C79  ( .A1(\UUT/byp_controlB[0] ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N22 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_7  ( .A(\UUT/Mcontrol/st_logic/N22 ), .ZN(
        \UUT/Mcontrol/st_logic/N23 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_8  ( .A(\UUT/m_mem_command[MR] ), .ZN(
        \UUT/Mcontrol/st_logic/N24 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_9  ( .A(
        \UUT/Mcontrol/st_logic/branch_uses_main_mem_result ), .ZN(
        \UUT/Mcontrol/st_logic/N25 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C85  ( .A1(\UUT/Mcontrol/x_mul_command [4]), 
        .A2(\UUT/Mcontrol/x_mul_command [5]), .ZN(\UUT/Mcontrol/st_logic/N28 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C86  ( .A1(\UUT/Mcontrol/x_mul_command [3]), 
        .A2(\UUT/Mcontrol/st_logic/N28 ), .ZN(\UUT/Mcontrol/st_logic/N29 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C87  ( .A1(\UUT/Mcontrol/st_logic/N26 ), .A2(
        \UUT/Mcontrol/st_logic/N29 ), .ZN(\UUT/Mcontrol/st_logic/N30 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C88  ( .A1(\UUT/Mcontrol/st_logic/N27 ), .A2(
        \UUT/Mcontrol/st_logic/N30 ), .ZN(\UUT/Mcontrol/st_logic/N31 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C89  ( .A1(\UUT/Mcontrol/x_mul_command [0]), 
        .A2(\UUT/Mcontrol/st_logic/N31 ), .ZN(\UUT/Mcontrol/st_logic/N32 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_12  ( .A(\UUT/Mcontrol/st_logic/N32 ), .ZN(
        \UUT/Mcontrol/st_logic/N33 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C94  ( .A1(\UUT/Mcontrol/x_mul_command [4]), 
        .A2(\UUT/Mcontrol/x_mul_command [5]), .ZN(\UUT/Mcontrol/st_logic/N35 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C95  ( .A1(\UUT/Mcontrol/x_mul_command [3]), 
        .A2(\UUT/Mcontrol/st_logic/N35 ), .ZN(\UUT/Mcontrol/st_logic/N36 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C96  ( .A1(\UUT/Mcontrol/st_logic/N26 ), .A2(
        \UUT/Mcontrol/st_logic/N36 ), .ZN(\UUT/Mcontrol/st_logic/N37 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C97  ( .A1(\UUT/Mcontrol/st_logic/N27 ), .A2(
        \UUT/Mcontrol/st_logic/N37 ), .ZN(\UUT/Mcontrol/st_logic/N38 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C98  ( .A1(\UUT/Mcontrol/st_logic/N34 ), .A2(
        \UUT/Mcontrol/st_logic/N38 ), .ZN(\UUT/Mcontrol/st_logic/N39 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_14  ( .A(\UUT/Mcontrol/st_logic/N39 ), .ZN(
        \UUT/Mcontrol/st_logic/N40 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_15  ( .A(
        \UUT/Mcontrol/st_logic/branch_uses_main_exe_result ), .ZN(
        \UUT/Mcontrol/st_logic/N41 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C104  ( .A1(\UUT/Mcontrol/st_logic/N42 ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N44 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_17  ( .A(\UUT/Mcontrol/st_logic/N44 ), .ZN(
        \UUT/Mcontrol/st_logic/N45 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_18  ( .A(
        \UUT/Mcontrol/st_logic/branch_uses_regb ), .ZN(
        \UUT/Mcontrol/st_logic/N46 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C110  ( .A1(\UUT/Mcontrol/st_logic/N47 ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N49 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_20  ( .A(\UUT/Mcontrol/st_logic/N49 ), .ZN(
        \UUT/Mcontrol/st_logic/N50 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_21  ( .A(
        \UUT/Mcontrol/st_logic/branch_uses_rega ), .ZN(
        \UUT/Mcontrol/st_logic/N51 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C115  ( .A1(\UUT/byp_controlB[0] ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N53 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_22  ( .A(\UUT/Mcontrol/st_logic/N53 ), .ZN(
        \UUT/Mcontrol/st_logic/N54 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C120  ( .A1(\UUT/byp_controlA[0] ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N56 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_23  ( .A(\UUT/Mcontrol/st_logic/N56 ), .ZN(
        \UUT/Mcontrol/st_logic/N57 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_24  ( .A(\UUT/Mcontrol/d_jump_type[2] ), 
        .ZN(\UUT/Mcontrol/st_logic/N58 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C126  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N60 ), .ZN(\UUT/Mcontrol/st_logic/N61 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C128  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N62 ), .ZN(\UUT/Mcontrol/st_logic/N63 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_25  ( .A(\UUT/Mcontrol/st_logic/N63 ), .ZN(
        \UUT/Mcontrol/st_logic/N64 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_26  ( .A(\UUT/Mcontrol/d_jump_type[0] ), 
        .ZN(\UUT/Mcontrol/st_logic/N65 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C134  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N67 ), .ZN(\UUT/Mcontrol/st_logic/N68 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C136  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N69 ), .ZN(\UUT/Mcontrol/st_logic/N70 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_27  ( .A(\UUT/Mcontrol/st_logic/N70 ), .ZN(
        \UUT/Mcontrol/st_logic/N71 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C141  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N73 ), .ZN(\UUT/Mcontrol/st_logic/N74 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C143  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N75 ), .ZN(\UUT/Mcontrol/st_logic/N76 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_28  ( .A(\UUT/Mcontrol/st_logic/N76 ), .ZN(
        \UUT/Mcontrol/st_logic/N77 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C149  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N79 ), .ZN(\UUT/Mcontrol/st_logic/N80 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C151  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N81 ), .ZN(\UUT/Mcontrol/st_logic/N82 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_29  ( .A(\UUT/Mcontrol/st_logic/N82 ), .ZN(
        \UUT/Mcontrol/st_logic/N83 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C155  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N85 ), .ZN(\UUT/Mcontrol/st_logic/N86 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C157  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N87 ), .ZN(\UUT/Mcontrol/st_logic/N88 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_30  ( .A(\UUT/Mcontrol/st_logic/N88 ), .ZN(
        \UUT/Mcontrol/st_logic/N89 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C163  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N92 ), .ZN(\UUT/Mcontrol/st_logic/N93 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C164  ( .A1(\UUT/Mcontrol/st_logic/N90 ), .A2(
        \UUT/Mcontrol/st_logic/N93 ), .ZN(\UUT/Mcontrol/st_logic/N94 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C165  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N94 ), .ZN(\UUT/Mcontrol/st_logic/N95 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_32  ( .A(\UUT/Mcontrol/st_logic/N95 ), .ZN(
        \UUT/Mcontrol/st_logic/N96 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C171  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N98 ), .ZN(\UUT/Mcontrol/st_logic/N99 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C172  ( .A1(\UUT/Mcontrol/st_logic/N90 ), .A2(
        \UUT/Mcontrol/st_logic/N99 ), .ZN(\UUT/Mcontrol/st_logic/N100 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C173  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N100 ), .ZN(\UUT/Mcontrol/st_logic/N101 )
         );
  INV_X2 \UUT/Mcontrol/st_logic/I_33  ( .A(\UUT/Mcontrol/st_logic/N101 ), .ZN(
        \UUT/Mcontrol/st_logic/N102 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C179  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N105 ), .ZN(\UUT/Mcontrol/st_logic/N106 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C181  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N107 ), .ZN(\UUT/Mcontrol/st_logic/N108 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_35  ( .A(\UUT/Mcontrol/st_logic/N108 ), .ZN(
        \UUT/Mcontrol/st_logic/N109 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C193  ( .A1(\UUT/Mcontrol/st_logic/N15 ), 
        .A2(\UUT/Mcontrol/st_logic/N110 ), .ZN(\UUT/Mcontrol/st_logic/N2 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C194  ( .A1(\UUT/Mcontrol/st_logic/N19 ), .A2(
        \UUT/Mcontrol/st_logic/N23 ), .ZN(\UUT/Mcontrol/st_logic/N110 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C195  ( .A1(\UUT/Mcontrol/st_logic/N114 ), 
        .A2(\UUT/Mcontrol/st_logic/N109 ), .ZN(\UUT/Mcontrol/st_logic/N3 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C196  ( .A1(\UUT/Mcontrol/st_logic/N113 ), 
        .A2(\UUT/Mcontrol/st_logic/N102 ), .ZN(\UUT/Mcontrol/st_logic/N114 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C197  ( .A1(\UUT/Mcontrol/st_logic/N112 ), 
        .A2(\UUT/Mcontrol/st_logic/N96 ), .ZN(\UUT/Mcontrol/st_logic/N113 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C198  ( .A1(\UUT/Mcontrol/st_logic/N111 ), 
        .A2(\UUT/Mcontrol/st_logic/N89 ), .ZN(\UUT/Mcontrol/st_logic/N112 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C199  ( .A1(\UUT/Mcontrol/st_logic/N77 ), .A2(
        \UUT/Mcontrol/st_logic/N83 ), .ZN(\UUT/Mcontrol/st_logic/N111 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C200  ( .A1(\UUT/Mcontrol/st_logic/N64 ), .A2(
        \UUT/Mcontrol/st_logic/N71 ), .ZN(\UUT/Mcontrol/st_logic/N4 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C201  ( .A1(\UUT/Mcontrol/st_logic/N115 ), 
        .A2(\UUT/Mcontrol/st_logic/N116 ), .ZN(\UUT/Mcontrol/st_logic/N5 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C202  ( .A1(\UUT/Mcontrol/st_logic/N45 ), 
        .A2(\UUT/Mcontrol/st_logic/N46 ), .ZN(\UUT/Mcontrol/st_logic/N115 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C203  ( .A1(\UUT/Mcontrol/st_logic/N50 ), 
        .A2(\UUT/Mcontrol/st_logic/N51 ), .ZN(\UUT/Mcontrol/st_logic/N116 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C204  ( .A1(\UUT/Mcontrol/st_logic/N24 ), 
        .A2(\UUT/Mcontrol/st_logic/N25 ), .ZN(\UUT/Mcontrol/st_logic/N6 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C205  ( .A1(\UUT/Mcontrol/st_logic/N117 ), 
        .A2(\UUT/Mcontrol/st_logic/N118 ), .ZN(\UUT/Mcontrol/st_logic/N7 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C206  ( .A1(\UUT/Mcontrol/st_logic/N54 ), 
        .A2(\UUT/Mcontrol/st_logic/N46 ), .ZN(\UUT/Mcontrol/st_logic/N117 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C207  ( .A1(\UUT/Mcontrol/st_logic/N57 ), 
        .A2(\UUT/Mcontrol/st_logic/N51 ), .ZN(\UUT/Mcontrol/st_logic/N118 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C208  ( .A1(\UUT/Mcontrol/st_logic/N119 ), 
        .A2(\UUT/Mcontrol/st_logic/N41 ), .ZN(\UUT/Mcontrol/st_logic/N8 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C209  ( .A1(\UUT/Mcontrol/st_logic/N33 ), .A2(
        \UUT/Mcontrol/st_logic/N40 ), .ZN(\UUT/Mcontrol/st_logic/N119 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C211  ( .A1(\UUT/Mcontrol/st_logic/N120 ), 
        .A2(\UUT/Mcontrol/st_logic/N14 ), .ZN(\UUT/Mcontrol/st_logic/N10 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C212  ( .A1(\UUT/Mcontrol/st_logic/N12 ), .A2(
        \UUT/Mcontrol/st_logic/N13 ), .ZN(\UUT/Mcontrol/st_logic/N120 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C19  ( .A1(\UUT/Mcontrol/x_rd[3] ), .A2(
        \UUT/Mcontrol/x_rd[4] ), .ZN(\UUT/Mcontrol/bp_logicB/N5 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C20  ( .A1(\UUT/Mcontrol/x_rd[2] ), .A2(
        \UUT/Mcontrol/bp_logicB/N5 ), .ZN(\UUT/Mcontrol/bp_logicB/N6 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C21  ( .A1(\UUT/Mcontrol/x_rd[1] ), .A2(
        \UUT/Mcontrol/bp_logicB/N6 ), .ZN(\UUT/Mcontrol/bp_logicB/N7 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C22  ( .A1(\UUT/Mcontrol/x_rd[0] ), .A2(
        \UUT/Mcontrol/bp_logicB/N7 ), .ZN(\UUT/Mcontrol/bp_logicB/N8 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C26  ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), 
        .A2(\UUT/Mcontrol/m_sampled_xrd[4] ), .ZN(\UUT/Mcontrol/bp_logicB/N10 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C27  ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N10 ), .ZN(\UUT/Mcontrol/bp_logicB/N11 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C28  ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N11 ), .ZN(\UUT/Mcontrol/bp_logicB/N12 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C29  ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N12 ), .ZN(\UUT/Mcontrol/bp_logicB/N13 )
         );
  INV_X2 \UUT/Mcontrol/bp_logicB/I_3  ( .A(\UUT/m_we ), .ZN(
        \UUT/Mcontrol/bp_logicB/N14 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C36  ( .A1(\UUT/Mcontrol/bp_logicB/N15 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N9 ), .ZN(
        \UUT/Mcontrol/bp_logicB/exec_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C37  ( .A1(\UUT/Mcontrol/bp_logicB/N2 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N8 ), .ZN(\UUT/Mcontrol/bp_logicB/N15 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C38  ( .A1(\UUT/Mcontrol/bp_logicB/N16 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N14 ), .ZN(
        \UUT/Mcontrol/bp_logicB/memory_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C39  ( .A1(\UUT/Mcontrol/bp_logicB/N3 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N13 ), .ZN(\UUT/Mcontrol/bp_logicB/N16 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C19  ( .A1(\UUT/Mcontrol/x_rd[3] ), .A2(
        \UUT/Mcontrol/x_rd[4] ), .ZN(\UUT/Mcontrol/bp_logicA/N5 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C20  ( .A1(\UUT/Mcontrol/x_rd[2] ), .A2(
        \UUT/Mcontrol/bp_logicA/N5 ), .ZN(\UUT/Mcontrol/bp_logicA/N6 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C21  ( .A1(\UUT/Mcontrol/x_rd[1] ), .A2(
        \UUT/Mcontrol/bp_logicA/N6 ), .ZN(\UUT/Mcontrol/bp_logicA/N7 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C22  ( .A1(\UUT/Mcontrol/x_rd[0] ), .A2(
        \UUT/Mcontrol/bp_logicA/N7 ), .ZN(\UUT/Mcontrol/bp_logicA/N8 ) );
  INV_X2 \UUT/Mcontrol/bp_logicA/I_1  ( .A(\UUT/x_we ), .ZN(
        \UUT/Mcontrol/bp_logicA/N9 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C26  ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), 
        .A2(\UUT/Mcontrol/m_sampled_xrd[4] ), .ZN(\UUT/Mcontrol/bp_logicA/N10 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C27  ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N10 ), .ZN(\UUT/Mcontrol/bp_logicA/N11 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C28  ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N11 ), .ZN(\UUT/Mcontrol/bp_logicA/N12 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C29  ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N12 ), .ZN(\UUT/Mcontrol/bp_logicA/N13 )
         );
  INV_X2 \UUT/Mcontrol/bp_logicA/I_3  ( .A(\UUT/m_we ), .ZN(
        \UUT/Mcontrol/bp_logicA/N14 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C36  ( .A1(\UUT/Mcontrol/bp_logicA/N15 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N9 ), .ZN(
        \UUT/Mcontrol/bp_logicA/exec_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C37  ( .A1(\UUT/Mcontrol/bp_logicA/N2 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N8 ), .ZN(\UUT/Mcontrol/bp_logicA/N15 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C38  ( .A1(\UUT/Mcontrol/bp_logicA/N16 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N14 ), .ZN(
        \UUT/Mcontrol/bp_logicA/memory_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C39  ( .A1(\UUT/Mcontrol/bp_logicA/N3 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N13 ), .ZN(\UUT/Mcontrol/bp_logicA/N16 )
         );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_0  ( .A(\UUT/Mcontrol/d_jump_type[3] ), .ZN(\UUT/Mcontrol/st_logic/N103 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C198  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N114 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N115 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_3  ( .A(\UUT/Mcontrol/d_jump_type[0] ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N120 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C208  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N122 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N123 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_10  ( .A(
        \UUT/Mcontrol/d_jump_type[2] ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N223 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C318  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N226 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N227 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C319  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N227 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N228 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C320  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N228 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N229 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_12  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N229 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N230 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C326  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N232 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N233 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C327  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N233 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N234 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C328  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N234 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N235 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C333  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N238 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N239 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C334  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N239 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N240 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C335  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N240 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N241 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_14  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N241 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N242 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C340  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N244 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N245 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C342  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N246 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N247 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_15  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N247 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N248 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C346  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N250 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N251 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C348  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N252 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N253 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_16  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N253 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N254 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C354  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N256 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N257 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C356  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N258 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N259 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_17  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N259 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N260 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C361  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N262 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N263 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C363  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N264 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N265 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_18  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N265 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N266 ) );
  AND2_X2 \UUT/Mcontrol/Nextpc_decoding/C397  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N222 ), .A2(n6860), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N32 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_0  ( .A(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1875 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_1  ( .A(
        \UUT/Mcontrol/d_instr [30]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1876 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_2  ( .A(
        \UUT/Mcontrol/d_sampled_finstr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1877 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2052  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1878 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1879 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2053  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1879 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1880 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2054  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1880 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1881 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2055  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1881 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1882 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2058  ( .A1(
        \UUT/Mcontrol/d_instr [4]), .A2(\UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1883 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2059  ( .A1(
        \UUT/Mcontrol/d_instr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1883 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1884 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2060  ( .A1(
        \UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1884 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1885 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2061  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1885 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1886 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2062  ( .A1(
        \UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1886 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1887 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_4  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1887 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1888 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2068  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1889 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1890 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2069  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1890 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1891 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2070  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1891 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1892 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2071  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1892 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1893 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2074  ( .A1(
        \UUT/Mcontrol/d_instr [4]), .A2(\UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1894 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2075  ( .A1(
        \UUT/Mcontrol/d_instr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1894 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1895 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2076  ( .A1(
        \UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1895 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1896 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2077  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1896 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1897 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2078  ( .A1(
        \UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1897 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1898 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_6  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1898 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1899 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_7  ( .A(
        \UUT/Mcontrol/d_instr [4]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1900 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_8  ( .A(
        \UUT/Mcontrol/d_instr [0]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1901 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2082  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1900 ), .A2(
        \UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1902 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2083  ( .A1(
        \UUT/Mcontrol/d_instr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1902 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1903 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2084  ( .A1(
        \UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1903 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1904 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2085  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1904 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1905 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2086  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1901 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1905 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1906 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_9  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1906 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1907 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2088  ( .A1(
        \UUT/Mcontrol/d_instr [4]), .A2(\UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1908 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2089  ( .A1(
        \UUT/Mcontrol/d_instr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1908 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1909 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2090  ( .A1(
        \UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1909 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1910 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2091  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1910 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1911 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2092  ( .A1(
        \UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1911 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1912 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_10  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1912 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1913 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2094  ( .A1(
        \UUT/Mcontrol/d_instr [6]), .A2(\UUT/Mcontrol/d_instr [7]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1914 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_11  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1914 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1915 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2100  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1916 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1917 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2101  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1917 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1918 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2102  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1918 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1919 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2103  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1919 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1920 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_13  ( .A(
        \UUT/Mcontrol/d_instr [27]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1921 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2109  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1923 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1924 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2110  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1924 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1925 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2111  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1925 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1926 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2112  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1926 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1927 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_15  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1927 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1928 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2117  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1929 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1930 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2118  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1930 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1931 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2119  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1931 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1932 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2120  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1932 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1933 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_16  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1933 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1934 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2125  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1935 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1936 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2126  ( .A1(n6539), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1936 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1937 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2127  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1937 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1938 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2128  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1938 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1939 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_17  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1939 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1940 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2132  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1941 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1942 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2133  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1942 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1943 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2134  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1943 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1944 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2142  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1947 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1948 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2143  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1948 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1949 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2144  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1949 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1950 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2145  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1950 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1951 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_19  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1951 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1952 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2151  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1953 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1954 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2152  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1954 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1955 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2153  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1955 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1956 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2154  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1956 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1957 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_20  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1957 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1958 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2160  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1959 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1960 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2161  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1960 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1961 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2162  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1961 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1962 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2163  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1962 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1963 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2168  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1965 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1966 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2169  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1966 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1967 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2170  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1967 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1968 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2171  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1968 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1969 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2177  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1971 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1972 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2178  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1972 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1973 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2179  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1973 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1974 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2180  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1974 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1975 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2186  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1977 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1978 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2187  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1978 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1979 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2188  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1979 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1980 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2189  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1980 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1981 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2194  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1983 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1984 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2195  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1984 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1985 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2196  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1985 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1986 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2197  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1986 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1987 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_26  ( .A(n6541), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1989 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2204  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1990 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1991 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2205  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1991 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1992 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2206  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1992 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1993 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2207  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1993 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1994 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2214  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1996 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1997 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2215  ( .A1(n6541), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1997 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1998 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2216  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1998 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1999 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2222  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2002 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2003 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2223  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2003 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2004 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2224  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2004 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2005 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2231  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2008 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2009 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2232  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2009 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2010 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2240  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2014 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2015 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2241  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2015 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2016 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2242  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2016 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2017 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2248  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2020 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2021 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2249  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2021 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2022 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2250  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2022 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2023 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2256  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2026 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2027 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2257  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2027 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2028 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2258  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2028 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2029 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2259  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2029 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2030 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2263  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2032 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2033 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2264  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2033 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2034 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2265  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2034 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2035 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2270  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2038 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2039 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2271  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2039 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2040 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2272  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2040 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2041 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2279  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2044 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2045 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2280  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2045 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2046 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2281  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2046 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2047 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2287  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2050 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2051 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2288  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2051 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2052 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2289  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2052 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2053 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2290  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2053 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2054 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2295  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2056 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2057 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2296  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2057 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2058 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2297  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2058 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2059 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2298  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2059 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2060 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2302  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2062 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2063 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2303  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2063 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2064 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2304  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2064 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2065 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2305  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2065 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2066 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2310  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2068 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2069 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2311  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2069 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2070 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2312  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2070 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2071 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2317  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2074 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2075 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2318  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2075 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2076 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2319  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2076 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2077 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2324  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2080 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2081 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2325  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2081 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2082 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2326  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2082 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2083 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2327  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2083 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2084 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2330  ( .A1(
        \UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2086 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2087 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2331  ( .A1(n6540), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2087 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2088 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2332  ( .A1(
        \UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2088 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2089 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2606  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1913 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1915 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N62 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2608  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1882 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1888 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1871 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2610  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1893 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1899 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1873 ) );
  AND2_X2 \UUT/Mcontrol/C112  ( .A1(\UUT/Mcontrol/N19 ), .A2(net54843), .ZN(
        I_BUSY) );
  INV_X2 \UUT/BYP_BRANCH_MUXB/I_1  ( .A(\UUT/byp_controlB[2] ), .ZN(
        \UUT/BYP_BRANCH_MUXB/N39 ) );
  OR2_X2 \UUT/regfile/C1388  ( .A1(\UUT/rs1_addr [3]), .A2(\UUT/rs1_addr [4]), 
        .ZN(\UUT/regfile/N260 ) );
  OR2_X2 \UUT/regfile/C1389  ( .A1(\UUT/rs1_addr [2]), .A2(\UUT/regfile/N260 ), 
        .ZN(\UUT/regfile/N261 ) );
  OR2_X2 \UUT/regfile/C1390  ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/regfile/N261 ), 
        .ZN(\UUT/regfile/N262 ) );
  OR2_X2 \UUT/regfile/C1394  ( .A1(\UUT/rs2_addr [3]), .A2(\UUT/rs2_addr [4]), 
        .ZN(\UUT/regfile/N265 ) );
  OR2_X2 \UUT/regfile/C1395  ( .A1(\UUT/rs2_addr [2]), .A2(\UUT/regfile/N265 ), 
        .ZN(\UUT/regfile/N266 ) );
  OR2_X2 \UUT/regfile/C1396  ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/regfile/N266 ), 
        .ZN(\UUT/regfile/N267 ) );
  OR2_X2 \UUT/regfile/C1401  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N272 ) );
  OR2_X2 \UUT/regfile/C1402  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N272 ), 
        .ZN(\UUT/regfile/N273 ) );
  OR2_X2 \UUT/regfile/C1408  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N279 ) );
  OR2_X2 \UUT/regfile/C1409  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N279 ), 
        .ZN(\UUT/regfile/N280 ) );
  OR2_X2 \UUT/regfile/C1416  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N285 ) );
  OR2_X2 \UUT/regfile/C1417  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N285 ), 
        .ZN(\UUT/regfile/N286 ) );
  INV_X2 \UUT/regfile/I_7  ( .A(\UUT/rd_addr [2]), .ZN(\UUT/regfile/N290 ) );
  OR2_X2 \UUT/regfile/C1423  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N292 ) );
  OR2_X2 \UUT/regfile/C1424  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N292 ), .ZN(\UUT/regfile/N293 ) );
  OR2_X2 \UUT/regfile/C1431  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N298 ) );
  OR2_X2 \UUT/regfile/C1432  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N298 ), .ZN(\UUT/regfile/N299 ) );
  OR2_X2 \UUT/regfile/C1439  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N304 ) );
  OR2_X2 \UUT/regfile/C1440  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N304 ), .ZN(\UUT/regfile/N305 ) );
  OR2_X2 \UUT/regfile/C1448  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N310 ) );
  OR2_X2 \UUT/regfile/C1449  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N310 ), .ZN(\UUT/regfile/N311 ) );
  INV_X2 \UUT/regfile/I_12  ( .A(\UUT/rd_addr [3]), .ZN(\UUT/regfile/N315 ) );
  OR2_X2 \UUT/regfile/C1455  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N317 ) );
  OR2_X2 \UUT/regfile/C1456  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N317 ), 
        .ZN(\UUT/regfile/N318 ) );
  OR2_X2 \UUT/regfile/C1463  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N323 ) );
  OR2_X2 \UUT/regfile/C1464  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N323 ), 
        .ZN(\UUT/regfile/N324 ) );
  OR2_X2 \UUT/regfile/C1471  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N329 ) );
  OR2_X2 \UUT/regfile/C1472  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N329 ), 
        .ZN(\UUT/regfile/N330 ) );
  OR2_X2 \UUT/regfile/C1480  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N335 ) );
  OR2_X2 \UUT/regfile/C1481  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N335 ), 
        .ZN(\UUT/regfile/N336 ) );
  OR2_X2 \UUT/regfile/C1488  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N341 ) );
  OR2_X2 \UUT/regfile/C1489  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N341 ), .ZN(\UUT/regfile/N342 ) );
  OR2_X2 \UUT/regfile/C1497  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N347 ) );
  OR2_X2 \UUT/regfile/C1498  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N347 ), .ZN(\UUT/regfile/N348 ) );
  OR2_X2 \UUT/regfile/C1506  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N353 ) );
  OR2_X2 \UUT/regfile/C1507  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N353 ), .ZN(\UUT/regfile/N354 ) );
  OR2_X2 \UUT/regfile/C1516  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N359 ) );
  OR2_X2 \UUT/regfile/C1517  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N359 ), .ZN(\UUT/regfile/N360 ) );
  INV_X2 \UUT/regfile/I_21  ( .A(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N455 )
         );
  OR2_X2 \UUT/regfile/C1523  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N366 ) );
  OR2_X2 \UUT/regfile/C1524  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N366 ), 
        .ZN(\UUT/regfile/N367 ) );
  OR2_X2 \UUT/regfile/C1531  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N372 ) );
  OR2_X2 \UUT/regfile/C1532  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N372 ), 
        .ZN(\UUT/regfile/N373 ) );
  OR2_X2 \UUT/regfile/C1539  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N378 ) );
  OR2_X2 \UUT/regfile/C1540  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N378 ), 
        .ZN(\UUT/regfile/N379 ) );
  OR2_X2 \UUT/regfile/C1548  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N384 ) );
  OR2_X2 \UUT/regfile/C1549  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N384 ), 
        .ZN(\UUT/regfile/N385 ) );
  OR2_X2 \UUT/regfile/C1556  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N390 ) );
  OR2_X2 \UUT/regfile/C1557  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N390 ), .ZN(\UUT/regfile/N391 ) );
  OR2_X2 \UUT/regfile/C1565  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N396 ) );
  OR2_X2 \UUT/regfile/C1566  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N396 ), .ZN(\UUT/regfile/N397 ) );
  OR2_X2 \UUT/regfile/C1574  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N402 ) );
  OR2_X2 \UUT/regfile/C1575  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N402 ), .ZN(\UUT/regfile/N403 ) );
  OR2_X2 \UUT/regfile/C1584  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N408 ) );
  OR2_X2 \UUT/regfile/C1585  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N408 ), .ZN(\UUT/regfile/N409 ) );
  OR2_X2 \UUT/regfile/C1592  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N414 ) );
  OR2_X2 \UUT/regfile/C1593  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N414 ), 
        .ZN(\UUT/regfile/N415 ) );
  OR2_X2 \UUT/regfile/C1601  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N420 ) );
  OR2_X2 \UUT/regfile/C1602  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N420 ), 
        .ZN(\UUT/regfile/N421 ) );
  OR2_X2 \UUT/regfile/C1610  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N426 ) );
  OR2_X2 \UUT/regfile/C1611  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N426 ), 
        .ZN(\UUT/regfile/N427 ) );
  OR2_X2 \UUT/regfile/C1620  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N432 ) );
  OR2_X2 \UUT/regfile/C1621  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N432 ), 
        .ZN(\UUT/regfile/N433 ) );
  OR2_X2 \UUT/regfile/C1629  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N438 ) );
  OR2_X2 \UUT/regfile/C1630  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N438 ), .ZN(\UUT/regfile/N439 ) );
  OR2_X2 \UUT/regfile/C1639  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N444 ) );
  OR2_X2 \UUT/regfile/C1640  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N444 ), .ZN(\UUT/regfile/N445 ) );
  OR2_X2 \UUT/regfile/C1649  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N450 ) );
  OR2_X2 \UUT/regfile/C1650  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N450 ), .ZN(\UUT/regfile/N451 ) );
  OR2_X2 \UUT/regfile/C1660  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N456 ) );
  OR2_X2 \UUT/regfile/C1661  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N456 ), .ZN(\UUT/regfile/N457 ) );
  INV_X2 \UUT/I_2  ( .A(dmem_read), .ZN(\UUT/N76 ) );
  INV_X2 \UUT/I_3  ( .A(dmem_write), .ZN(\UUT/N77 ) );
  OR2_X2 \UUT/C150  ( .A1(\UUT/N76 ), .A2(\UUT/N77 ), .ZN(\UUT/N3 ) );
  AND2_X2 C271 ( .A1(N40), .A2(N41), .ZN(N178) );
  AND2_X2 C270 ( .A1(N178), .A2(N172), .ZN(N42) );
  AND2_X2 C268 ( .A1(N37), .A2(N38), .ZN(N177) );
  AND2_X2 C267 ( .A1(N177), .A2(N171), .ZN(N43) );
  AND2_X2 C265 ( .A1(N33), .A2(N34), .ZN(N176) );
  AND2_X2 C264 ( .A1(N176), .A2(N168), .ZN(N35) );
  AND2_X2 C262 ( .A1(N29), .A2(N30), .ZN(N175) );
  AND2_X2 C261 ( .A1(N175), .A2(N165), .ZN(N31) );
  AND2_X2 C259 ( .A1(N24), .A2(N25), .ZN(N174) );
  AND2_X2 C258 ( .A1(N174), .A2(N26), .ZN(N27) );
  AND2_X2 C256 ( .A1(N19), .A2(N20), .ZN(N173) );
  AND2_X2 C255 ( .A1(N173), .A2(N21), .ZN(N22) );
  INV_X2 I_19 ( .A(I_BUSY), .ZN(iram_rd) );
  AND2_X2 C246 ( .A1(D_ADDR_OUTBUS[0]), .A2(D_ADDR_OUTBUS[1]), .ZN(N172) );
  INV_X2 I_18 ( .A(N170), .ZN(N171) );
  OR2_X2 C244 ( .A1(D_ADDR_OUTBUS[0]), .A2(N169), .ZN(N170) );
  INV_X2 I_17 ( .A(D_ADDR_OUTBUS[1]), .ZN(N169) );
  INV_X2 I_16 ( .A(N167), .ZN(N168) );
  OR2_X2 C241 ( .A1(N166), .A2(D_ADDR_OUTBUS[1]), .ZN(N167) );
  INV_X2 I_15 ( .A(D_ADDR_OUTBUS[0]), .ZN(N166) );
  INV_X2 I_14 ( .A(N164), .ZN(N165) );
  OR2_X2 C238 ( .A1(D_ADDR_OUTBUS[0]), .A2(D_ADDR_OUTBUS[1]), .ZN(N164) );
  INV_X2 I_13 ( .A(N13), .ZN(N41) );
  INV_X2 I_12 ( .A(N12), .ZN(N40) );
  INV_X2 I_11 ( .A(N11), .ZN(N38) );
  INV_X2 I_10 ( .A(N10), .ZN(N37) );
  INV_X2 I_9 ( .A(N9), .ZN(N34) );
  INV_X2 I_8 ( .A(N8), .ZN(N33) );
  INV_X2 I_7 ( .A(N7), .ZN(N30) );
  INV_X2 I_6 ( .A(N6), .ZN(N29) );
  INV_X2 I_5 ( .A(N5), .ZN(N26) );
  INV_X2 I_4 ( .A(N4), .ZN(N25) );
  INV_X2 I_3 ( .A(N3), .ZN(N24) );
  INV_X2 I_2 ( .A(N2), .ZN(N21) );
  INV_X2 I_1 ( .A(N1), .ZN(N20) );
  INV_X2 I_0 ( .A(N0), .ZN(N19) );
  DFFS_X1 \localbus/c2_op_reg[MASTER]  ( .D(\localbus/c1_op[MASTER] ), .CK(CLK), .SN(\UUT/Mcontrol/int_reset ), .Q(\localbus/c2_op[MASTER] ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[0]  ( .D(n4335), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[0] ), .QN(
        \UUT/Mpath/the_alu/N84 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[31]  ( .D(n4334), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [31]) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[2]  ( .D(n4333), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [2]), .QN(
        \UUT/Mpath/N111 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[0]  ( .D(n4332), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[0] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[0]  ( .D(n4331), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5677) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[0]  ( .D(n4330), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[32] ), 
        .QN(n5709) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[31]  ( .D(n4328), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5455) );
  DFFR_X1 \localbus/c2_op_reg[SLAVE][1]  ( .D(1'b0), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\localbus/c2_op[SLAVE][1] ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[10]  ( .D(n4325), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[10] ), .QN(
        \UUT/Mpath/the_alu/N64 ) );
  DFFR_X1 \localbus/c2_op_reg[SLAVE][0]  ( .D(\localbus/c1_op[SLAVE][0] ), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\localbus/c2_op[SLAVE][0] ), .QN(\localbus/N219 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[8]  ( .D(n4324), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[8] ), .QN(
        \UUT/Mpath/the_alu/N68 ) );
  DFFS_X1 \localbus/c2_op_reg[SLAVE][2]  ( .D(\localbus/N227 ), .CK(CLK), .SN(
        \UUT/Mcontrol/int_reset ), .Q(\localbus/c2_op[SLAVE][2] ) );
  DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[0]  ( .D(n4322), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/mem_baddr [0]), .QN(
        \UUT/Mpath/the_memhandle/N240 ) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[0]  ( .D(n4321), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5527) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[63]  ( .D(n4320), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[63] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[62]  ( .D(n4319), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[62] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[61]  ( .D(n4318), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[61] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[60]  ( .D(n4317), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[60] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[59]  ( .D(n4316), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[59] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[58]  ( .D(n4315), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[58] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[57]  ( .D(n4314), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[57] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[56]  ( .D(n4313), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[56] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[55]  ( .D(n4312), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[55] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[54]  ( .D(n4311), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[54] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[53]  ( .D(n4310), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[53] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[52]  ( .D(n4309), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[52] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[51]  ( .D(n4308), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[51] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[49]  ( .D(n4306), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[49] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[48]  ( .D(n4305), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[48] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[47]  ( .D(n4304), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[47] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[46]  ( .D(n4303), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[46] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[45]  ( .D(n4302), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[45] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[44]  ( .D(n4301), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[44] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[43]  ( .D(n4300), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[43] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[42]  ( .D(n4299), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[42] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[41]  ( .D(n4298), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[41] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[40]  ( .D(n4297), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[40] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[39]  ( .D(n4296), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[39] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[38]  ( .D(n4295), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[38] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[37]  ( .D(n4294), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[37] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[36]  ( .D(n4293), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[36] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[35]  ( .D(n4292), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[35] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[34]  ( .D(n4291), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[34] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[33]  ( .D(n4290), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[33] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[32]  ( .D(n4289), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[32] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[31]  ( .D(n4288), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[31] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[30]  ( .D(n4287), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[30] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[29]  ( .D(n4286), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[29] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[28]  ( .D(n4285), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[28] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[27]  ( .D(n4284), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[27] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[26]  ( .D(n4283), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[26] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[25]  ( .D(n4282), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[25] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[24]  ( .D(n4281), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[24] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[23]  ( .D(n4280), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[23] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[22]  ( .D(n4279), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[22] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[21]  ( .D(n4278), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[21] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[20]  ( .D(n4277), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[20] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[19]  ( .D(n4276), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[19] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[18]  ( .D(n4275), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[18] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[17]  ( .D(n4274), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[17] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[16]  ( .D(n4273), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[16] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[15]  ( .D(n4272), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[15] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[14]  ( .D(n4271), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[14] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[13]  ( .D(n4270), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[13] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[12]  ( .D(n4269), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[12] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[11]  ( .D(n4268), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[11] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[10]  ( .D(n4267), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[10] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[9]  ( .D(n4266), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[9] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[8]  ( .D(n4265), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[8] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[7]  ( .D(n4264), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[7] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[6]  ( .D(n4263), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[6] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[5]  ( .D(n4262), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[5] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[4]  ( .D(n4261), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[4] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[3]  ( .D(n4260), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[3] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[2]  ( .D(n4259), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[2] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[1]  ( .D(n4258), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[1] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[0]  ( .D(n4257), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[0] ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[0]  ( .D(n4255), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [0]), 
        .QN(\UUT/Mcontrol/st_logic/N34 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[30]  ( .D(n4254), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [30]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[29]  ( .D(n4253), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [29]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[28]  ( .D(n4252), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [28]), .QN(n2785)
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[27]  ( .D(n4251), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [27]), .QN(n2784)
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[26]  ( .D(n4250), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [26]), .QN(n2783)
         );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[SIGN]  ( .D(n4249), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[SIGN] ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MW]  ( .D(n4248), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[MW] ), .QN(n2781) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MR]  ( .D(n4247), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[MR] ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MH]  ( .D(n4246), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[MH] ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MB]  ( .D(n4245), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[MB] ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[25]  ( .D(n4244), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [25]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[24]  ( .D(n4243), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [24]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[23]  ( .D(n4242), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [23]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[22]  ( .D(n4241), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [22]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[21]  ( .D(n4240), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [21]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[20]  ( .D(n4239), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [20]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[19]  ( .D(n4238), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [19]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[18]  ( .D(n4237), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [18]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[17]  ( .D(n4236), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [17]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[16]  ( .D(n4235), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [16]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[15]  ( .D(n4234), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [15]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[14]  ( .D(n4233), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [14]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[13]  ( .D(n4232), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [13]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[12]  ( .D(n4231), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [12]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[11]  ( .D(n4230), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [11]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[10]  ( .D(n4229), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [10]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[9]  ( .D(n4228), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [9]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[8]  ( .D(n4227), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [8]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[7]  ( .D(n4226), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [7]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[6]  ( .D(n4225), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [6]) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[5]  ( .D(n4224), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [5]) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[5]  ( .D(n4223), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [5]), 
        .QN(n2756) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[5]  ( .D(n4222), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[5] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[5]  ( .D(n4221), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[5] ), .QN(n2754) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[4]  ( .D(n4220), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [4]) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[4]  ( .D(n4219), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [4]), 
        .QN(n2752) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[4]  ( .D(n4218), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[4] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[4]  ( .D(n4217), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[4] ), .QN(n2750) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[3]  ( .D(n4216), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [3]) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[3]  ( .D(n4215), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [3]), 
        .QN(n2748) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[3]  ( .D(n4214), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[3] ), .QN(\UUT/Mpath/the_mult/N192 )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[3]  ( .D(n4213), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[3] ), .QN(\UUT/Mpath/the_mult/N229 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[2]  ( .D(n4212), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [2]) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[2]  ( .D(n4211), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mcontrol/st_logic/N26 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[2]  ( .D(n4210), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[2] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[2]  ( .D(n4209), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[2] ), .QN(\UUT/Mpath/the_mult/N244 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[1]  ( .D(n4208), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [1]) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[1]  ( .D(n4207), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mcontrol/st_logic/N27 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[1]  ( .D(n4206), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[1] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[1]  ( .D(n4205), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[1] ), .QN(\UUT/Mpath/the_mult/N230 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[0]  ( .D(n4204), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [0]) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[0]  ( .D(n4203), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[0] ), .QN(\UUT/Mpath/the_mult/N193 )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[0]  ( .D(n4202), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[0] ), .QN(\UUT/Mpath/the_mult/N231 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[4]  ( .D(n4201), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[4] ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[4]  ( .D(n4200), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[4] ), .QN(
        n2741) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[3]  ( .D(n4199), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[3] ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[3]  ( .D(n4198), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[3] ), .QN(
        n2739) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[2]  ( .D(n4197), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[2] ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[2]  ( .D(n4196), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[2] ), .QN(
        n2737) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[1]  ( .D(n4195), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[1] ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[1]  ( .D(n4194), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[1] ), .QN(
        n2735) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[0]  ( .D(n4193), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[0] ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[0]  ( .D(n4192), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[0] ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[10]  ( .D(n4191), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [10]), .QN(
        n2732) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_rf_we_reg  ( .D(n4190), .CK(CLK), .SN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/x_we ), .QN(
        \UUT/Mcontrol/bp_logicB/N9 ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_rf_we_reg  ( .D(n4189), .CK(CLK), .SN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/m_we ), .QN(n5413) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[0]  ( .D(n4188), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[0] ), 
        .QN(n5676) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[0]  ( .D(n4187), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5092) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[10]  ( .D(n4186), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5091) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[31]  ( .D(n4185), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5068) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[8]  ( .D(n4184), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5062) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[0]  ( .D(n4183), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4644) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[10]  ( .D(n4182), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4643) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[31]  ( .D(n4181), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4620) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[8]  ( .D(n4180), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4614) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[0]  ( .D(n4179), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][0] ), .QN(n4580)
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[10]  ( .D(n4178), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][10] ), .QN(n4579) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[31]  ( .D(n4177), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][31] ), .QN(n4556) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[8]  ( .D(n4176), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][8] ), .QN(n4550)
         );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[0]  ( .D(n4175), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4516) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[10]  ( .D(n4174), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4515) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[31]  ( .D(n4173), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4492) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[8]  ( .D(n4172), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4486) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[0]  ( .D(n4171), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4452) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[10]  ( .D(n4170), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4451) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[31]  ( .D(n4169), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4428) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[8]  ( .D(n4168), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4422) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[0]  ( .D(n4167), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5380) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[10]  ( .D(n4166), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5379) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[31]  ( .D(n4165), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5356) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[8]  ( .D(n4164), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5350) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[0]  ( .D(n4163), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5316) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[10]  ( .D(n4162), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5315) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[31]  ( .D(n4161), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5292) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[8]  ( .D(n4160), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5286) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[0]  ( .D(n4159), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5252) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[10]  ( .D(n4158), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5251) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[31]  ( .D(n4157), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5228) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[8]  ( .D(n4156), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5222) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[0]  ( .D(n4155), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5188) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[10]  ( .D(n4154), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5187) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[31]  ( .D(n4153), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5164) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[8]  ( .D(n4152), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5158) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[0]  ( .D(n4151), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][0] ), .QN(n5124) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[10]  ( .D(n4150), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][10] ), .QN(
        n5123) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[31]  ( .D(n4149), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][31] ), .QN(
        n5100) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[8]  ( .D(n4148), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][8] ), .QN(n5094) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[0]  ( .D(n4147), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][0] ), .QN(n5028) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[10]  ( .D(n4146), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][10] ), .QN(
        n5027) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[31]  ( .D(n4145), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][31] ), .QN(
        n5004) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[8]  ( .D(n4144), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][8] ), .QN(n4998) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[0]  ( .D(n4143), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4964) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[10]  ( .D(n4142), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4963) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[31]  ( .D(n4141), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4940) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[8]  ( .D(n4140), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4934) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[0]  ( .D(n4139), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][0] ), .QN(n4900) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[10]  ( .D(n4138), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][10] ), .QN(
        n4899) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[31]  ( .D(n4137), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][31] ), .QN(
        n4876) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[8]  ( .D(n4136), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][8] ), .QN(n4870) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[0]  ( .D(n4135), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4836) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[10]  ( .D(n4134), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4835) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[31]  ( .D(n4133), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4812) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[8]  ( .D(n4132), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4806) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[0]  ( .D(n4131), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][0] ), .QN(n4772) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[10]  ( .D(n4130), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][10] ), .QN(
        n4771) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[31]  ( .D(n4129), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][31] ), .QN(
        n4748) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[8]  ( .D(n4128), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][8] ), .QN(n4742) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[0]  ( .D(n4127), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4676) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[10]  ( .D(n4126), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4675) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[31]  ( .D(n4125), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4652) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[8]  ( .D(n4124), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4646) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[0]  ( .D(n4123), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4740) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[10]  ( .D(n4122), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4739) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[31]  ( .D(n4121), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4716) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[8]  ( .D(n4120), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4710) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[0]  ( .D(n4119), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][0] ), .QN(n4612)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[10]  ( .D(n4118), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][10] ), .QN(n4611) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[31]  ( .D(n4117), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][31] ), .QN(n4588) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[8]  ( .D(n4116), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][8] ), .QN(n4582)
         );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[0]  ( .D(n4115), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4548) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[10]  ( .D(n4114), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4547) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[31]  ( .D(n4113), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4524) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[8]  ( .D(n4112), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4518) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[0]  ( .D(n4111), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4484) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[10]  ( .D(n4110), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4483) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[31]  ( .D(n4109), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4460) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[8]  ( .D(n4108), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4454) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[0]  ( .D(n4107), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5412) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[10]  ( .D(n4106), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5411) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[31]  ( .D(n4105), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5388) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[8]  ( .D(n4104), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5382) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[0]  ( .D(n4103), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5348) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[10]  ( .D(n4102), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5347) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[31]  ( .D(n4101), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5324) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[8]  ( .D(n4100), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5318) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[0]  ( .D(n4099), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5284) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[10]  ( .D(n4098), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5283) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[31]  ( .D(n4097), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5260) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[8]  ( .D(n4096), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5254) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[0]  ( .D(n4095), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5220) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[10]  ( .D(n4094), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5219) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[31]  ( .D(n4093), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5196) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[8]  ( .D(n4092), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5190) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[0]  ( .D(n4091), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][0] ), .QN(n5156) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[10]  ( .D(n4090), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][10] ), .QN(
        n5155) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[31]  ( .D(n4089), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][31] ), .QN(
        n5132) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[8]  ( .D(n4088), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][8] ), .QN(n5126) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[0]  ( .D(n4087), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][0] ), .QN(n5060) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[10]  ( .D(n4086), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][10] ), .QN(
        n5059) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[31]  ( .D(n4085), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][31] ), .QN(
        n5036) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[8]  ( .D(n4084), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][8] ), .QN(n5030) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[0]  ( .D(n4083), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4996) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[10]  ( .D(n4082), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4995) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[31]  ( .D(n4081), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4972) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[8]  ( .D(n4080), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4966) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[0]  ( .D(n4079), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][0] ), .QN(n4932) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[10]  ( .D(n4078), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][10] ), .QN(
        n4931) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[31]  ( .D(n4077), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][31] ), .QN(
        n4908) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[8]  ( .D(n4076), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][8] ), .QN(n4902) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[0]  ( .D(n4075), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4868) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[10]  ( .D(n4074), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4867) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[31]  ( .D(n4073), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4844) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[8]  ( .D(n4072), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4838) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[0]  ( .D(n4071), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][0] ), .QN(n4804) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[10]  ( .D(n4070), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][10] ), .QN(
        n4803) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[31]  ( .D(n4069), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][31] ), .QN(
        n4780) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[8]  ( .D(n4068), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][8] ), .QN(n4774) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[0]  ( .D(n4067), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4708) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[10]  ( .D(n4066), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4707) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[31]  ( .D(n4065), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4684) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[8]  ( .D(n4064), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4678) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[SIGN]  ( .D(n4063), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/m_mem_command[SIGN] ), .QN(
        \UUT/Mpath/the_memhandle/N235 ) );
  DFFR_X1 \localbus/c2_op_reg[OP][0]  ( .D(\UUT/Mcontrol/st_logic/N15 ), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(\localbus/N293 ) );
  DFFR_X1 \localbus/c2_op_reg[OP][1]  ( .D(\localbus/c1_op[OP][1] ), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\localbus/c2_op[OP][1] ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MH]  ( .D(n4059), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mpath/the_memhandle/N238 ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MB]  ( .D(n4058), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mpath/the_memhandle/N236 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[31]  ( .D(n4056), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[31] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[31]  ( .D(n4055), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5629) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[31]  ( .D(n4054), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[31] ), .QN(
        n5628) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[1]  ( .D(n4053), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [1]), .QN(
        \UUT/Mpath/N116 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[0]  ( .D(n4052), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [0]), .QN(
        \UUT/Mpath/N112 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[2]  ( .D(n4051), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [2]), .QN(
        \UUT/Mpath/the_shift/N104 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[1]  ( .D(n4050), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [1]), .QN(
        \UUT/Mpath/the_shift/N112 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[0]  ( .D(n4049), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [0]), .QN(
        \UUT/Mpath/the_shift/N105 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][5]  ( .D(n4048), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][5] ), .QN(
        \UUT/Mpath/the_alu/N466 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][4]  ( .D(n4047), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][4] ), .QN(
        \UUT/Mpath/the_alu/N453 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][3]  ( .D(n4046), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][3] ), .QN(n2730) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][2]  ( .D(n4045), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][2] ), .QN(n2729) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][1]  ( .D(n4044), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][1] ), .QN(
        \UUT/Mpath/the_alu/N467 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][0]  ( .D(n4043), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][0] ), .QN(
        \UUT/Mpath/the_alu/N468 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[9]  ( .D(n4042), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [9]), .QN(
        n2728) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[23]  ( .D(n4041), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [23]), .QN(
        n2727) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[0]  ( .D(n4040), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[0] ) );
  DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[0]  ( .D(n4039), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [0]), .QN(
        n2725) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[1]  ( .D(n4038), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[1] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[2]  ( .D(n4037), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[2] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[3]  ( .D(n4036), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[3] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[4]  ( .D(n4035), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[4] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[5]  ( .D(n4034), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[5] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[6]  ( .D(n4033), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[6] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[7]  ( .D(n4032), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[7] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[8]  ( .D(n4031), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[8] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[9]  ( .D(n4030), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[9] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[10]  ( .D(n4029), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[10] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[11]  ( .D(n4028), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[11] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[12]  ( .D(n4027), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[12] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[13]  ( .D(n4026), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[13] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[14]  ( .D(n4025), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[14] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[15]  ( .D(n4024), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[15] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[16]  ( .D(n4023), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[16] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[17]  ( .D(n4022), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[17] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[18]  ( .D(n4021), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[18] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[19]  ( .D(n4020), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[19] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[20]  ( .D(n4019), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[20] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[21]  ( .D(n4018), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[21] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[22]  ( .D(n4017), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[22] ) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[23]  ( .D(n4016), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_jar[23] ) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[23]  ( .D(n4015), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5482) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[30]  ( .D(n4013), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5458) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[30]  ( .D(n4012), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4429) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[30]  ( .D(n4011), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4461) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[30]  ( .D(n4010), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4493) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[30]  ( .D(n4009), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4525) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[30]  ( .D(n4008), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][30] ), .QN(n4557) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[30]  ( .D(n4007), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][30] ), .QN(n4589) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[30]  ( .D(n4006), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4621) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[30]  ( .D(n4005), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4653) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[30]  ( .D(n4004), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4685) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[30]  ( .D(n4003), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4717) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[30]  ( .D(n4002), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][30] ), .QN(
        n4749) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[30]  ( .D(n4001), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][30] ), .QN(
        n4781) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[30]  ( .D(n4000), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4813) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[30]  ( .D(n3999), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4845) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[30]  ( .D(n3998), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][30] ), .QN(
        n4877) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[30]  ( .D(n3997), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][30] ), .QN(
        n4909) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[30]  ( .D(n3996), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4941) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[30]  ( .D(n3995), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4973) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[30]  ( .D(n3994), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][30] ), .QN(
        n5005) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[30]  ( .D(n3993), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][30] ), .QN(
        n5037) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[30]  ( .D(n3992), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5069) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[30]  ( .D(n3991), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][30] ), .QN(
        n5101) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[30]  ( .D(n3990), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][30] ), .QN(
        n5133) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[30]  ( .D(n3989), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5165) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[30]  ( .D(n3988), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5197) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[30]  ( .D(n3987), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5229) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[30]  ( .D(n3986), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5261) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[30]  ( .D(n3985), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5293) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[30]  ( .D(n3984), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5325) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[30]  ( .D(n3983), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5357) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[30]  ( .D(n3982), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5389) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[30]  ( .D(n3980), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[30] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[30]  ( .D(n3979), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5631) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[30]  ( .D(n3978), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[30] ), .QN(
        n5630) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[30]  ( .D(n3977), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[62] ), .QN(
        n5686) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[30]  ( .D(n3976), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[30] ), .QN(
        \UUT/Mpath/the_alu/N24 ) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[29]  ( .D(n3975), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5464) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[29]  ( .D(n3974), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4431) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[29]  ( .D(n3973), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4463) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[29]  ( .D(n3972), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4495) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[29]  ( .D(n3971), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4527) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[29]  ( .D(n3970), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][29] ), .QN(n4559) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[29]  ( .D(n3969), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][29] ), .QN(n4591) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[29]  ( .D(n3968), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4623) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[29]  ( .D(n3967), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4655) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[29]  ( .D(n3966), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4687) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[29]  ( .D(n3965), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4719) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[29]  ( .D(n3964), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][29] ), .QN(
        n4751) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[29]  ( .D(n3963), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][29] ), .QN(
        n4783) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[29]  ( .D(n3962), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4815) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[29]  ( .D(n3961), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4847) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[29]  ( .D(n3960), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][29] ), .QN(
        n4879) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[29]  ( .D(n3959), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][29] ), .QN(
        n4911) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[29]  ( .D(n3958), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4943) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[29]  ( .D(n3957), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4975) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[29]  ( .D(n3956), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][29] ), .QN(
        n5007) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[29]  ( .D(n3955), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][29] ), .QN(
        n5039) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[29]  ( .D(n3954), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5071) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[29]  ( .D(n3953), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][29] ), .QN(
        n5103) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[29]  ( .D(n3952), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][29] ), .QN(
        n5135) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[29]  ( .D(n3951), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5167) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[29]  ( .D(n3950), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5199) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[29]  ( .D(n3949), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5231) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[29]  ( .D(n3948), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5263) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[29]  ( .D(n3947), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5295) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[29]  ( .D(n3946), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5327) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[29]  ( .D(n3945), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5359) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[29]  ( .D(n3944), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5391) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[28]  ( .D(n3942), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5467) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[28]  ( .D(n3941), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4432) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[28]  ( .D(n3940), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4464) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[28]  ( .D(n3939), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4496) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[28]  ( .D(n3938), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4528) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[28]  ( .D(n3937), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][28] ), .QN(n4560) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[28]  ( .D(n3936), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][28] ), .QN(n4592) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[28]  ( .D(n3935), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4624) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[28]  ( .D(n3934), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4656) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[28]  ( .D(n3933), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4688) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[28]  ( .D(n3932), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4720) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[28]  ( .D(n3931), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][28] ), .QN(
        n4752) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[28]  ( .D(n3930), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][28] ), .QN(
        n4784) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[28]  ( .D(n3929), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4816) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[28]  ( .D(n3928), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4848) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[28]  ( .D(n3927), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][28] ), .QN(
        n4880) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[28]  ( .D(n3926), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][28] ), .QN(
        n4912) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[28]  ( .D(n3925), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4944) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[28]  ( .D(n3924), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4976) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[28]  ( .D(n3923), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][28] ), .QN(
        n5008) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[28]  ( .D(n3922), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][28] ), .QN(
        n5040) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[28]  ( .D(n3921), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5072) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[28]  ( .D(n3920), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][28] ), .QN(
        n5104) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[28]  ( .D(n3919), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][28] ), .QN(
        n5136) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[28]  ( .D(n3918), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5168) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[28]  ( .D(n3917), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5200) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[28]  ( .D(n3916), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5232) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[28]  ( .D(n3915), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5264) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[28]  ( .D(n3914), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5296) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[28]  ( .D(n3913), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5328) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[28]  ( .D(n3912), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5360) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[28]  ( .D(n3911), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5392) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[27]  ( .D(n3909), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5470) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[27]  ( .D(n3908), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4433) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[27]  ( .D(n3907), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4465) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[27]  ( .D(n3906), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4497) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[27]  ( .D(n3905), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4529) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[27]  ( .D(n3904), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][27] ), .QN(n4561) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[27]  ( .D(n3903), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][27] ), .QN(n4593) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[27]  ( .D(n3902), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4625) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[27]  ( .D(n3901), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4657) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[27]  ( .D(n3900), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4689) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[27]  ( .D(n3899), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4721) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[27]  ( .D(n3898), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][27] ), .QN(
        n4753) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[27]  ( .D(n3897), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][27] ), .QN(
        n4785) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[27]  ( .D(n3896), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4817) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[27]  ( .D(n3895), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4849) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[27]  ( .D(n3894), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][27] ), .QN(
        n4881) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[27]  ( .D(n3893), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][27] ), .QN(
        n4913) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[27]  ( .D(n3892), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4945) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[27]  ( .D(n3891), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4977) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[27]  ( .D(n3890), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][27] ), .QN(
        n5009) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[27]  ( .D(n3889), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][27] ), .QN(
        n5041) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[27]  ( .D(n3888), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5073) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[27]  ( .D(n3887), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][27] ), .QN(
        n5105) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[27]  ( .D(n3886), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][27] ), .QN(
        n5137) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[27]  ( .D(n3885), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5169) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[27]  ( .D(n3884), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5201) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[27]  ( .D(n3883), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5233) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[27]  ( .D(n3882), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5265) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[27]  ( .D(n3881), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5297) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[27]  ( .D(n3880), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5329) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[27]  ( .D(n3879), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5361) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[27]  ( .D(n3878), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5393) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[26]  ( .D(n3876), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5473) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[26]  ( .D(n3875), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4434) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[26]  ( .D(n3874), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4466) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[26]  ( .D(n3873), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4498) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[26]  ( .D(n3872), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4530) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[26]  ( .D(n3871), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][26] ), .QN(n4562) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[26]  ( .D(n3870), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][26] ), .QN(n4594) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[26]  ( .D(n3869), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4626) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[26]  ( .D(n3868), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4658) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[26]  ( .D(n3867), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4690) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[26]  ( .D(n3866), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4722) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[26]  ( .D(n3865), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][26] ), .QN(
        n4754) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[26]  ( .D(n3864), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][26] ), .QN(
        n4786) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[26]  ( .D(n3863), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4818) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[26]  ( .D(n3862), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4850) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[26]  ( .D(n3861), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][26] ), .QN(
        n4882) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[26]  ( .D(n3860), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][26] ), .QN(
        n4914) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[26]  ( .D(n3859), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4946) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[26]  ( .D(n3858), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4978) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[26]  ( .D(n3857), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][26] ), .QN(
        n5010) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[26]  ( .D(n3856), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][26] ), .QN(
        n5042) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[26]  ( .D(n3855), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5074) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[26]  ( .D(n3854), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][26] ), .QN(
        n5106) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[26]  ( .D(n3853), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][26] ), .QN(
        n5138) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[26]  ( .D(n3852), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5170) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[26]  ( .D(n3851), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5202) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[26]  ( .D(n3850), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5234) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[26]  ( .D(n3849), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5266) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[26]  ( .D(n3848), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5298) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[26]  ( .D(n3847), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5330) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[26]  ( .D(n3846), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5362) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[26]  ( .D(n3845), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5394) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[25]  ( .D(n3843), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5476) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[25]  ( .D(n3842), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4435) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[25]  ( .D(n3841), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4467) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[25]  ( .D(n3840), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4499) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[25]  ( .D(n3839), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4531) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[25]  ( .D(n3838), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][25] ), .QN(n4563) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[25]  ( .D(n3837), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][25] ), .QN(n4595) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[25]  ( .D(n3836), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4627) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[25]  ( .D(n3835), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4659) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[25]  ( .D(n3834), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4691) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[25]  ( .D(n3833), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4723) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[25]  ( .D(n3832), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][25] ), .QN(
        n4755) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[25]  ( .D(n3831), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][25] ), .QN(
        n4787) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[25]  ( .D(n3830), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4819) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[25]  ( .D(n3829), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4851) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[25]  ( .D(n3828), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][25] ), .QN(
        n4883) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[25]  ( .D(n3827), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][25] ), .QN(
        n4915) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[25]  ( .D(n3826), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4947) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[25]  ( .D(n3825), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4979) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[25]  ( .D(n3824), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][25] ), .QN(
        n5011) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[25]  ( .D(n3823), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][25] ), .QN(
        n5043) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[25]  ( .D(n3822), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5075) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[25]  ( .D(n3821), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][25] ), .QN(
        n5107) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[25]  ( .D(n3820), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][25] ), .QN(
        n5139) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[25]  ( .D(n3819), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5171) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[25]  ( .D(n3818), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5203) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[25]  ( .D(n3817), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5235) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[25]  ( .D(n3816), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5267) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[25]  ( .D(n3815), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5299) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[25]  ( .D(n3814), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5331) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[25]  ( .D(n3813), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5363) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[25]  ( .D(n3812), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5395) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[1]  ( .D(n3810), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5494) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[1]  ( .D(n3809), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[1] ), .QN(
        \UUT/Mpath/the_alu/N82 ) );
  DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[1]  ( .D(n3808), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/mem_baddr [1]), .QN(
        \UUT/Mpath/the_memhandle/N239 ) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[23]  ( .D(n3807), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4437) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[23]  ( .D(n3806), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4469) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[23]  ( .D(n3805), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4501) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[23]  ( .D(n3804), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4533) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[23]  ( .D(n3803), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][23] ), .QN(n4565) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[23]  ( .D(n3802), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][23] ), .QN(n4597) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[23]  ( .D(n3801), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4629) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[23]  ( .D(n3800), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4661) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[23]  ( .D(n3799), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4693) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[23]  ( .D(n3798), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4725) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[23]  ( .D(n3797), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][23] ), .QN(
        n4757) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[23]  ( .D(n3796), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][23] ), .QN(
        n4789) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[23]  ( .D(n3795), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4821) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[23]  ( .D(n3794), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4853) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[23]  ( .D(n3793), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][23] ), .QN(
        n4885) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[23]  ( .D(n3792), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][23] ), .QN(
        n4917) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[23]  ( .D(n3791), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4949) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[23]  ( .D(n3790), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4981) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[23]  ( .D(n3789), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][23] ), .QN(
        n5013) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[23]  ( .D(n3788), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][23] ), .QN(
        n5045) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[23]  ( .D(n3787), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5077) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[23]  ( .D(n3786), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][23] ), .QN(
        n5109) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[23]  ( .D(n3785), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][23] ), .QN(
        n5141) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[23]  ( .D(n3784), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5173) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[23]  ( .D(n3783), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5205) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[23]  ( .D(n3782), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5237) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[23]  ( .D(n3781), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5269) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[23]  ( .D(n3780), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5301) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[23]  ( .D(n3779), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5333) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[23]  ( .D(n3778), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5365) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[23]  ( .D(n3777), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5397) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[23]  ( .D(n3775), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[23] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[23]  ( .D(n3774), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5647) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[23]  ( .D(n3773), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[23] ), .QN(
        n5646) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[23]  ( .D(n3772), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[55] ), .QN(
        n5694) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[1]  ( .D(n3771), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4441) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[1]  ( .D(n3770), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4473) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[1]  ( .D(n3769), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4505) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[1]  ( .D(n3768), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4537) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[1]  ( .D(n3767), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][1] ), .QN(n4569)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[1]  ( .D(n3766), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][1] ), .QN(n4601)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[1]  ( .D(n3765), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4633) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[1]  ( .D(n3764), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4665) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[1]  ( .D(n3763), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4697) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[1]  ( .D(n3762), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4729) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[1]  ( .D(n3761), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][1] ), .QN(n4761) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[1]  ( .D(n3760), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][1] ), .QN(n4793) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[1]  ( .D(n3759), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4825) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[1]  ( .D(n3758), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4857) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[1]  ( .D(n3757), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][1] ), .QN(n4889) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[1]  ( .D(n3756), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][1] ), .QN(n4921) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[1]  ( .D(n3755), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4953) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[1]  ( .D(n3754), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4985) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[1]  ( .D(n3753), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][1] ), .QN(n5017) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[1]  ( .D(n3752), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][1] ), .QN(n5049) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[1]  ( .D(n3751), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5081) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[1]  ( .D(n3750), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][1] ), .QN(n5113) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[1]  ( .D(n3749), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][1] ), .QN(n5145) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[1]  ( .D(n3748), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5177) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[1]  ( .D(n3747), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5209) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[1]  ( .D(n3746), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5241) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[1]  ( .D(n3745), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5273) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[1]  ( .D(n3744), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5305) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[1]  ( .D(n3743), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5337) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[1]  ( .D(n3742), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5369) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[1]  ( .D(n3741), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5401) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[1]  ( .D(n3739), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[1] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[1]  ( .D(n3738), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5655) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[1]  ( .D(n3737), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[1] ), 
        .QN(n5654) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[1]  ( .D(n3736), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[33] ), 
        .QN(n5698) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[1]  ( .D(n3734), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [1])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[2]  ( .D(n3733), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5461) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[2]  ( .D(n3732), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4430) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[2]  ( .D(n3731), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4462) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[2]  ( .D(n3730), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4494) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[2]  ( .D(n3729), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4526) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[2]  ( .D(n3728), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][2] ), .QN(n4558)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[2]  ( .D(n3727), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][2] ), .QN(n4590)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[2]  ( .D(n3726), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4622) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[2]  ( .D(n3725), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4654) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[2]  ( .D(n3724), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4686) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[2]  ( .D(n3723), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4718) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[2]  ( .D(n3722), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][2] ), .QN(n4750) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[2]  ( .D(n3721), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][2] ), .QN(n4782) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[2]  ( .D(n3720), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4814) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[2]  ( .D(n3719), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4846) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[2]  ( .D(n3718), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][2] ), .QN(n4878) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[2]  ( .D(n3717), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][2] ), .QN(n4910) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[2]  ( .D(n3716), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4942) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[2]  ( .D(n3715), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4974) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[2]  ( .D(n3714), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][2] ), .QN(n5006) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[2]  ( .D(n3713), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][2] ), .QN(n5038) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[2]  ( .D(n3712), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5070) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[2]  ( .D(n3711), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][2] ), .QN(n5102) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[2]  ( .D(n3710), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][2] ), .QN(n5134) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[2]  ( .D(n3709), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5166) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[2]  ( .D(n3708), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5198) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[2]  ( .D(n3707), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5230) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[2]  ( .D(n3706), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5262) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[2]  ( .D(n3705), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5294) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[2]  ( .D(n3704), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5326) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[2]  ( .D(n3703), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5358) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[2]  ( .D(n3702), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5390) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[2]  ( .D(n3700), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[2] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[2]  ( .D(n3699), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5633) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[2]  ( .D(n3698), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[2] ), 
        .QN(n5632) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[2]  ( .D(n3697), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[34] ), 
        .QN(n5687) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[2]  ( .D(n3696), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[2] ), .QN(
        \UUT/Mpath/the_alu/N80 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[2]  ( .D(n3695), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [2])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[2]  ( .D(n3694), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [2]), .QN(
        n2694) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[3]  ( .D(n3693), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5452) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[3]  ( .D(n3692), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4427) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[3]  ( .D(n3691), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4459) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[3]  ( .D(n3690), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4491) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[3]  ( .D(n3689), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4523) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[3]  ( .D(n3688), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][3] ), .QN(n4555)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[3]  ( .D(n3687), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][3] ), .QN(n4587)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[3]  ( .D(n3686), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4619) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[3]  ( .D(n3685), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4651) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[3]  ( .D(n3684), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4683) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[3]  ( .D(n3683), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4715) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[3]  ( .D(n3682), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][3] ), .QN(n4747) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[3]  ( .D(n3681), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][3] ), .QN(n4779) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[3]  ( .D(n3680), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4811) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[3]  ( .D(n3679), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4843) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[3]  ( .D(n3678), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][3] ), .QN(n4875) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[3]  ( .D(n3677), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][3] ), .QN(n4907) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[3]  ( .D(n3676), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4939) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[3]  ( .D(n3675), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4971) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[3]  ( .D(n3674), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][3] ), .QN(n5003) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[3]  ( .D(n3673), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][3] ), .QN(n5035) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[3]  ( .D(n3672), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5067) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[3]  ( .D(n3671), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][3] ), .QN(n5099) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[3]  ( .D(n3670), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][3] ), .QN(n5131) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[3]  ( .D(n3669), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5163) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[3]  ( .D(n3668), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5195) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[3]  ( .D(n3667), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5227) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[3]  ( .D(n3666), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5259) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[3]  ( .D(n3665), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5291) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[3]  ( .D(n3664), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5323) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[3]  ( .D(n3663), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5355) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[3]  ( .D(n3662), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5387) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[3]  ( .D(n3660), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[3] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[3]  ( .D(n3659), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5627) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[3]  ( .D(n3658), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[3] ), 
        .QN(n5626) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[3]  ( .D(n3657), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[35] ), 
        .QN(n5684) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[3]  ( .D(n3656), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[3] ), .QN(
        \UUT/Mpath/the_alu/N78 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[3]  ( .D(n3655), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [3])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[3]  ( .D(n3654), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [3]), .QN(
        n2691) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[4]  ( .D(n3653), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5449) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[4]  ( .D(n3652), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4426) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[4]  ( .D(n3651), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4458) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[4]  ( .D(n3650), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4490) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[4]  ( .D(n3649), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4522) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[4]  ( .D(n3648), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][4] ), .QN(n4554)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[4]  ( .D(n3647), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][4] ), .QN(n4586)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[4]  ( .D(n3646), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4618) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[4]  ( .D(n3645), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4650) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[4]  ( .D(n3644), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4682) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[4]  ( .D(n3643), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4714) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[4]  ( .D(n3642), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][4] ), .QN(n4746) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[4]  ( .D(n3641), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][4] ), .QN(n4778) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[4]  ( .D(n3640), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4810) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[4]  ( .D(n3639), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4842) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[4]  ( .D(n3638), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][4] ), .QN(n4874) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[4]  ( .D(n3637), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][4] ), .QN(n4906) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[4]  ( .D(n3636), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4938) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[4]  ( .D(n3635), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4970) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[4]  ( .D(n3634), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][4] ), .QN(n5002) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[4]  ( .D(n3633), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][4] ), .QN(n5034) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[4]  ( .D(n3632), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5066) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[4]  ( .D(n3631), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][4] ), .QN(n5098) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[4]  ( .D(n3630), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][4] ), .QN(n5130) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[4]  ( .D(n3629), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5162) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[4]  ( .D(n3628), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5194) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[4]  ( .D(n3627), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5226) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[4]  ( .D(n3626), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5258) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[4]  ( .D(n3625), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5290) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[4]  ( .D(n3624), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5322) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[4]  ( .D(n3623), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5354) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[4]  ( .D(n3622), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5386) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[4]  ( .D(n3620), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[4] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[4]  ( .D(n3619), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5625) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[4]  ( .D(n3618), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[4] ), 
        .QN(n5624) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[4]  ( .D(n3617), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[36] ), 
        .QN(n5683) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[4]  ( .D(n3616), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[4] ), .QN(
        \UUT/Mpath/the_alu/N76 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[4]  ( .D(n3615), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [4])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[4]  ( .D(n3614), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [4]), .QN(
        n2688) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[5]  ( .D(n3613), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5446) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[5]  ( .D(n3612), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4425) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[5]  ( .D(n3611), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4457) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[5]  ( .D(n3610), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4489) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[5]  ( .D(n3609), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4521) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[5]  ( .D(n3608), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][5] ), .QN(n4553)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[5]  ( .D(n3607), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][5] ), .QN(n4585)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[5]  ( .D(n3606), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4617) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[5]  ( .D(n3605), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4649) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[5]  ( .D(n3604), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4681) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[5]  ( .D(n3603), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4713) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[5]  ( .D(n3602), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][5] ), .QN(n4745) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[5]  ( .D(n3601), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][5] ), .QN(n4777) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[5]  ( .D(n3600), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4809) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[5]  ( .D(n3599), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4841) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[5]  ( .D(n3598), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][5] ), .QN(n4873) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[5]  ( .D(n3597), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][5] ), .QN(n4905) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[5]  ( .D(n3596), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4937) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[5]  ( .D(n3595), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4969) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[5]  ( .D(n3594), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][5] ), .QN(n5001) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[5]  ( .D(n3593), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][5] ), .QN(n5033) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[5]  ( .D(n3592), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5065) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[5]  ( .D(n3591), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][5] ), .QN(n5097) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[5]  ( .D(n3590), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][5] ), .QN(n5129) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[5]  ( .D(n3589), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5161) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[5]  ( .D(n3588), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5193) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[5]  ( .D(n3587), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5225) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[5]  ( .D(n3586), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5257) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[5]  ( .D(n3585), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5289) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[5]  ( .D(n3584), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5321) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[5]  ( .D(n3583), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5353) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[5]  ( .D(n3582), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5385) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[5]  ( .D(n3580), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[5] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[5]  ( .D(n3579), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5623) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[5]  ( .D(n3578), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[5] ), 
        .QN(n5622) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[5]  ( .D(n3577), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[37] ), 
        .QN(n5682) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[5]  ( .D(n3575), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [5])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[6]  ( .D(n3573), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5443) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[6]  ( .D(n3572), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4424) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[6]  ( .D(n3571), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4456) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[6]  ( .D(n3570), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4488) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[6]  ( .D(n3569), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4520) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[6]  ( .D(n3568), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][6] ), .QN(n4552)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[6]  ( .D(n3567), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][6] ), .QN(n4584)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[6]  ( .D(n3566), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4616) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[6]  ( .D(n3565), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4648) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[6]  ( .D(n3564), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4680) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[6]  ( .D(n3563), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4712) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[6]  ( .D(n3562), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][6] ), .QN(n4744) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[6]  ( .D(n3561), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][6] ), .QN(n4776) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[6]  ( .D(n3560), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4808) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[6]  ( .D(n3559), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4840) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[6]  ( .D(n3558), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][6] ), .QN(n4872) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[6]  ( .D(n3557), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][6] ), .QN(n4904) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[6]  ( .D(n3556), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4936) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[6]  ( .D(n3555), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4968) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[6]  ( .D(n3554), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][6] ), .QN(n5000) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[6]  ( .D(n3553), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][6] ), .QN(n5032) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[6]  ( .D(n3552), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5064) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[6]  ( .D(n3551), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][6] ), .QN(n5096) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[6]  ( .D(n3550), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][6] ), .QN(n5128) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[6]  ( .D(n3549), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5160) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[6]  ( .D(n3548), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5192) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[6]  ( .D(n3547), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5224) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[6]  ( .D(n3546), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5256) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[6]  ( .D(n3545), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5288) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[6]  ( .D(n3544), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5320) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[6]  ( .D(n3543), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5352) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[6]  ( .D(n3542), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5384) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[6]  ( .D(n3540), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[6] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[6]  ( .D(n3539), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5621) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[6]  ( .D(n3538), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[6] ), 
        .QN(n5620) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[6]  ( .D(n3537), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[38] ), 
        .QN(n5681) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[6]  ( .D(n3536), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[6] ), .QN(
        \UUT/Mpath/the_alu/N72 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[6]  ( .D(n3535), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [6])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[6]  ( .D(n3534), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [6]), .QN(
        n2682) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[7]  ( .D(n3533), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5440) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[7]  ( .D(n3532), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4423) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[7]  ( .D(n3531), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4455) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[7]  ( .D(n3530), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4487) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[7]  ( .D(n3529), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4519) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[7]  ( .D(n3528), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][7] ), .QN(n4551)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[7]  ( .D(n3527), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][7] ), .QN(n4583)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[7]  ( .D(n3526), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4615) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[7]  ( .D(n3525), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4647) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[7]  ( .D(n3524), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4679) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[7]  ( .D(n3523), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4711) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[7]  ( .D(n3522), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][7] ), .QN(n4743) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[7]  ( .D(n3521), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][7] ), .QN(n4775) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[7]  ( .D(n3520), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4807) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[7]  ( .D(n3519), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4839) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[7]  ( .D(n3518), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][7] ), .QN(n4871) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[7]  ( .D(n3517), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][7] ), .QN(n4903) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[7]  ( .D(n3516), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4935) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[7]  ( .D(n3515), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4967) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[7]  ( .D(n3514), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][7] ), .QN(n4999) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[7]  ( .D(n3513), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][7] ), .QN(n5031) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[7]  ( .D(n3512), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5063) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[7]  ( .D(n3511), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][7] ), .QN(n5095) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[7]  ( .D(n3510), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][7] ), .QN(n5127) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[7]  ( .D(n3509), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5159) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[7]  ( .D(n3508), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5191) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[7]  ( .D(n3507), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5223) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[7]  ( .D(n3506), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5255) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[7]  ( .D(n3505), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5287) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[7]  ( .D(n3504), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5319) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[7]  ( .D(n3503), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5351) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[7]  ( .D(n3502), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5383) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[7]  ( .D(n3500), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[7] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[7]  ( .D(n3499), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5619) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[7]  ( .D(n3498), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[7] ), 
        .QN(n5618) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[7]  ( .D(n3497), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[39] ), 
        .QN(n5680) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[7]  ( .D(n3496), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[7] ), .QN(
        \UUT/Mpath/the_alu/N70 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[7]  ( .D(n3495), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [7])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[7]  ( .D(n3494), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [7]), .QN(
        n2679) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[8]  ( .D(n3493), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5437) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[8]  ( .D(n3491), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[8] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[8]  ( .D(n3490), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5617) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[8]  ( .D(n3489), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[8] ), 
        .QN(n5616) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[8]  ( .D(n3488), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[40] ), 
        .QN(n5679) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[8]  ( .D(n3487), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [8]), .QN(
        n2677) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[9]  ( .D(n3486), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5433) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[9]  ( .D(n3485), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4421) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[9]  ( .D(n3484), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4453) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[9]  ( .D(n3483), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4485) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[9]  ( .D(n3482), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4517) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[9]  ( .D(n3481), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][9] ), .QN(n4549)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[9]  ( .D(n3480), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][9] ), .QN(n4581)
         );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[9]  ( .D(n3479), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4613) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[9]  ( .D(n3478), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4645) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[9]  ( .D(n3477), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4677) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[9]  ( .D(n3476), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4709) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[9]  ( .D(n3475), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][9] ), .QN(n4741) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[9]  ( .D(n3474), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][9] ), .QN(n4773) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[9]  ( .D(n3473), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4805) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[9]  ( .D(n3472), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4837) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[9]  ( .D(n3471), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][9] ), .QN(n4869) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[9]  ( .D(n3470), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][9] ), .QN(n4901) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[9]  ( .D(n3469), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4933) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[9]  ( .D(n3468), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4965) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[9]  ( .D(n3467), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][9] ), .QN(n4997) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[9]  ( .D(n3466), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][9] ), .QN(n5029) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[9]  ( .D(n3465), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5061) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[9]  ( .D(n3464), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][9] ), .QN(n5093) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[9]  ( .D(n3463), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][9] ), .QN(n5125) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[9]  ( .D(n3462), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5157) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[9]  ( .D(n3461), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5189) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[9]  ( .D(n3460), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5221) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[9]  ( .D(n3459), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5253) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[9]  ( .D(n3458), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5285) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[9]  ( .D(n3457), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5317) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[9]  ( .D(n3456), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5349) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[9]  ( .D(n3455), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5381) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[9]  ( .D(n3453), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[9] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[9]  ( .D(n3452), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5615) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[9]  ( .D(n3451), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[9] ), 
        .QN(n5614) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[9]  ( .D(n3450), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[41] ), 
        .QN(n5678) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[9]  ( .D(n3449), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[9] ), .QN(
        \UUT/Mpath/the_alu/N66 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[9]  ( .D(n3448), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [9])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[10]  ( .D(n3447), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5524) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[10]  ( .D(n3445), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[10] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[10]  ( .D(n3444), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5675) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[10]  ( .D(n3443), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[10] ), .QN(
        n5674) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[10]  ( .D(n3442), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[42] ), .QN(
        n5708) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[11]  ( .D(n3441), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5521) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[11]  ( .D(n3440), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4450) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[11]  ( .D(n3439), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4482) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[11]  ( .D(n3438), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4514) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[11]  ( .D(n3437), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4546) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[11]  ( .D(n3436), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][11] ), .QN(n4578) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[11]  ( .D(n3435), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][11] ), .QN(n4610) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[11]  ( .D(n3434), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4642) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[11]  ( .D(n3433), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4674) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[11]  ( .D(n3432), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4706) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[11]  ( .D(n3431), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4738) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[11]  ( .D(n3430), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][11] ), .QN(
        n4770) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[11]  ( .D(n3429), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][11] ), .QN(
        n4802) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[11]  ( .D(n3428), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4834) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[11]  ( .D(n3427), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4866) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[11]  ( .D(n3426), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][11] ), .QN(
        n4898) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[11]  ( .D(n3425), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][11] ), .QN(
        n4930) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[11]  ( .D(n3424), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4962) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[11]  ( .D(n3423), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4994) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[11]  ( .D(n3422), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][11] ), .QN(
        n5026) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[11]  ( .D(n3421), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][11] ), .QN(
        n5058) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[11]  ( .D(n3420), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5090) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[11]  ( .D(n3419), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][11] ), .QN(
        n5122) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[11]  ( .D(n3418), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][11] ), .QN(
        n5154) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[11]  ( .D(n3417), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5186) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[11]  ( .D(n3416), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5218) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[11]  ( .D(n3415), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5250) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[11]  ( .D(n3414), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5282) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[11]  ( .D(n3413), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5314) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[11]  ( .D(n3412), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5346) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[11]  ( .D(n3411), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5378) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[11]  ( .D(n3410), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5410) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[11]  ( .D(n3408), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[11] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[11]  ( .D(n3407), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5673) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[11]  ( .D(n3406), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[11] ), .QN(
        n5672) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[11]  ( .D(n3405), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[43] ), .QN(
        n5707) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[11]  ( .D(n3403), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [11])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[11]  ( .D(n3402), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [11]), .QN(
        n2671) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[12]  ( .D(n3401), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5518) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[12]  ( .D(n3400), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4449) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[12]  ( .D(n3399), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4481) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[12]  ( .D(n3398), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4513) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[12]  ( .D(n3397), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4545) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[12]  ( .D(n3396), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][12] ), .QN(n4577) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[12]  ( .D(n3395), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][12] ), .QN(n4609) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[12]  ( .D(n3394), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4641) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[12]  ( .D(n3393), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4673) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[12]  ( .D(n3392), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4705) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[12]  ( .D(n3391), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4737) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[12]  ( .D(n3390), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][12] ), .QN(
        n4769) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[12]  ( .D(n3389), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][12] ), .QN(
        n4801) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[12]  ( .D(n3388), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4833) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[12]  ( .D(n3387), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4865) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[12]  ( .D(n3386), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][12] ), .QN(
        n4897) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[12]  ( .D(n3385), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][12] ), .QN(
        n4929) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[12]  ( .D(n3384), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4961) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[12]  ( .D(n3383), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4993) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[12]  ( .D(n3382), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][12] ), .QN(
        n5025) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[12]  ( .D(n3381), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][12] ), .QN(
        n5057) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[12]  ( .D(n3380), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5089) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[12]  ( .D(n3379), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][12] ), .QN(
        n5121) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[12]  ( .D(n3378), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][12] ), .QN(
        n5153) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[12]  ( .D(n3377), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5185) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[12]  ( .D(n3376), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5217) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[12]  ( .D(n3375), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5249) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[12]  ( .D(n3374), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5281) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[12]  ( .D(n3373), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5313) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[12]  ( .D(n3372), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5345) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[12]  ( .D(n3371), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5377) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[12]  ( .D(n3370), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5409) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[12]  ( .D(n3368), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[12] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[12]  ( .D(n3367), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5671) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[12]  ( .D(n3366), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[12] ), .QN(
        n5670) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[12]  ( .D(n3365), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[44] ), .QN(
        n5706) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[12]  ( .D(n3363), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [12])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[12]  ( .D(n3362), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [12]), .QN(
        n2668) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[13]  ( .D(n3361), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5515) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[13]  ( .D(n3360), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4448) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[13]  ( .D(n3359), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4480) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[13]  ( .D(n3358), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4512) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[13]  ( .D(n3357), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4544) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[13]  ( .D(n3356), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][13] ), .QN(n4576) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[13]  ( .D(n3355), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][13] ), .QN(n4608) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[13]  ( .D(n3354), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4640) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[13]  ( .D(n3353), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4672) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[13]  ( .D(n3352), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4704) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[13]  ( .D(n3351), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4736) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[13]  ( .D(n3350), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][13] ), .QN(
        n4768) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[13]  ( .D(n3349), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][13] ), .QN(
        n4800) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[13]  ( .D(n3348), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4832) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[13]  ( .D(n3347), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4864) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[13]  ( .D(n3346), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][13] ), .QN(
        n4896) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[13]  ( .D(n3345), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][13] ), .QN(
        n4928) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[13]  ( .D(n3344), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4960) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[13]  ( .D(n3343), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4992) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[13]  ( .D(n3342), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][13] ), .QN(
        n5024) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[13]  ( .D(n3341), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][13] ), .QN(
        n5056) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[13]  ( .D(n3340), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5088) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[13]  ( .D(n3339), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][13] ), .QN(
        n5120) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[13]  ( .D(n3338), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][13] ), .QN(
        n5152) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[13]  ( .D(n3337), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5184) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[13]  ( .D(n3336), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5216) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[13]  ( .D(n3335), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5248) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[13]  ( .D(n3334), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5280) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[13]  ( .D(n3333), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5312) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[13]  ( .D(n3332), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5344) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[13]  ( .D(n3331), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5376) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[13]  ( .D(n3330), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5408) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[13]  ( .D(n3328), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[13] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[13]  ( .D(n3327), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5669) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[13]  ( .D(n3326), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[13] ), .QN(
        n5668) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[13]  ( .D(n3325), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[45] ), .QN(
        n5705) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[13]  ( .D(n3323), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [13]), .QN(
        n2666) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[13]  ( .D(n3322), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [13])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[14]  ( .D(n3321), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5512) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[14]  ( .D(n3320), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4447) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[14]  ( .D(n3319), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4479) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[14]  ( .D(n3318), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4511) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[14]  ( .D(n3317), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4543) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[14]  ( .D(n3316), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][14] ), .QN(n4575) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[14]  ( .D(n3315), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][14] ), .QN(n4607) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[14]  ( .D(n3314), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4639) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[14]  ( .D(n3313), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4671) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[14]  ( .D(n3312), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4703) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[14]  ( .D(n3311), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4735) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[14]  ( .D(n3310), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][14] ), .QN(
        n4767) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[14]  ( .D(n3309), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][14] ), .QN(
        n4799) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[14]  ( .D(n3308), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4831) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[14]  ( .D(n3307), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4863) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[14]  ( .D(n3306), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][14] ), .QN(
        n4895) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[14]  ( .D(n3305), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][14] ), .QN(
        n4927) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[14]  ( .D(n3304), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4959) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[14]  ( .D(n3303), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4991) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[14]  ( .D(n3302), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][14] ), .QN(
        n5023) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[14]  ( .D(n3301), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][14] ), .QN(
        n5055) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[14]  ( .D(n3300), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5087) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[14]  ( .D(n3299), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][14] ), .QN(
        n5119) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[14]  ( .D(n3298), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][14] ), .QN(
        n5151) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[14]  ( .D(n3297), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5183) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[14]  ( .D(n3296), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5215) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[14]  ( .D(n3295), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5247) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[14]  ( .D(n3294), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5279) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[14]  ( .D(n3293), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5311) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[14]  ( .D(n3292), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5343) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[14]  ( .D(n3291), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5375) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[14]  ( .D(n3290), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5407) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[14]  ( .D(n3288), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[14] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[14]  ( .D(n3287), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5667) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[14]  ( .D(n3286), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[14] ), .QN(
        n5666) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[14]  ( .D(n3285), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[46] ), .QN(
        n5704) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[14]  ( .D(n3283), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [14]), .QN(
        n2663) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[14]  ( .D(n3282), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [14])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[15]  ( .D(n3281), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5509) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[15]  ( .D(n3280), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4446) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[15]  ( .D(n3279), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4478) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[15]  ( .D(n3278), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4510) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[15]  ( .D(n3277), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4542) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[15]  ( .D(n3276), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][15] ), .QN(n4574) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[15]  ( .D(n3275), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][15] ), .QN(n4606) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[15]  ( .D(n3274), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4638) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[15]  ( .D(n3273), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4670) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[15]  ( .D(n3272), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4702) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[15]  ( .D(n3271), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4734) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[15]  ( .D(n3270), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][15] ), .QN(
        n4766) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[15]  ( .D(n3269), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][15] ), .QN(
        n4798) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[15]  ( .D(n3268), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4830) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[15]  ( .D(n3267), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4862) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[15]  ( .D(n3266), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][15] ), .QN(
        n4894) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[15]  ( .D(n3265), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][15] ), .QN(
        n4926) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[15]  ( .D(n3264), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4958) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[15]  ( .D(n3263), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4990) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[15]  ( .D(n3262), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][15] ), .QN(
        n5022) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[15]  ( .D(n3261), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][15] ), .QN(
        n5054) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[15]  ( .D(n3260), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5086) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[15]  ( .D(n3259), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][15] ), .QN(
        n5118) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[15]  ( .D(n3258), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][15] ), .QN(
        n5150) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[15]  ( .D(n3257), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5182) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[15]  ( .D(n3256), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5214) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[15]  ( .D(n3255), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5246) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[15]  ( .D(n3254), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5278) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[15]  ( .D(n3253), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5310) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[15]  ( .D(n3252), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5342) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[15]  ( .D(n3251), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5374) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[15]  ( .D(n3250), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5406) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[15]  ( .D(n3248), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[15] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[15]  ( .D(n3247), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5665) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[15]  ( .D(n3246), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[15] ), .QN(
        n5664) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[15]  ( .D(n3245), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[47] ), .QN(
        n5703) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[15]  ( .D(n3242), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [15])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[16]  ( .D(n3241), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5506) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[16]  ( .D(n3240), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4445) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[16]  ( .D(n3239), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4477) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[16]  ( .D(n3238), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4509) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[16]  ( .D(n3237), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4541) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[16]  ( .D(n3236), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][16] ), .QN(n4573) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[16]  ( .D(n3235), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][16] ), .QN(n4605) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[16]  ( .D(n3234), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4637) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[16]  ( .D(n3233), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4669) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[16]  ( .D(n3232), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4701) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[16]  ( .D(n3231), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4733) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[16]  ( .D(n3230), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][16] ), .QN(
        n4765) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[16]  ( .D(n3229), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][16] ), .QN(
        n4797) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[16]  ( .D(n3228), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4829) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[16]  ( .D(n3227), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4861) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[16]  ( .D(n3226), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][16] ), .QN(
        n4893) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[16]  ( .D(n3225), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][16] ), .QN(
        n4925) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[16]  ( .D(n3224), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4957) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[16]  ( .D(n3223), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4989) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[16]  ( .D(n3222), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][16] ), .QN(
        n5021) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[16]  ( .D(n3221), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][16] ), .QN(
        n5053) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[16]  ( .D(n3220), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5085) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[16]  ( .D(n3219), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][16] ), .QN(
        n5117) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[16]  ( .D(n3218), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][16] ), .QN(
        n5149) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[16]  ( .D(n3217), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5181) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[16]  ( .D(n3216), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5213) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[16]  ( .D(n3215), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5245) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[16]  ( .D(n3214), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5277) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[16]  ( .D(n3213), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5309) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[16]  ( .D(n3212), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5341) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[16]  ( .D(n3211), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5373) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[16]  ( .D(n3210), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5405) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[16]  ( .D(n3208), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[16] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[16]  ( .D(n3207), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5663) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[16]  ( .D(n3206), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[16] ), .QN(
        n5662) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[16]  ( .D(n3205), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[48] ), .QN(
        n5702) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[16]  ( .D(n3203), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [16]), .QN(
        n2657) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[16]  ( .D(n3202), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [16])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[17]  ( .D(n3201), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5503) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[17]  ( .D(n3200), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4444) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[17]  ( .D(n3199), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4476) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[17]  ( .D(n3198), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4508) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[17]  ( .D(n3197), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4540) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[17]  ( .D(n3196), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][17] ), .QN(n4572) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[17]  ( .D(n3195), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][17] ), .QN(n4604) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[17]  ( .D(n3194), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4636) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[17]  ( .D(n3193), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4668) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[17]  ( .D(n3192), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4700) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[17]  ( .D(n3191), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4732) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[17]  ( .D(n3190), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][17] ), .QN(
        n4764) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[17]  ( .D(n3189), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][17] ), .QN(
        n4796) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[17]  ( .D(n3188), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4828) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[17]  ( .D(n3187), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4860) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[17]  ( .D(n3186), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][17] ), .QN(
        n4892) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[17]  ( .D(n3185), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][17] ), .QN(
        n4924) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[17]  ( .D(n3184), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4956) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[17]  ( .D(n3183), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4988) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[17]  ( .D(n3182), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][17] ), .QN(
        n5020) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[17]  ( .D(n3181), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][17] ), .QN(
        n5052) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[17]  ( .D(n3180), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5084) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[17]  ( .D(n3179), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][17] ), .QN(
        n5116) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[17]  ( .D(n3178), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][17] ), .QN(
        n5148) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[17]  ( .D(n3177), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5180) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[17]  ( .D(n3176), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5212) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[17]  ( .D(n3175), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5244) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[17]  ( .D(n3174), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5276) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[17]  ( .D(n3173), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5308) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[17]  ( .D(n3172), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5340) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[17]  ( .D(n3171), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5372) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[17]  ( .D(n3170), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5404) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[17]  ( .D(n3168), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[17] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[17]  ( .D(n3167), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5661) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[17]  ( .D(n3166), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[17] ), .QN(
        n5660) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[17]  ( .D(n3165), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[49] ), .QN(
        n5701) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[17]  ( .D(n3163), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [17]), .QN(
        n2654) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[17]  ( .D(n3162), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [17])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[18]  ( .D(n3161), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5500) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[18]  ( .D(n3160), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4443) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[18]  ( .D(n3159), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4475) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[18]  ( .D(n3158), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4507) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[18]  ( .D(n3157), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4539) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[18]  ( .D(n3156), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][18] ), .QN(n4571) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[18]  ( .D(n3155), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][18] ), .QN(n4603) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[18]  ( .D(n3154), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4635) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[18]  ( .D(n3153), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4667) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[18]  ( .D(n3152), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4699) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[18]  ( .D(n3151), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4731) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[18]  ( .D(n3150), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][18] ), .QN(
        n4763) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[18]  ( .D(n3149), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][18] ), .QN(
        n4795) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[18]  ( .D(n3148), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4827) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[18]  ( .D(n3147), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4859) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[18]  ( .D(n3146), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][18] ), .QN(
        n4891) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[18]  ( .D(n3145), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][18] ), .QN(
        n4923) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[18]  ( .D(n3144), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4955) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[18]  ( .D(n3143), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4987) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[18]  ( .D(n3142), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][18] ), .QN(
        n5019) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[18]  ( .D(n3141), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][18] ), .QN(
        n5051) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[18]  ( .D(n3140), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5083) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[18]  ( .D(n3139), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][18] ), .QN(
        n5115) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[18]  ( .D(n3138), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][18] ), .QN(
        n5147) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[18]  ( .D(n3137), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5179) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[18]  ( .D(n3136), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5211) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[18]  ( .D(n3135), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5243) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[18]  ( .D(n3134), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5275) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[18]  ( .D(n3133), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5307) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[18]  ( .D(n3132), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5339) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[18]  ( .D(n3131), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5371) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[18]  ( .D(n3130), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5403) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[18]  ( .D(n3128), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[18] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[18]  ( .D(n3127), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5659) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[18]  ( .D(n3126), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[18] ), .QN(
        n5658) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[18]  ( .D(n3125), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[50] ), .QN(
        n5700) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[18]  ( .D(n3122), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [18])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[19]  ( .D(n3121), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5497) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[19]  ( .D(n3120), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4442) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[19]  ( .D(n3119), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4474) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[19]  ( .D(n3118), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4506) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[19]  ( .D(n3117), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4538) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[19]  ( .D(n3116), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][19] ), .QN(n4570) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[19]  ( .D(n3115), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][19] ), .QN(n4602) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[19]  ( .D(n3114), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4634) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[19]  ( .D(n3113), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4666) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[19]  ( .D(n3112), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4698) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[19]  ( .D(n3111), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4730) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[19]  ( .D(n3110), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][19] ), .QN(
        n4762) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[19]  ( .D(n3109), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][19] ), .QN(
        n4794) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[19]  ( .D(n3108), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4826) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[19]  ( .D(n3107), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4858) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[19]  ( .D(n3106), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][19] ), .QN(
        n4890) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[19]  ( .D(n3105), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][19] ), .QN(
        n4922) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[19]  ( .D(n3104), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4954) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[19]  ( .D(n3103), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4986) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[19]  ( .D(n3102), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][19] ), .QN(
        n5018) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[19]  ( .D(n3101), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][19] ), .QN(
        n5050) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[19]  ( .D(n3100), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5082) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[19]  ( .D(n3099), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][19] ), .QN(
        n5114) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[19]  ( .D(n3098), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][19] ), .QN(
        n5146) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[19]  ( .D(n3097), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5178) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[19]  ( .D(n3096), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5210) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[19]  ( .D(n3095), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5242) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[19]  ( .D(n3094), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5274) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[19]  ( .D(n3093), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5306) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[19]  ( .D(n3092), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5338) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[19]  ( .D(n3091), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5370) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[19]  ( .D(n3090), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5402) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[19]  ( .D(n3088), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[19] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[19]  ( .D(n3087), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5657) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[19]  ( .D(n3086), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[19] ), .QN(
        n5656) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[19]  ( .D(n3085), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[51] ), .QN(
        n5699) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[19]  ( .D(n3083), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [19]), .QN(
        n2648) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[19]  ( .D(n3082), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [19])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[20]  ( .D(n3081), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5491) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[20]  ( .D(n3080), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4440) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[20]  ( .D(n3079), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4472) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[20]  ( .D(n3078), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4504) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[20]  ( .D(n3077), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4536) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[20]  ( .D(n3076), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][20] ), .QN(n4568) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[20]  ( .D(n3075), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][20] ), .QN(n4600) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[20]  ( .D(n3074), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4632) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[20]  ( .D(n3073), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4664) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[20]  ( .D(n3072), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4696) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[20]  ( .D(n3071), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4728) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[20]  ( .D(n3070), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][20] ), .QN(
        n4760) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[20]  ( .D(n3069), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][20] ), .QN(
        n4792) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[20]  ( .D(n3068), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4824) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[20]  ( .D(n3067), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4856) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[20]  ( .D(n3066), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][20] ), .QN(
        n4888) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[20]  ( .D(n3065), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][20] ), .QN(
        n4920) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[20]  ( .D(n3064), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4952) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[20]  ( .D(n3063), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4984) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[20]  ( .D(n3062), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][20] ), .QN(
        n5016) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[20]  ( .D(n3061), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][20] ), .QN(
        n5048) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[20]  ( .D(n3060), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5080) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[20]  ( .D(n3059), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][20] ), .QN(
        n5112) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[20]  ( .D(n3058), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][20] ), .QN(
        n5144) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[20]  ( .D(n3057), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5176) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[20]  ( .D(n3056), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5208) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[20]  ( .D(n3055), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5240) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[20]  ( .D(n3054), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5272) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[20]  ( .D(n3053), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5304) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[20]  ( .D(n3052), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5336) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[20]  ( .D(n3051), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5368) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[20]  ( .D(n3050), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5400) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[20]  ( .D(n3048), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[20] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[20]  ( .D(n3047), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5653) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[20]  ( .D(n3046), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[20] ), .QN(
        n5652) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[20]  ( .D(n3045), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[52] ), .QN(
        n5697) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[20]  ( .D(n3043), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [20]), .QN(
        n2645) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[20]  ( .D(n3042), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [20])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[21]  ( .D(n3041), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5488) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[21]  ( .D(n3040), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4439) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[21]  ( .D(n3039), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4471) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[21]  ( .D(n3038), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4503) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[21]  ( .D(n3037), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4535) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[21]  ( .D(n3036), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][21] ), .QN(n4567) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[21]  ( .D(n3035), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][21] ), .QN(n4599) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[21]  ( .D(n3034), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4631) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[21]  ( .D(n3033), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4663) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[21]  ( .D(n3032), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4695) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[21]  ( .D(n3031), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4727) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[21]  ( .D(n3030), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][21] ), .QN(
        n4759) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[21]  ( .D(n3029), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][21] ), .QN(
        n4791) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[21]  ( .D(n3028), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4823) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[21]  ( .D(n3027), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4855) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[21]  ( .D(n3026), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][21] ), .QN(
        n4887) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[21]  ( .D(n3025), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][21] ), .QN(
        n4919) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[21]  ( .D(n3024), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4951) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[21]  ( .D(n3023), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4983) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[21]  ( .D(n3022), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][21] ), .QN(
        n5015) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[21]  ( .D(n3021), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][21] ), .QN(
        n5047) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[21]  ( .D(n3020), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5079) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[21]  ( .D(n3019), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][21] ), .QN(
        n5111) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[21]  ( .D(n3018), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][21] ), .QN(
        n5143) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[21]  ( .D(n3017), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5175) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[21]  ( .D(n3016), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5207) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[21]  ( .D(n3015), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5239) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[21]  ( .D(n3014), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5271) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[21]  ( .D(n3013), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5303) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[21]  ( .D(n3012), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5335) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[21]  ( .D(n3011), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5367) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[21]  ( .D(n3010), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5399) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[21]  ( .D(n3008), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[21] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[21]  ( .D(n3007), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5651) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[21]  ( .D(n3006), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[21] ), .QN(
        n5650) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[21]  ( .D(n3005), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[53] ), .QN(
        n5696) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[21]  ( .D(n3003), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [21]), .QN(
        n2642) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[21]  ( .D(n3002), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [21])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[22]  ( .D(n3001), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5485) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[22]  ( .D(n3000), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4438) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[22]  ( .D(n2999), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4470) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[22]  ( .D(n2998), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4502) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[22]  ( .D(n2997), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4534) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[22]  ( .D(n2996), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][22] ), .QN(n4566) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[22]  ( .D(n2995), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][22] ), .QN(n4598) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[22]  ( .D(n2994), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4630) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[22]  ( .D(n2993), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4662) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[22]  ( .D(n2992), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4694) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[22]  ( .D(n2991), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4726) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[22]  ( .D(n2990), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][22] ), .QN(
        n4758) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[22]  ( .D(n2989), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][22] ), .QN(
        n4790) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[22]  ( .D(n2988), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4822) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[22]  ( .D(n2987), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4854) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[22]  ( .D(n2986), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][22] ), .QN(
        n4886) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[22]  ( .D(n2985), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][22] ), .QN(
        n4918) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[22]  ( .D(n2984), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4950) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[22]  ( .D(n2983), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4982) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[22]  ( .D(n2982), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][22] ), .QN(
        n5014) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[22]  ( .D(n2981), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][22] ), .QN(
        n5046) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[22]  ( .D(n2980), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5078) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[22]  ( .D(n2979), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][22] ), .QN(
        n5110) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[22]  ( .D(n2978), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][22] ), .QN(
        n5142) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[22]  ( .D(n2977), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5174) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[22]  ( .D(n2976), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5206) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[22]  ( .D(n2975), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5238) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[22]  ( .D(n2974), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5270) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[22]  ( .D(n2973), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5302) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[22]  ( .D(n2972), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5334) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[22]  ( .D(n2971), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5366) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[22]  ( .D(n2970), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5398) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[22]  ( .D(n2968), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[22] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[22]  ( .D(n2967), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5649) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[22]  ( .D(n2966), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[22] ), .QN(
        n5648) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[22]  ( .D(n2965), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[54] ), .QN(
        n5695) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[22]  ( .D(n2963), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [22]), .QN(
        n2639) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[22]  ( .D(n2962), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [22])
         );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[24]  ( .D(n2961), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5479) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[24]  ( .D(n2960), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4436) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[24]  ( .D(n2959), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4468) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[24]  ( .D(n2958), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4500) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[24]  ( .D(n2957), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4532) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[24]  ( .D(n2956), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][24] ), .QN(n4564) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[24]  ( .D(n2955), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][24] ), .QN(n4596) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[24]  ( .D(n2954), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4628) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[24]  ( .D(n2953), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4660) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[24]  ( .D(n2952), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4692) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[24]  ( .D(n2951), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4724) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[24]  ( .D(n2950), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][24] ), .QN(
        n4756) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[24]  ( .D(n2949), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][24] ), .QN(
        n4788) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[24]  ( .D(n2948), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4820) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[24]  ( .D(n2947), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4852) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[24]  ( .D(n2946), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][24] ), .QN(
        n4884) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[24]  ( .D(n2945), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][24] ), .QN(
        n4916) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[24]  ( .D(n2944), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4948) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[24]  ( .D(n2943), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4980) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[24]  ( .D(n2942), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][24] ), .QN(
        n5012) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[24]  ( .D(n2941), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][24] ), .QN(
        n5044) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[24]  ( .D(n2940), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5076) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[24]  ( .D(n2939), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][24] ), .QN(
        n5108) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[24]  ( .D(n2938), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][24] ), .QN(
        n5140) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[24]  ( .D(n2937), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5172) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[24]  ( .D(n2936), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5204) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[24]  ( .D(n2935), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5236) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[24]  ( .D(n2934), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5268) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[24]  ( .D(n2933), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5300) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[24]  ( .D(n2932), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5332) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[24]  ( .D(n2931), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5364) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[24]  ( .D(n2930), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5396) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[24]  ( .D(n2928), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[24] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[24]  ( .D(n2927), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5645) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[24]  ( .D(n2926), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[24] ), .QN(
        n5644) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[24]  ( .D(n2925), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[56] ), .QN(
        n5693) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[24]  ( .D(n2923), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [24])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[25]  ( .D(n2922), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[25] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[25]  ( .D(n2921), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5643) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[25]  ( .D(n2920), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[25] ), .QN(
        n5642) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[25]  ( .D(n2919), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[57] ), .QN(
        n5692) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[25]  ( .D(n2917), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [25])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[26]  ( .D(n2916), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[26] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[26]  ( .D(n2915), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5641) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[26]  ( .D(n2914), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[26] ), .QN(
        n5640) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[26]  ( .D(n2913), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[58] ), .QN(
        n5691) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[26]  ( .D(n2911), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [26])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[27]  ( .D(n2910), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[27] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[27]  ( .D(n2909), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5639) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[27]  ( .D(n2908), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[27] ), .QN(
        n5638) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[27]  ( .D(n2907), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[59] ), .QN(
        n5690) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[27]  ( .D(n2905), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [27])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[28]  ( .D(n2904), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[28] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[28]  ( .D(n2903), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5637) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[28]  ( .D(n2902), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[28] ), .QN(
        n5636) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[28]  ( .D(n2901), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[60] ), .QN(
        n5689) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[28]  ( .D(n2899), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [28])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[29]  ( .D(n2898), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[29] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[29]  ( .D(n2897), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n5635) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[29]  ( .D(n2896), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[29] ), .QN(
        n5634) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[29]  ( .D(n2895), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[61] ), .QN(
        n5688) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[29]  ( .D(n2894), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[29] ), .QN(
        \UUT/Mpath/the_alu/N26 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[29]  ( .D(n2893), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [29])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[30]  ( .D(n2892), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [30])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[23]  ( .D(n2891), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [23])
         );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[31]  ( .D(n2890), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[31] ), 
        .QN(n2623) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[30]  ( .D(n2889), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[30] ), 
        .QN(n2622) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[29]  ( .D(n2888), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[29] ), 
        .QN(n2621) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[28]  ( .D(n2887), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[28] ), 
        .QN(n2620) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[27]  ( .D(n2886), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[27] ), 
        .QN(n2619) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[26]  ( .D(n2885), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[26] ), 
        .QN(n2618) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[25]  ( .D(n2884), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[25] ), 
        .QN(n2617) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[24]  ( .D(n2883), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[24] ), 
        .QN(n2616) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[23]  ( .D(n2882), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[23] ), 
        .QN(n2615) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[22]  ( .D(n2881), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[22] ), 
        .QN(n2614) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[21]  ( .D(n2880), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[21] ), 
        .QN(n2613) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[20]  ( .D(n2879), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[20] ), 
        .QN(n2612) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[19]  ( .D(n2878), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[19] ), 
        .QN(n2611) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[18]  ( .D(n2877), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[18] ), 
        .QN(n2610) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[17]  ( .D(n2876), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[17] ), 
        .QN(n2609) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[16]  ( .D(n2875), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[16] ), 
        .QN(n2608) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[15]  ( .D(n2874), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
        .QN(n2607) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[14]  ( .D(n2873), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
        .QN(n2606) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[13]  ( .D(n2872), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
        .QN(n2605) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[12]  ( .D(n2871), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
        .QN(n2604) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[11]  ( .D(n2870), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
        .QN(n2603) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[10]  ( .D(n2869), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
        .QN(n2602) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[9]  ( .D(n2868), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_memhandle/smdr_out[9] ), .QN(n2601) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[8]  ( .D(n2867), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_memhandle/smdr_out[8] ), .QN(n2600) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[7]  ( .D(n2866), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[7]), .QN(n4380) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[6]  ( .D(n2865), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[6]), .QN(n4381) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[5]  ( .D(n2864), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[5]), .QN(n4382) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[4]  ( .D(n2863), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[4]), .QN(n4383) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[3]  ( .D(n2862), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[3]), .QN(n4384) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[2]  ( .D(n2861), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[2]), .QN(n4387) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[1]  ( .D(n2860), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[1]), .QN(n4398) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[0]  ( .D(n2859), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[0]), .QN(n4409) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[8]  ( .D(n2858), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [8])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[10]  ( .D(n2857), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [10])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[31]  ( .D(n2856), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [31])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[0]  ( .D(n2855), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [0])
         );
  OAI221_X1 U3 ( .B1(n68), .B2(n69), .C1(n70), .C2(n71), .A(n72), .ZN(n2855)
         );
  NAND2_X1 U4 ( .A1(\UUT/Mpath/the_mult/x_operand2 [0]), .A2(n6409), .ZN(n72)
         );
  OAI21_X1 U5 ( .B1(n74), .B2(n6409), .A(n75), .ZN(n2856) );
  NAND2_X1 U6 ( .A1(\UUT/Mpath/the_mult/x_operand2 [31]), .A2(n6409), .ZN(n75)
         );
  OAI221_X1 U7 ( .B1(n76), .B2(n69), .C1(n77), .C2(n71), .A(n78), .ZN(n2857)
         );
  NAND2_X1 U8 ( .A1(\UUT/Mpath/the_mult/x_operand2 [10]), .A2(n6409), .ZN(n78)
         );
  OAI221_X1 U9 ( .B1(n79), .B2(n69), .C1(n80), .C2(n71), .A(n81), .ZN(n2858)
         );
  NAND2_X1 U10 ( .A1(\UUT/Mpath/the_mult/x_operand2 [8]), .A2(n6409), .ZN(n81)
         );
  OAI22_X1 U11 ( .A1(n4409), .A2(n82), .B1(n70), .B2(n83), .ZN(n2859) );
  OAI22_X1 U12 ( .A1(n4398), .A2(n82), .B1(n84), .B2(n83), .ZN(n2860) );
  OAI22_X1 U13 ( .A1(n4387), .A2(n82), .B1(n85), .B2(n83), .ZN(n2861) );
  OAI22_X1 U14 ( .A1(n4384), .A2(n82), .B1(n86), .B2(n83), .ZN(n2862) );
  OAI22_X1 U15 ( .A1(n4383), .A2(n82), .B1(n87), .B2(n83), .ZN(n2863) );
  OAI22_X1 U16 ( .A1(n4382), .A2(n82), .B1(n88), .B2(n83), .ZN(n2864) );
  OAI22_X1 U48 ( .A1(n4381), .A2(n82), .B1(n89), .B2(n83), .ZN(n2865) );
  OAI22_X1 U49 ( .A1(n4380), .A2(n82), .B1(n90), .B2(n83), .ZN(n2866) );
  OAI22_X1 U50 ( .A1(n82), .A2(n2600), .B1(n80), .B2(n83), .ZN(n2867) );
  OAI22_X1 U51 ( .A1(n82), .A2(n2601), .B1(n91), .B2(n83), .ZN(n2868) );
  OAI22_X1 U52 ( .A1(n82), .A2(n2602), .B1(n77), .B2(n83), .ZN(n2869) );
  OAI22_X1 U53 ( .A1(n82), .A2(n2603), .B1(n92), .B2(n83), .ZN(n2870) );
  OAI22_X1 U54 ( .A1(n82), .A2(n2604), .B1(n93), .B2(n83), .ZN(n2871) );
  OAI22_X1 U55 ( .A1(n82), .A2(n2605), .B1(n94), .B2(n83), .ZN(n2872) );
  OAI22_X1 U56 ( .A1(n82), .A2(n2606), .B1(n95), .B2(n83), .ZN(n2873) );
  OAI22_X1 U57 ( .A1(n82), .A2(n2607), .B1(n96), .B2(n83), .ZN(n2874) );
  OAI22_X1 U58 ( .A1(n82), .A2(n2608), .B1(n97), .B2(n83), .ZN(n2875) );
  OAI22_X1 U59 ( .A1(n82), .A2(n2609), .B1(n98), .B2(n83), .ZN(n2876) );
  OAI22_X1 U60 ( .A1(n82), .A2(n2610), .B1(n99), .B2(n83), .ZN(n2877) );
  OAI22_X1 U61 ( .A1(n82), .A2(n2611), .B1(n100), .B2(n83), .ZN(n2878) );
  OAI22_X1 U62 ( .A1(n82), .A2(n2612), .B1(n101), .B2(n83), .ZN(n2879) );
  OAI22_X1 U63 ( .A1(n82), .A2(n2613), .B1(n102), .B2(n83), .ZN(n2880) );
  OAI22_X1 U64 ( .A1(n82), .A2(n2614), .B1(n103), .B2(n83), .ZN(n2881) );
  OAI22_X1 U65 ( .A1(n82), .A2(n2615), .B1(n104), .B2(n83), .ZN(n2882) );
  OAI22_X1 U66 ( .A1(n82), .A2(n2616), .B1(n105), .B2(n83), .ZN(n2883) );
  INV_X1 U67 ( .A(n106), .ZN(n105) );
  OAI22_X1 U68 ( .A1(n82), .A2(n2617), .B1(n107), .B2(n83), .ZN(n2884) );
  INV_X1 U69 ( .A(n108), .ZN(n107) );
  OAI22_X1 U70 ( .A1(n82), .A2(n2618), .B1(n109), .B2(n83), .ZN(n2885) );
  INV_X1 U71 ( .A(n110), .ZN(n109) );
  OAI22_X1 U72 ( .A1(n82), .A2(n2619), .B1(n111), .B2(n83), .ZN(n2886) );
  OAI22_X1 U73 ( .A1(n82), .A2(n2620), .B1(n112), .B2(n83), .ZN(n2887) );
  OAI22_X1 U74 ( .A1(n82), .A2(n2621), .B1(n113), .B2(n83), .ZN(n2888) );
  OAI22_X1 U75 ( .A1(n82), .A2(n2622), .B1(n114), .B2(n83), .ZN(n2889) );
  OAI22_X1 U76 ( .A1(n82), .A2(n2623), .B1(n115), .B2(n83), .ZN(n2890) );
  OAI221_X1 U79 ( .B1(n117), .B2(n69), .C1(n104), .C2(n71), .A(n118), .ZN(
        n2891) );
  NAND2_X1 U80 ( .A1(\UUT/Mpath/the_mult/x_operand2 [23]), .A2(n6409), .ZN(
        n118) );
  OAI221_X1 U81 ( .B1(n119), .B2(n6409), .C1(n114), .C2(n71), .A(n120), .ZN(
        n2892) );
  NAND2_X1 U82 ( .A1(\UUT/Mpath/the_mult/x_operand2 [30]), .A2(n6409), .ZN(
        n120) );
  OAI221_X1 U83 ( .B1(n121), .B2(n6409), .C1(n113), .C2(n71), .A(n122), .ZN(
        n2893) );
  NAND2_X1 U84 ( .A1(\UUT/Mpath/the_mult/x_operand2 [29]), .A2(n6409), .ZN(
        n122) );
  OAI222_X1 U85 ( .A1(n113), .A2(n123), .B1(net54933), .B2(n121), .C1(
        \UUT/Mpath/the_alu/N26 ), .C2(net54893), .ZN(n2894) );
  AOI21_X1 U86 ( .B1(\UUT/Mcontrol/d_sampled_finstr [13]), .B2(n125), .A(n126), 
        .ZN(n121) );
  INV_X1 U87 ( .A(n127), .ZN(n113) );
  OAI222_X1 U88 ( .A1(n128), .A2(n129), .B1(n130), .B2(n131), .C1(n5463), .C2(
        n132), .ZN(n127) );
  OAI221_X1 U91 ( .B1(n140), .B2(n141), .C1(n5634), .C2(n142), .A(n143), .ZN(
        n2896) );
  AOI22_X1 U92 ( .A1(n144), .A2(n138), .B1(\UUT/Mpath/the_mult/Mad_out [29]), 
        .B2(n145), .ZN(n143) );
  INV_X1 U93 ( .A(n5635), .ZN(n138) );
  OAI22_X1 U94 ( .A1(net54903), .A2(n146), .B1(n5635), .B2(net54873), .ZN(
        n2897) );
  OAI22_X1 U95 ( .A1(n147), .A2(n146), .B1(n148), .B2(n6409), .ZN(n2898) );
  INV_X1 U96 ( .A(\UUT/Mpath/the_mult/x_operand1[29] ), .ZN(n146) );
  OAI221_X1 U97 ( .B1(n149), .B2(n6409), .C1(n112), .C2(n71), .A(n150), .ZN(
        n2899) );
  NAND2_X1 U98 ( .A1(\UUT/Mpath/the_mult/x_operand2 [28]), .A2(n6409), .ZN(
        n150) );
  OAI222_X1 U99 ( .A1(n112), .A2(n123), .B1(net54933), .B2(n149), .C1(
        \UUT/Mpath/the_alu/N28 ), .C2(net54893), .ZN(n2900) );
  AOI21_X1 U100 ( .B1(\UUT/Mcontrol/d_sampled_finstr [12]), .B2(n125), .A(n126), .ZN(n149) );
  INV_X1 U101 ( .A(n151), .ZN(n112) );
  OAI222_X1 U102 ( .A1(n152), .A2(n129), .B1(n153), .B2(n131), .C1(n5466), 
        .C2(n132), .ZN(n151) );
  OAI221_X1 U105 ( .B1(n140), .B2(n157), .C1(n5636), .C2(n142), .A(n158), .ZN(
        n2902) );
  AOI22_X1 U106 ( .A1(n144), .A2(n156), .B1(\UUT/Mpath/the_mult/Mad_out [28]), 
        .B2(n145), .ZN(n158) );
  INV_X1 U107 ( .A(n5637), .ZN(n156) );
  OAI22_X1 U108 ( .A1(net54905), .A2(n159), .B1(n5637), .B2(net54875), .ZN(
        n2903) );
  OAI22_X1 U109 ( .A1(n147), .A2(n159), .B1(n160), .B2(n6409), .ZN(n2904) );
  INV_X1 U110 ( .A(\UUT/Mpath/the_mult/x_operand1[28] ), .ZN(n159) );
  OAI221_X1 U111 ( .B1(n161), .B2(n6409), .C1(n111), .C2(n71), .A(n162), .ZN(
        n2905) );
  NAND2_X1 U112 ( .A1(\UUT/Mpath/the_mult/x_operand2 [27]), .A2(n6409), .ZN(
        n162) );
  OAI222_X1 U113 ( .A1(n111), .A2(n123), .B1(net54933), .B2(n161), .C1(
        \UUT/Mpath/the_alu/N30 ), .C2(net54893), .ZN(n2906) );
  AOI21_X1 U114 ( .B1(\UUT/Mcontrol/d_sampled_finstr [11]), .B2(n125), .A(n126), .ZN(n161) );
  INV_X1 U115 ( .A(n163), .ZN(n111) );
  OAI222_X1 U116 ( .A1(n164), .A2(n129), .B1(n165), .B2(n131), .C1(n5469), 
        .C2(n132), .ZN(n163) );
  OAI221_X1 U117 ( .B1(n133), .B2(n166), .C1(n5690), .C2(n135), .A(n167), .ZN(
        n2907) );
  AOI22_X1 U118 ( .A1(n137), .A2(n168), .B1(\UUT/Mpath/the_mult/Mad_out [59]), 
        .B2(n139), .ZN(n167) );
  OAI221_X1 U119 ( .B1(n140), .B2(n169), .C1(n5638), .C2(n142), .A(n170), .ZN(
        n2908) );
  AOI22_X1 U120 ( .A1(n144), .A2(n168), .B1(\UUT/Mpath/the_mult/Mad_out [27]), 
        .B2(n145), .ZN(n170) );
  INV_X1 U121 ( .A(n5639), .ZN(n168) );
  OAI22_X1 U122 ( .A1(net54903), .A2(n171), .B1(n5639), .B2(net54875), .ZN(
        n2909) );
  OAI22_X1 U123 ( .A1(n147), .A2(n171), .B1(n172), .B2(n6409), .ZN(n2910) );
  INV_X1 U124 ( .A(\UUT/Mpath/the_mult/x_operand1[27] ), .ZN(n171) );
  OAI21_X1 U125 ( .B1(n173), .B2(n6409), .A(n174), .ZN(n2911) );
  NAND2_X1 U126 ( .A1(\UUT/Mpath/the_mult/x_operand2 [26]), .A2(n6409), .ZN(
        n174) );
  OAI22_X1 U127 ( .A1(\UUT/Mpath/the_alu/N32 ), .A2(net54879), .B1(net54919), 
        .B2(n173), .ZN(n2912) );
  AOI211_X1 U128 ( .C1(n175), .C2(n110), .A(n176), .B(n177), .ZN(n173) );
  INV_X1 U129 ( .A(n178), .ZN(n177) );
  AOI22_X1 U130 ( .A1(n179), .A2(\UUT/Mcontrol/d_sampled_finstr [24]), .B1(
        n125), .B2(\UUT/Mcontrol/d_sampled_finstr [10]), .ZN(n178) );
  OAI222_X1 U131 ( .A1(n180), .A2(n129), .B1(n181), .B2(n131), .C1(n5472), 
        .C2(n132), .ZN(n110) );
  OAI221_X1 U132 ( .B1(n133), .B2(n182), .C1(n5691), .C2(n135), .A(n183), .ZN(
        n2913) );
  AOI22_X1 U133 ( .A1(n137), .A2(n184), .B1(\UUT/Mpath/the_mult/Mad_out [58]), 
        .B2(n139), .ZN(n183) );
  OAI221_X1 U134 ( .B1(n140), .B2(n185), .C1(n5640), .C2(n142), .A(n186), .ZN(
        n2914) );
  AOI22_X1 U135 ( .A1(n144), .A2(n184), .B1(\UUT/Mpath/the_mult/Mad_out [26]), 
        .B2(n145), .ZN(n186) );
  INV_X1 U136 ( .A(n5641), .ZN(n184) );
  OAI22_X1 U137 ( .A1(net54907), .A2(n187), .B1(n5641), .B2(net54873), .ZN(
        n2915) );
  OAI22_X1 U138 ( .A1(n147), .A2(n187), .B1(n188), .B2(n6409), .ZN(n2916) );
  INV_X1 U139 ( .A(\UUT/Mpath/the_mult/x_operand1[26] ), .ZN(n187) );
  OAI21_X1 U140 ( .B1(n189), .B2(n6409), .A(n190), .ZN(n2917) );
  NAND2_X1 U141 ( .A1(\UUT/Mpath/the_mult/x_operand2 [25]), .A2(n6409), .ZN(
        n190) );
  OAI22_X1 U142 ( .A1(\UUT/Mpath/the_alu/N34 ), .A2(net54879), .B1(net54919), 
        .B2(n189), .ZN(n2918) );
  AOI211_X1 U143 ( .C1(n175), .C2(n108), .A(n176), .B(n191), .ZN(n189) );
  INV_X1 U144 ( .A(n192), .ZN(n191) );
  AOI22_X1 U145 ( .A1(n179), .A2(\UUT/Mcontrol/d_sampled_finstr [23]), .B1(
        n125), .B2(\UUT/Mcontrol/d_sampled_finstr [9]), .ZN(n192) );
  OAI222_X1 U146 ( .A1(n193), .A2(n129), .B1(n194), .B2(n131), .C1(n5475), 
        .C2(n132), .ZN(n108) );
  OAI221_X1 U147 ( .B1(n133), .B2(n195), .C1(n5692), .C2(n135), .A(n196), .ZN(
        n2919) );
  AOI22_X1 U148 ( .A1(n137), .A2(n197), .B1(\UUT/Mpath/the_mult/Mad_out [57]), 
        .B2(n139), .ZN(n196) );
  OAI221_X1 U149 ( .B1(n140), .B2(n198), .C1(n5642), .C2(n142), .A(n199), .ZN(
        n2920) );
  AOI22_X1 U150 ( .A1(n144), .A2(n197), .B1(\UUT/Mpath/the_mult/Mad_out [25]), 
        .B2(n145), .ZN(n199) );
  INV_X1 U151 ( .A(n5643), .ZN(n197) );
  OAI22_X1 U152 ( .A1(net54905), .A2(n200), .B1(n5643), .B2(net54875), .ZN(
        n2921) );
  OAI22_X1 U153 ( .A1(n147), .A2(n200), .B1(n201), .B2(n6409), .ZN(n2922) );
  INV_X1 U154 ( .A(\UUT/Mpath/the_mult/x_operand1[25] ), .ZN(n200) );
  OAI21_X1 U155 ( .B1(n202), .B2(n6409), .A(n203), .ZN(n2923) );
  NAND2_X1 U156 ( .A1(\UUT/Mpath/the_mult/x_operand2 [24]), .A2(n6409), .ZN(
        n203) );
  OAI22_X1 U157 ( .A1(\UUT/Mpath/the_alu/N36 ), .A2(net54879), .B1(net54923), 
        .B2(n202), .ZN(n2924) );
  AOI211_X1 U158 ( .C1(n175), .C2(n106), .A(n176), .B(n204), .ZN(n202) );
  INV_X1 U159 ( .A(n205), .ZN(n204) );
  AOI22_X1 U160 ( .A1(n179), .A2(\UUT/Mcontrol/d_sampled_finstr [22]), .B1(
        n125), .B2(\UUT/Mcontrol/d_sampled_finstr [8]), .ZN(n205) );
  NOR2_X1 U161 ( .A1(n206), .A2(n5872), .ZN(n179) );
  INV_X1 U162 ( .A(n207), .ZN(n206) );
  OAI222_X1 U163 ( .A1(n208), .A2(n129), .B1(n209), .B2(n131), .C1(n5478), 
        .C2(n132), .ZN(n106) );
  OAI221_X1 U164 ( .B1(n133), .B2(n210), .C1(n5693), .C2(n135), .A(n211), .ZN(
        n2925) );
  AOI22_X1 U165 ( .A1(n137), .A2(n212), .B1(\UUT/Mpath/the_mult/Mad_out [56]), 
        .B2(n139), .ZN(n211) );
  OAI221_X1 U166 ( .B1(n140), .B2(n213), .C1(n5644), .C2(n142), .A(n214), .ZN(
        n2926) );
  AOI22_X1 U167 ( .A1(n144), .A2(n212), .B1(\UUT/Mpath/the_mult/Mad_out [24]), 
        .B2(n145), .ZN(n214) );
  INV_X1 U168 ( .A(n5645), .ZN(n212) );
  OAI22_X1 U169 ( .A1(net54905), .A2(n215), .B1(n5645), .B2(net54875), .ZN(
        n2927) );
  OAI22_X1 U170 ( .A1(n147), .A2(n215), .B1(n216), .B2(n6409), .ZN(n2928) );
  INV_X1 U171 ( .A(\UUT/Mpath/the_mult/x_operand1[24] ), .ZN(n215) );
  OAI22_X1 U172 ( .A1(\UUT/Mpath/the_alu/N35 ), .A2(net54879), .B1(net54919), 
        .B2(n216), .ZN(n2929) );
  INV_X1 U173 ( .A(n217), .ZN(n216) );
  OAI222_X1 U174 ( .A1(n5530), .A2(n209), .B1(n5528), .B2(n208), .C1(n6364), 
        .C2(n5421), .ZN(n217) );
  OAI22_X1 U175 ( .A1(n5396), .A2(n6407), .B1(n209), .B2(n219), .ZN(n2930) );
  OAI22_X1 U176 ( .A1(n5364), .A2(n6410), .B1(n209), .B2(n221), .ZN(n2931) );
  OAI22_X1 U177 ( .A1(n5332), .A2(n6401), .B1(n209), .B2(n223), .ZN(n2932) );
  OAI22_X1 U178 ( .A1(n5300), .A2(n6406), .B1(n209), .B2(n225), .ZN(n2933) );
  OAI22_X1 U179 ( .A1(n5268), .A2(n6399), .B1(n209), .B2(n227), .ZN(n2934) );
  OAI22_X1 U180 ( .A1(n5236), .A2(n6404), .B1(n209), .B2(n229), .ZN(n2935) );
  OAI22_X1 U181 ( .A1(n5204), .A2(n6398), .B1(n209), .B2(n231), .ZN(n2936) );
  OAI22_X1 U182 ( .A1(n5172), .A2(n6396), .B1(n209), .B2(n233), .ZN(n2937) );
  OAI22_X1 U183 ( .A1(n5140), .A2(n6393), .B1(n209), .B2(n235), .ZN(n2938) );
  OAI22_X1 U184 ( .A1(n5108), .A2(n6391), .B1(n209), .B2(n237), .ZN(n2939) );
  OAI22_X1 U185 ( .A1(n5076), .A2(n6390), .B1(n209), .B2(n239), .ZN(n2940) );
  OAI22_X1 U186 ( .A1(n5044), .A2(n6388), .B1(n209), .B2(n241), .ZN(n2941) );
  OAI22_X1 U187 ( .A1(n5012), .A2(n6385), .B1(n209), .B2(n243), .ZN(n2942) );
  OAI22_X1 U188 ( .A1(n4980), .A2(n6383), .B1(n209), .B2(n245), .ZN(n2943) );
  OAI22_X1 U189 ( .A1(n4948), .A2(n6382), .B1(n209), .B2(n247), .ZN(n2944) );
  OAI22_X1 U190 ( .A1(n4916), .A2(n6380), .B1(n209), .B2(n249), .ZN(n2945) );
  OAI22_X1 U191 ( .A1(n4884), .A2(n6384), .B1(n209), .B2(n251), .ZN(n2946) );
  OAI22_X1 U192 ( .A1(n4852), .A2(n6381), .B1(n209), .B2(n253), .ZN(n2947) );
  OAI22_X1 U193 ( .A1(n4820), .A2(n6387), .B1(n209), .B2(n255), .ZN(n2948) );
  OAI22_X1 U194 ( .A1(n4788), .A2(n6386), .B1(n209), .B2(n257), .ZN(n2949) );
  OAI22_X1 U195 ( .A1(n4756), .A2(n6392), .B1(n209), .B2(n259), .ZN(n2950) );
  OAI22_X1 U196 ( .A1(n4724), .A2(n6394), .B1(n209), .B2(n261), .ZN(n2951) );
  OAI22_X1 U197 ( .A1(n4692), .A2(n6389), .B1(n209), .B2(n263), .ZN(n2952) );
  OAI22_X1 U198 ( .A1(n4660), .A2(n6395), .B1(n209), .B2(n265), .ZN(n2953) );
  OAI22_X1 U199 ( .A1(n4628), .A2(n6400), .B1(n209), .B2(n267), .ZN(n2954) );
  OAI22_X1 U200 ( .A1(n4596), .A2(n6402), .B1(n209), .B2(n269), .ZN(n2955) );
  OAI22_X1 U201 ( .A1(n4564), .A2(n6397), .B1(n209), .B2(n271), .ZN(n2956) );
  OAI22_X1 U202 ( .A1(n4532), .A2(n6403), .B1(n209), .B2(n273), .ZN(n2957) );
  OAI22_X1 U203 ( .A1(n4500), .A2(n6408), .B1(n209), .B2(n275), .ZN(n2958) );
  OAI22_X1 U204 ( .A1(n4468), .A2(n6405), .B1(n209), .B2(n277), .ZN(n2959) );
  OAI22_X1 U205 ( .A1(n4436), .A2(n6411), .B1(n209), .B2(n279), .ZN(n2960) );
  OAI22_X1 U208 ( .A1(n5479), .A2(net54881), .B1(net54921), .B2(n208), .ZN(
        n2961) );
  AOI221_X1 U209 ( .B1(n283), .B2(n284), .C1(n5605), .C2(n285), .A(n286), .ZN(
        n208) );
  INV_X1 U210 ( .A(n287), .ZN(n286) );
  AOI222_X1 U211 ( .A1(n288), .A2(n289), .B1(n6379), .B2(n5606), .C1(
        \UUT/Mpath/the_mult/x_mult_out[24] ), .C2(n291), .ZN(n287) );
  INV_X1 U212 ( .A(n5644), .ZN(n289) );
  INV_X1 U213 ( .A(n5693), .ZN(n283) );
  OAI221_X1 U214 ( .B1(n292), .B2(n69), .C1(n103), .C2(n71), .A(n293), .ZN(
        n2962) );
  NAND2_X1 U215 ( .A1(\UUT/Mpath/the_mult/x_operand2 [22]), .A2(n6409), .ZN(
        n293) );
  OAI222_X1 U218 ( .A1(n103), .A2(n123), .B1(n292), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N40 ), .C2(net54893), .ZN(n2964) );
  INV_X1 U219 ( .A(n301), .ZN(n103) );
  OAI222_X1 U220 ( .A1(n302), .A2(n129), .B1(n303), .B2(n131), .C1(n5484), 
        .C2(n132), .ZN(n301) );
  OAI221_X1 U221 ( .B1(n133), .B2(n304), .C1(n5695), .C2(n135), .A(n305), .ZN(
        n2965) );
  AOI22_X1 U222 ( .A1(n137), .A2(n306), .B1(\UUT/Mpath/the_mult/Mad_out [54]), 
        .B2(n139), .ZN(n305) );
  OAI221_X1 U223 ( .B1(n140), .B2(n307), .C1(n5648), .C2(n142), .A(n308), .ZN(
        n2966) );
  AOI22_X1 U224 ( .A1(n144), .A2(n306), .B1(\UUT/Mpath/the_mult/Mad_out [22]), 
        .B2(n145), .ZN(n308) );
  INV_X1 U225 ( .A(n5649), .ZN(n306) );
  OAI22_X1 U226 ( .A1(net54905), .A2(n309), .B1(n5649), .B2(net54873), .ZN(
        n2967) );
  OAI221_X1 U227 ( .B1(n302), .B2(n310), .C1(n147), .C2(n309), .A(n311), .ZN(
        n2968) );
  AOI22_X1 U228 ( .A1(n312), .A2(n313), .B1(n314), .B2(n315), .ZN(n311) );
  INV_X1 U229 ( .A(\UUT/Mpath/the_mult/x_operand1[22] ), .ZN(n309) );
  OAI221_X1 U230 ( .B1(n302), .B2(n316), .C1(\UUT/Mpath/the_alu/N39 ), .C2(
        net54885), .A(n317), .ZN(n2969) );
  AOI22_X1 U231 ( .A1(n318), .A2(n313), .B1(n319), .B2(n315), .ZN(n317) );
  OAI22_X1 U232 ( .A1(n5398), .A2(n6407), .B1(n303), .B2(n219), .ZN(n2970) );
  OAI22_X1 U233 ( .A1(n5366), .A2(n6410), .B1(n303), .B2(n221), .ZN(n2971) );
  OAI22_X1 U234 ( .A1(n5334), .A2(n6401), .B1(n303), .B2(n223), .ZN(n2972) );
  OAI22_X1 U235 ( .A1(n5302), .A2(n6406), .B1(n303), .B2(n225), .ZN(n2973) );
  OAI22_X1 U236 ( .A1(n5270), .A2(n6399), .B1(n303), .B2(n227), .ZN(n2974) );
  OAI22_X1 U237 ( .A1(n5238), .A2(n6404), .B1(n303), .B2(n229), .ZN(n2975) );
  OAI22_X1 U238 ( .A1(n5206), .A2(n6398), .B1(n303), .B2(n231), .ZN(n2976) );
  OAI22_X1 U239 ( .A1(n5174), .A2(n6396), .B1(n303), .B2(n233), .ZN(n2977) );
  OAI22_X1 U240 ( .A1(n5142), .A2(n6393), .B1(n303), .B2(n235), .ZN(n2978) );
  OAI22_X1 U241 ( .A1(n5110), .A2(n6391), .B1(n303), .B2(n237), .ZN(n2979) );
  OAI22_X1 U242 ( .A1(n5078), .A2(n6390), .B1(n303), .B2(n239), .ZN(n2980) );
  OAI22_X1 U243 ( .A1(n5046), .A2(n6388), .B1(n303), .B2(n241), .ZN(n2981) );
  OAI22_X1 U244 ( .A1(n5014), .A2(n6385), .B1(n303), .B2(n243), .ZN(n2982) );
  OAI22_X1 U245 ( .A1(n4982), .A2(n6383), .B1(n303), .B2(n245), .ZN(n2983) );
  OAI22_X1 U246 ( .A1(n4950), .A2(n6382), .B1(n303), .B2(n247), .ZN(n2984) );
  OAI22_X1 U247 ( .A1(n4918), .A2(n6380), .B1(n303), .B2(n249), .ZN(n2985) );
  OAI22_X1 U248 ( .A1(n4886), .A2(n6384), .B1(n303), .B2(n251), .ZN(n2986) );
  OAI22_X1 U249 ( .A1(n4854), .A2(n6381), .B1(n303), .B2(n253), .ZN(n2987) );
  OAI22_X1 U250 ( .A1(n4822), .A2(n6387), .B1(n303), .B2(n255), .ZN(n2988) );
  OAI22_X1 U251 ( .A1(n4790), .A2(n6386), .B1(n303), .B2(n257), .ZN(n2989) );
  OAI22_X1 U252 ( .A1(n4758), .A2(n6392), .B1(n303), .B2(n259), .ZN(n2990) );
  OAI22_X1 U253 ( .A1(n4726), .A2(n6394), .B1(n303), .B2(n261), .ZN(n2991) );
  OAI22_X1 U254 ( .A1(n4694), .A2(n6389), .B1(n303), .B2(n263), .ZN(n2992) );
  OAI22_X1 U255 ( .A1(n4662), .A2(n6395), .B1(n303), .B2(n265), .ZN(n2993) );
  OAI22_X1 U256 ( .A1(n4630), .A2(n6400), .B1(n303), .B2(n267), .ZN(n2994) );
  OAI22_X1 U257 ( .A1(n4598), .A2(n6402), .B1(n303), .B2(n269), .ZN(n2995) );
  OAI22_X1 U258 ( .A1(n4566), .A2(n6397), .B1(n303), .B2(n271), .ZN(n2996) );
  OAI22_X1 U259 ( .A1(n4534), .A2(n6403), .B1(n303), .B2(n273), .ZN(n2997) );
  OAI22_X1 U260 ( .A1(n4502), .A2(n6408), .B1(n303), .B2(n275), .ZN(n2998) );
  OAI22_X1 U261 ( .A1(n4470), .A2(n6405), .B1(n303), .B2(n277), .ZN(n2999) );
  OAI22_X1 U262 ( .A1(n4438), .A2(n6411), .B1(n303), .B2(n279), .ZN(n3000) );
  OAI221_X1 U264 ( .B1(n5772), .B2(n281), .C1(n5710), .C2(n5485), .A(n282), 
        .ZN(n315) );
  OAI22_X1 U265 ( .A1(n5485), .A2(net54881), .B1(net54921), .B2(n302), .ZN(
        n3001) );
  INV_X1 U266 ( .A(n320), .ZN(n302) );
  OAI211_X1 U267 ( .C1(n5648), .C2(n321), .A(n322), .B(n323), .ZN(n320) );
  AOI222_X1 U268 ( .A1(n285), .A2(n324), .B1(\UUT/Mpath/out_jar[22] ), .B2(
        n325), .C1(n284), .C2(n326), .ZN(n323) );
  INV_X1 U269 ( .A(n5695), .ZN(n326) );
  AOI22_X1 U270 ( .A1(n6379), .A2(n6100), .B1(
        \UUT/Mpath/the_mult/x_mult_out[22] ), .B2(n291), .ZN(n322) );
  OAI221_X1 U271 ( .B1(n327), .B2(n69), .C1(n102), .C2(n71), .A(n328), .ZN(
        n3002) );
  NAND2_X1 U272 ( .A1(\UUT/Mpath/the_mult/x_operand2 [21]), .A2(n6409), .ZN(
        n328) );
  OAI222_X1 U275 ( .A1(n102), .A2(n123), .B1(n327), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N42 ), .C2(net54893), .ZN(n3004) );
  INV_X1 U276 ( .A(n330), .ZN(n102) );
  OAI222_X1 U277 ( .A1(n331), .A2(n129), .B1(n332), .B2(n131), .C1(n5487), 
        .C2(n132), .ZN(n330) );
  OAI221_X1 U278 ( .B1(n133), .B2(n333), .C1(n5696), .C2(n135), .A(n334), .ZN(
        n3005) );
  AOI22_X1 U279 ( .A1(n137), .A2(n335), .B1(\UUT/Mpath/the_mult/Mad_out [53]), 
        .B2(n139), .ZN(n334) );
  OAI221_X1 U280 ( .B1(n140), .B2(n336), .C1(n5650), .C2(n142), .A(n337), .ZN(
        n3006) );
  AOI22_X1 U281 ( .A1(n144), .A2(n335), .B1(\UUT/Mpath/the_mult/Mad_out [21]), 
        .B2(n145), .ZN(n337) );
  INV_X1 U282 ( .A(n5651), .ZN(n335) );
  OAI22_X1 U283 ( .A1(net54905), .A2(n338), .B1(n5651), .B2(net54875), .ZN(
        n3007) );
  OAI221_X1 U284 ( .B1(n331), .B2(n310), .C1(n147), .C2(n338), .A(n339), .ZN(
        n3008) );
  AOI22_X1 U285 ( .A1(n312), .A2(n340), .B1(n314), .B2(n341), .ZN(n339) );
  INV_X1 U286 ( .A(\UUT/Mpath/the_mult/x_operand1[21] ), .ZN(n338) );
  OAI221_X1 U287 ( .B1(n331), .B2(n316), .C1(\UUT/Mpath/the_alu/N41 ), .C2(
        net54885), .A(n342), .ZN(n3009) );
  AOI22_X1 U288 ( .A1(n318), .A2(n340), .B1(n319), .B2(n341), .ZN(n342) );
  OAI22_X1 U289 ( .A1(n5399), .A2(n218), .B1(n332), .B2(n219), .ZN(n3010) );
  OAI22_X1 U290 ( .A1(n5367), .A2(n220), .B1(n332), .B2(n221), .ZN(n3011) );
  OAI22_X1 U291 ( .A1(n5335), .A2(n222), .B1(n332), .B2(n223), .ZN(n3012) );
  OAI22_X1 U292 ( .A1(n5303), .A2(n224), .B1(n332), .B2(n225), .ZN(n3013) );
  OAI22_X1 U293 ( .A1(n5271), .A2(n226), .B1(n332), .B2(n227), .ZN(n3014) );
  OAI22_X1 U294 ( .A1(n5239), .A2(n228), .B1(n332), .B2(n229), .ZN(n3015) );
  OAI22_X1 U295 ( .A1(n5207), .A2(n230), .B1(n332), .B2(n231), .ZN(n3016) );
  OAI22_X1 U296 ( .A1(n5175), .A2(n232), .B1(n332), .B2(n233), .ZN(n3017) );
  OAI22_X1 U297 ( .A1(n5143), .A2(n234), .B1(n332), .B2(n235), .ZN(n3018) );
  OAI22_X1 U298 ( .A1(n5111), .A2(n236), .B1(n332), .B2(n237), .ZN(n3019) );
  OAI22_X1 U299 ( .A1(n5079), .A2(n238), .B1(n332), .B2(n239), .ZN(n3020) );
  OAI22_X1 U300 ( .A1(n5047), .A2(n240), .B1(n332), .B2(n241), .ZN(n3021) );
  OAI22_X1 U301 ( .A1(n5015), .A2(n242), .B1(n332), .B2(n243), .ZN(n3022) );
  OAI22_X1 U302 ( .A1(n4983), .A2(n244), .B1(n332), .B2(n245), .ZN(n3023) );
  OAI22_X1 U303 ( .A1(n4951), .A2(n246), .B1(n332), .B2(n247), .ZN(n3024) );
  OAI22_X1 U304 ( .A1(n4919), .A2(n248), .B1(n332), .B2(n249), .ZN(n3025) );
  OAI22_X1 U305 ( .A1(n4887), .A2(n250), .B1(n332), .B2(n251), .ZN(n3026) );
  OAI22_X1 U306 ( .A1(n4855), .A2(n252), .B1(n332), .B2(n253), .ZN(n3027) );
  OAI22_X1 U307 ( .A1(n4823), .A2(n254), .B1(n332), .B2(n255), .ZN(n3028) );
  OAI22_X1 U308 ( .A1(n4791), .A2(n256), .B1(n332), .B2(n257), .ZN(n3029) );
  OAI22_X1 U309 ( .A1(n4759), .A2(n258), .B1(n332), .B2(n259), .ZN(n3030) );
  OAI22_X1 U310 ( .A1(n4727), .A2(n260), .B1(n332), .B2(n261), .ZN(n3031) );
  OAI22_X1 U311 ( .A1(n4695), .A2(n262), .B1(n332), .B2(n263), .ZN(n3032) );
  OAI22_X1 U312 ( .A1(n4663), .A2(n264), .B1(n332), .B2(n265), .ZN(n3033) );
  OAI22_X1 U313 ( .A1(n4631), .A2(n266), .B1(n332), .B2(n267), .ZN(n3034) );
  OAI22_X1 U314 ( .A1(n4599), .A2(n268), .B1(n332), .B2(n269), .ZN(n3035) );
  OAI22_X1 U315 ( .A1(n4567), .A2(n270), .B1(n332), .B2(n271), .ZN(n3036) );
  OAI22_X1 U316 ( .A1(n4535), .A2(n272), .B1(n332), .B2(n273), .ZN(n3037) );
  OAI22_X1 U317 ( .A1(n4503), .A2(n274), .B1(n332), .B2(n275), .ZN(n3038) );
  OAI22_X1 U318 ( .A1(n4471), .A2(n276), .B1(n332), .B2(n277), .ZN(n3039) );
  OAI22_X1 U319 ( .A1(n4439), .A2(n278), .B1(n332), .B2(n279), .ZN(n3040) );
  OAI221_X1 U321 ( .B1(n5789), .B2(n281), .C1(n5710), .C2(n5488), .A(n282), 
        .ZN(n341) );
  OAI22_X1 U322 ( .A1(n5488), .A2(net54881), .B1(net54921), .B2(n331), .ZN(
        n3041) );
  INV_X1 U323 ( .A(n343), .ZN(n331) );
  OAI211_X1 U324 ( .C1(n5650), .C2(n321), .A(n344), .B(n345), .ZN(n343) );
  AOI222_X1 U325 ( .A1(n285), .A2(n346), .B1(\UUT/Mpath/out_jar[21] ), .B2(
        n325), .C1(n284), .C2(n347), .ZN(n345) );
  INV_X1 U326 ( .A(n5696), .ZN(n347) );
  AOI22_X1 U327 ( .A1(n6379), .A2(n6107), .B1(
        \UUT/Mpath/the_mult/x_mult_out[21] ), .B2(n291), .ZN(n344) );
  OAI221_X1 U328 ( .B1(n348), .B2(n69), .C1(n101), .C2(n71), .A(n349), .ZN(
        n3042) );
  NAND2_X1 U329 ( .A1(\UUT/Mpath/the_mult/x_operand2 [20]), .A2(n6409), .ZN(
        n349) );
  OAI222_X1 U332 ( .A1(n101), .A2(n123), .B1(n348), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N44 ), .C2(net54893), .ZN(n3044) );
  INV_X1 U333 ( .A(n351), .ZN(n101) );
  OAI222_X1 U334 ( .A1(n352), .A2(n129), .B1(n353), .B2(n131), .C1(n5490), 
        .C2(n132), .ZN(n351) );
  OAI221_X1 U335 ( .B1(n133), .B2(n354), .C1(n5697), .C2(n135), .A(n355), .ZN(
        n3045) );
  AOI22_X1 U336 ( .A1(n137), .A2(n356), .B1(\UUT/Mpath/the_mult/Mad_out [52]), 
        .B2(n139), .ZN(n355) );
  OAI221_X1 U337 ( .B1(n140), .B2(n357), .C1(n5652), .C2(n142), .A(n358), .ZN(
        n3046) );
  AOI22_X1 U338 ( .A1(n144), .A2(n356), .B1(\UUT/Mpath/the_mult/Mad_out [20]), 
        .B2(n145), .ZN(n358) );
  INV_X1 U339 ( .A(n5653), .ZN(n356) );
  OAI22_X1 U340 ( .A1(net54905), .A2(n359), .B1(n5653), .B2(net54873), .ZN(
        n3047) );
  OAI221_X1 U341 ( .B1(n352), .B2(n310), .C1(n147), .C2(n359), .A(n360), .ZN(
        n3048) );
  AOI22_X1 U342 ( .A1(n312), .A2(n361), .B1(n314), .B2(n362), .ZN(n360) );
  INV_X1 U343 ( .A(\UUT/Mpath/the_mult/x_operand1[20] ), .ZN(n359) );
  OAI221_X1 U344 ( .B1(n352), .B2(n316), .C1(\UUT/Mpath/the_alu/N43 ), .C2(
        net54887), .A(n363), .ZN(n3049) );
  AOI22_X1 U345 ( .A1(n318), .A2(n361), .B1(n319), .B2(n362), .ZN(n363) );
  OAI22_X1 U346 ( .A1(n5400), .A2(n6407), .B1(n353), .B2(n219), .ZN(n3050) );
  OAI22_X1 U347 ( .A1(n5368), .A2(n6410), .B1(n353), .B2(n221), .ZN(n3051) );
  OAI22_X1 U348 ( .A1(n5336), .A2(n6401), .B1(n353), .B2(n223), .ZN(n3052) );
  OAI22_X1 U349 ( .A1(n5304), .A2(n6406), .B1(n353), .B2(n225), .ZN(n3053) );
  OAI22_X1 U350 ( .A1(n5272), .A2(n6399), .B1(n353), .B2(n227), .ZN(n3054) );
  OAI22_X1 U351 ( .A1(n5240), .A2(n6404), .B1(n353), .B2(n229), .ZN(n3055) );
  OAI22_X1 U352 ( .A1(n5208), .A2(n6398), .B1(n353), .B2(n231), .ZN(n3056) );
  OAI22_X1 U353 ( .A1(n5176), .A2(n6396), .B1(n353), .B2(n233), .ZN(n3057) );
  OAI22_X1 U354 ( .A1(n5144), .A2(n6393), .B1(n353), .B2(n235), .ZN(n3058) );
  OAI22_X1 U355 ( .A1(n5112), .A2(n6391), .B1(n353), .B2(n237), .ZN(n3059) );
  OAI22_X1 U356 ( .A1(n5080), .A2(n6390), .B1(n353), .B2(n239), .ZN(n3060) );
  OAI22_X1 U357 ( .A1(n5048), .A2(n6388), .B1(n353), .B2(n241), .ZN(n3061) );
  OAI22_X1 U358 ( .A1(n5016), .A2(n6385), .B1(n353), .B2(n243), .ZN(n3062) );
  OAI22_X1 U359 ( .A1(n4984), .A2(n6383), .B1(n353), .B2(n245), .ZN(n3063) );
  OAI22_X1 U360 ( .A1(n4952), .A2(n6382), .B1(n353), .B2(n247), .ZN(n3064) );
  OAI22_X1 U361 ( .A1(n4920), .A2(n6380), .B1(n353), .B2(n249), .ZN(n3065) );
  OAI22_X1 U362 ( .A1(n4888), .A2(n6384), .B1(n353), .B2(n251), .ZN(n3066) );
  OAI22_X1 U363 ( .A1(n4856), .A2(n6381), .B1(n353), .B2(n253), .ZN(n3067) );
  OAI22_X1 U364 ( .A1(n4824), .A2(n6387), .B1(n353), .B2(n255), .ZN(n3068) );
  OAI22_X1 U365 ( .A1(n4792), .A2(n6386), .B1(n353), .B2(n257), .ZN(n3069) );
  OAI22_X1 U366 ( .A1(n4760), .A2(n6392), .B1(n353), .B2(n259), .ZN(n3070) );
  OAI22_X1 U367 ( .A1(n4728), .A2(n6394), .B1(n353), .B2(n261), .ZN(n3071) );
  OAI22_X1 U368 ( .A1(n4696), .A2(n6389), .B1(n353), .B2(n263), .ZN(n3072) );
  OAI22_X1 U369 ( .A1(n4664), .A2(n6395), .B1(n353), .B2(n265), .ZN(n3073) );
  OAI22_X1 U370 ( .A1(n4632), .A2(n6400), .B1(n353), .B2(n267), .ZN(n3074) );
  OAI22_X1 U371 ( .A1(n4600), .A2(n6402), .B1(n353), .B2(n269), .ZN(n3075) );
  OAI22_X1 U372 ( .A1(n4568), .A2(n6397), .B1(n353), .B2(n271), .ZN(n3076) );
  OAI22_X1 U373 ( .A1(n4536), .A2(n6403), .B1(n353), .B2(n273), .ZN(n3077) );
  OAI22_X1 U374 ( .A1(n4504), .A2(n6408), .B1(n353), .B2(n275), .ZN(n3078) );
  OAI22_X1 U375 ( .A1(n4472), .A2(n6405), .B1(n353), .B2(n277), .ZN(n3079) );
  OAI22_X1 U376 ( .A1(n4440), .A2(n6411), .B1(n353), .B2(n279), .ZN(n3080) );
  OAI221_X1 U378 ( .B1(n5802), .B2(n281), .C1(n5710), .C2(n5491), .A(n282), 
        .ZN(n362) );
  OAI22_X1 U379 ( .A1(n5491), .A2(net54883), .B1(net54921), .B2(n352), .ZN(
        n3081) );
  INV_X1 U380 ( .A(n364), .ZN(n352) );
  OAI211_X1 U381 ( .C1(n5652), .C2(n321), .A(n365), .B(n366), .ZN(n364) );
  AOI222_X1 U382 ( .A1(n285), .A2(n367), .B1(\UUT/Mpath/out_jar[20] ), .B2(
        n325), .C1(n284), .C2(n368), .ZN(n366) );
  INV_X1 U383 ( .A(n5697), .ZN(n368) );
  AOI22_X1 U384 ( .A1(n6379), .A2(n6114), .B1(
        \UUT/Mpath/the_mult/x_mult_out[20] ), .B2(n291), .ZN(n365) );
  OAI221_X1 U385 ( .B1(n369), .B2(n69), .C1(n100), .C2(n71), .A(n370), .ZN(
        n3082) );
  NAND2_X1 U386 ( .A1(\UUT/Mpath/the_mult/x_operand2 [19]), .A2(n6409), .ZN(
        n370) );
  INV_X1 U387 ( .A(n371), .ZN(n100) );
  INV_X1 U390 ( .A(\UUT/break_code[19] ), .ZN(n369) );
  OAI211_X1 U391 ( .C1(\UUT/Mpath/the_alu/N46 ), .C2(net54895), .A(n373), .B(
        n374), .ZN(n3084) );
  AOI222_X1 U392 ( .A1(n375), .A2(n371), .B1(n376), .B2(
        \UUT/Mcontrol/d_sampled_finstr [3]), .C1(n377), .C2(n6126), .ZN(n374)
         );
  OAI222_X1 U393 ( .A1(n378), .A2(n129), .B1(n379), .B2(n131), .C1(n5496), 
        .C2(n132), .ZN(n371) );
  OAI221_X1 U394 ( .B1(n133), .B2(n380), .C1(n5699), .C2(n135), .A(n381), .ZN(
        n3085) );
  AOI22_X1 U395 ( .A1(n137), .A2(n382), .B1(\UUT/Mpath/the_mult/Mad_out [51]), 
        .B2(n139), .ZN(n381) );
  OAI221_X1 U396 ( .B1(n140), .B2(n383), .C1(n5656), .C2(n142), .A(n384), .ZN(
        n3086) );
  AOI22_X1 U397 ( .A1(n144), .A2(n382), .B1(\UUT/Mpath/the_mult/Mad_out [19]), 
        .B2(n145), .ZN(n384) );
  INV_X1 U398 ( .A(n5657), .ZN(n382) );
  OAI22_X1 U399 ( .A1(net54905), .A2(n385), .B1(n5657), .B2(net54873), .ZN(
        n3087) );
  OAI221_X1 U400 ( .B1(n378), .B2(n310), .C1(n147), .C2(n385), .A(n386), .ZN(
        n3088) );
  AOI22_X1 U401 ( .A1(n312), .A2(n387), .B1(n314), .B2(n388), .ZN(n386) );
  INV_X1 U402 ( .A(\UUT/Mpath/the_mult/x_operand1[19] ), .ZN(n385) );
  OAI221_X1 U403 ( .B1(n378), .B2(n316), .C1(\UUT/Mpath/the_alu/N45 ), .C2(
        net54885), .A(n389), .ZN(n3089) );
  AOI22_X1 U404 ( .A1(n318), .A2(n387), .B1(n319), .B2(n388), .ZN(n389) );
  OAI22_X1 U405 ( .A1(n5402), .A2(n218), .B1(n379), .B2(n219), .ZN(n3090) );
  OAI22_X1 U406 ( .A1(n5370), .A2(n220), .B1(n379), .B2(n221), .ZN(n3091) );
  OAI22_X1 U407 ( .A1(n5338), .A2(n222), .B1(n379), .B2(n223), .ZN(n3092) );
  OAI22_X1 U408 ( .A1(n5306), .A2(n224), .B1(n379), .B2(n225), .ZN(n3093) );
  OAI22_X1 U409 ( .A1(n5274), .A2(n226), .B1(n379), .B2(n227), .ZN(n3094) );
  OAI22_X1 U410 ( .A1(n5242), .A2(n228), .B1(n379), .B2(n229), .ZN(n3095) );
  OAI22_X1 U411 ( .A1(n5210), .A2(n230), .B1(n379), .B2(n231), .ZN(n3096) );
  OAI22_X1 U412 ( .A1(n5178), .A2(n232), .B1(n379), .B2(n233), .ZN(n3097) );
  OAI22_X1 U413 ( .A1(n5146), .A2(n234), .B1(n379), .B2(n235), .ZN(n3098) );
  OAI22_X1 U414 ( .A1(n5114), .A2(n236), .B1(n379), .B2(n237), .ZN(n3099) );
  OAI22_X1 U415 ( .A1(n5082), .A2(n238), .B1(n379), .B2(n239), .ZN(n3100) );
  OAI22_X1 U416 ( .A1(n5050), .A2(n240), .B1(n379), .B2(n241), .ZN(n3101) );
  OAI22_X1 U417 ( .A1(n5018), .A2(n242), .B1(n379), .B2(n243), .ZN(n3102) );
  OAI22_X1 U418 ( .A1(n4986), .A2(n244), .B1(n379), .B2(n245), .ZN(n3103) );
  OAI22_X1 U419 ( .A1(n4954), .A2(n246), .B1(n379), .B2(n247), .ZN(n3104) );
  OAI22_X1 U420 ( .A1(n4922), .A2(n248), .B1(n379), .B2(n249), .ZN(n3105) );
  OAI22_X1 U421 ( .A1(n4890), .A2(n250), .B1(n379), .B2(n251), .ZN(n3106) );
  OAI22_X1 U422 ( .A1(n4858), .A2(n252), .B1(n379), .B2(n253), .ZN(n3107) );
  OAI22_X1 U423 ( .A1(n4826), .A2(n254), .B1(n379), .B2(n255), .ZN(n3108) );
  OAI22_X1 U424 ( .A1(n4794), .A2(n256), .B1(n379), .B2(n257), .ZN(n3109) );
  OAI22_X1 U425 ( .A1(n4762), .A2(n258), .B1(n379), .B2(n259), .ZN(n3110) );
  OAI22_X1 U426 ( .A1(n4730), .A2(n260), .B1(n379), .B2(n261), .ZN(n3111) );
  OAI22_X1 U427 ( .A1(n4698), .A2(n262), .B1(n379), .B2(n263), .ZN(n3112) );
  OAI22_X1 U428 ( .A1(n4666), .A2(n264), .B1(n379), .B2(n265), .ZN(n3113) );
  OAI22_X1 U429 ( .A1(n4634), .A2(n266), .B1(n379), .B2(n267), .ZN(n3114) );
  OAI22_X1 U430 ( .A1(n4602), .A2(n268), .B1(n379), .B2(n269), .ZN(n3115) );
  OAI22_X1 U431 ( .A1(n4570), .A2(n270), .B1(n379), .B2(n271), .ZN(n3116) );
  OAI22_X1 U432 ( .A1(n4538), .A2(n272), .B1(n379), .B2(n273), .ZN(n3117) );
  OAI22_X1 U433 ( .A1(n4506), .A2(n274), .B1(n379), .B2(n275), .ZN(n3118) );
  OAI22_X1 U434 ( .A1(n4474), .A2(n276), .B1(n379), .B2(n277), .ZN(n3119) );
  OAI22_X1 U435 ( .A1(n4442), .A2(n278), .B1(n379), .B2(n279), .ZN(n3120) );
  OAI221_X1 U437 ( .B1(n5815), .B2(n281), .C1(n5710), .C2(n5497), .A(n282), 
        .ZN(n388) );
  OAI22_X1 U438 ( .A1(n5497), .A2(net54883), .B1(net54921), .B2(n378), .ZN(
        n3121) );
  INV_X1 U439 ( .A(n390), .ZN(n378) );
  OAI211_X1 U440 ( .C1(n5656), .C2(n321), .A(n391), .B(n392), .ZN(n390) );
  AOI222_X1 U441 ( .A1(n285), .A2(n393), .B1(\UUT/Mpath/out_jar[19] ), .B2(
        n325), .C1(n284), .C2(n394), .ZN(n392) );
  INV_X1 U442 ( .A(n5699), .ZN(n394) );
  AOI22_X1 U443 ( .A1(n6379), .A2(n6124), .B1(
        \UUT/Mpath/the_mult/x_mult_out[19] ), .B2(n291), .ZN(n391) );
  OAI221_X1 U444 ( .B1(n395), .B2(n69), .C1(n99), .C2(n71), .A(n396), .ZN(
        n3122) );
  NAND2_X1 U445 ( .A1(\UUT/Mpath/the_mult/x_operand2 [18]), .A2(n6409), .ZN(
        n396) );
  INV_X1 U446 ( .A(n397), .ZN(n99) );
  INV_X1 U449 ( .A(\UUT/break_code[18] ), .ZN(n395) );
  OAI211_X1 U450 ( .C1(\UUT/Mpath/the_alu/N48 ), .C2(net54895), .A(n373), .B(
        n399), .ZN(n3124) );
  AOI222_X1 U451 ( .A1(n375), .A2(n397), .B1(n376), .B2(
        \UUT/Mcontrol/d_sampled_finstr [2]), .C1(n6135), .C2(n377), .ZN(n399)
         );
  OAI222_X1 U452 ( .A1(n400), .A2(n129), .B1(n401), .B2(n131), .C1(n5499), 
        .C2(n132), .ZN(n397) );
  OAI221_X1 U453 ( .B1(n133), .B2(n402), .C1(n5700), .C2(n135), .A(n403), .ZN(
        n3125) );
  AOI22_X1 U454 ( .A1(n137), .A2(n404), .B1(\UUT/Mpath/the_mult/Mad_out [50]), 
        .B2(n139), .ZN(n403) );
  OAI221_X1 U455 ( .B1(n140), .B2(n405), .C1(n5658), .C2(n142), .A(n406), .ZN(
        n3126) );
  AOI22_X1 U456 ( .A1(n144), .A2(n404), .B1(\UUT/Mpath/the_mult/Mad_out [18]), 
        .B2(n145), .ZN(n406) );
  INV_X1 U457 ( .A(n5659), .ZN(n404) );
  OAI22_X1 U458 ( .A1(net54907), .A2(n407), .B1(n5659), .B2(net54873), .ZN(
        n3127) );
  OAI221_X1 U459 ( .B1(n400), .B2(n310), .C1(n147), .C2(n407), .A(n408), .ZN(
        n3128) );
  AOI22_X1 U460 ( .A1(n312), .A2(n409), .B1(n314), .B2(n410), .ZN(n408) );
  INV_X1 U461 ( .A(\UUT/Mpath/the_mult/x_operand1[18] ), .ZN(n407) );
  OAI221_X1 U462 ( .B1(n400), .B2(n316), .C1(\UUT/Mpath/the_alu/N47 ), .C2(
        net54885), .A(n411), .ZN(n3129) );
  AOI22_X1 U463 ( .A1(n318), .A2(n409), .B1(n319), .B2(n410), .ZN(n411) );
  OAI22_X1 U464 ( .A1(n5403), .A2(n6407), .B1(n401), .B2(n219), .ZN(n3130) );
  OAI22_X1 U465 ( .A1(n5371), .A2(n6410), .B1(n401), .B2(n221), .ZN(n3131) );
  OAI22_X1 U466 ( .A1(n5339), .A2(n6401), .B1(n401), .B2(n223), .ZN(n3132) );
  OAI22_X1 U467 ( .A1(n5307), .A2(n6406), .B1(n401), .B2(n225), .ZN(n3133) );
  OAI22_X1 U468 ( .A1(n5275), .A2(n6399), .B1(n401), .B2(n227), .ZN(n3134) );
  OAI22_X1 U469 ( .A1(n5243), .A2(n6404), .B1(n401), .B2(n229), .ZN(n3135) );
  OAI22_X1 U470 ( .A1(n5211), .A2(n6398), .B1(n401), .B2(n231), .ZN(n3136) );
  OAI22_X1 U471 ( .A1(n5179), .A2(n6396), .B1(n401), .B2(n233), .ZN(n3137) );
  OAI22_X1 U472 ( .A1(n5147), .A2(n6393), .B1(n401), .B2(n235), .ZN(n3138) );
  OAI22_X1 U473 ( .A1(n5115), .A2(n6391), .B1(n401), .B2(n237), .ZN(n3139) );
  OAI22_X1 U474 ( .A1(n5083), .A2(n6390), .B1(n401), .B2(n239), .ZN(n3140) );
  OAI22_X1 U475 ( .A1(n5051), .A2(n6388), .B1(n401), .B2(n241), .ZN(n3141) );
  OAI22_X1 U476 ( .A1(n5019), .A2(n6385), .B1(n401), .B2(n243), .ZN(n3142) );
  OAI22_X1 U477 ( .A1(n4987), .A2(n6383), .B1(n401), .B2(n245), .ZN(n3143) );
  OAI22_X1 U478 ( .A1(n4955), .A2(n6382), .B1(n401), .B2(n247), .ZN(n3144) );
  OAI22_X1 U479 ( .A1(n4923), .A2(n6380), .B1(n401), .B2(n249), .ZN(n3145) );
  OAI22_X1 U480 ( .A1(n4891), .A2(n6384), .B1(n401), .B2(n251), .ZN(n3146) );
  OAI22_X1 U481 ( .A1(n4859), .A2(n6381), .B1(n401), .B2(n253), .ZN(n3147) );
  OAI22_X1 U482 ( .A1(n4827), .A2(n6387), .B1(n401), .B2(n255), .ZN(n3148) );
  OAI22_X1 U483 ( .A1(n4795), .A2(n6386), .B1(n401), .B2(n257), .ZN(n3149) );
  OAI22_X1 U484 ( .A1(n4763), .A2(n6392), .B1(n401), .B2(n259), .ZN(n3150) );
  OAI22_X1 U485 ( .A1(n4731), .A2(n6394), .B1(n401), .B2(n261), .ZN(n3151) );
  OAI22_X1 U486 ( .A1(n4699), .A2(n6389), .B1(n401), .B2(n263), .ZN(n3152) );
  OAI22_X1 U487 ( .A1(n4667), .A2(n6395), .B1(n401), .B2(n265), .ZN(n3153) );
  OAI22_X1 U488 ( .A1(n4635), .A2(n6400), .B1(n401), .B2(n267), .ZN(n3154) );
  OAI22_X1 U489 ( .A1(n4603), .A2(n6402), .B1(n401), .B2(n269), .ZN(n3155) );
  OAI22_X1 U490 ( .A1(n4571), .A2(n6397), .B1(n401), .B2(n271), .ZN(n3156) );
  OAI22_X1 U491 ( .A1(n4539), .A2(n6403), .B1(n401), .B2(n273), .ZN(n3157) );
  OAI22_X1 U492 ( .A1(n4507), .A2(n6408), .B1(n401), .B2(n275), .ZN(n3158) );
  OAI22_X1 U493 ( .A1(n4475), .A2(n6405), .B1(n401), .B2(n277), .ZN(n3159) );
  OAI22_X1 U494 ( .A1(n4443), .A2(n6411), .B1(n401), .B2(n279), .ZN(n3160) );
  OAI221_X1 U496 ( .B1(n5841), .B2(n281), .C1(n5710), .C2(n5500), .A(n282), 
        .ZN(n410) );
  OAI22_X1 U497 ( .A1(n5500), .A2(net54883), .B1(net54921), .B2(n400), .ZN(
        n3161) );
  INV_X1 U498 ( .A(n412), .ZN(n400) );
  OAI211_X1 U499 ( .C1(n5658), .C2(n321), .A(n413), .B(n414), .ZN(n412) );
  AOI222_X1 U500 ( .A1(n285), .A2(n415), .B1(\UUT/Mpath/out_jar[18] ), .B2(
        n325), .C1(n284), .C2(n416), .ZN(n414) );
  INV_X1 U501 ( .A(n5700), .ZN(n416) );
  AOI22_X1 U502 ( .A1(n6379), .A2(n6134), .B1(
        \UUT/Mpath/the_mult/x_mult_out[18] ), .B2(n291), .ZN(n413) );
  OAI221_X1 U503 ( .B1(n417), .B2(n69), .C1(n98), .C2(n71), .A(n418), .ZN(
        n3162) );
  NAND2_X1 U504 ( .A1(\UUT/Mpath/the_mult/x_operand2 [17]), .A2(n6409), .ZN(
        n418) );
  INV_X1 U505 ( .A(n419), .ZN(n98) );
  INV_X1 U508 ( .A(\UUT/break_code[17] ), .ZN(n417) );
  OAI211_X1 U509 ( .C1(\UUT/Mpath/the_alu/N50 ), .C2(net54895), .A(n373), .B(
        n421), .ZN(n3164) );
  AOI222_X1 U510 ( .A1(n375), .A2(n419), .B1(n376), .B2(
        \UUT/Mcontrol/d_sampled_finstr [1]), .C1(n6153), .C2(n377), .ZN(n421)
         );
  OAI222_X1 U511 ( .A1(n422), .A2(n129), .B1(n423), .B2(n131), .C1(n5502), 
        .C2(n132), .ZN(n419) );
  OAI221_X1 U512 ( .B1(n133), .B2(n424), .C1(n5701), .C2(n135), .A(n425), .ZN(
        n3165) );
  AOI22_X1 U513 ( .A1(n137), .A2(n426), .B1(\UUT/Mpath/the_mult/Mad_out [49]), 
        .B2(n139), .ZN(n425) );
  OAI221_X1 U514 ( .B1(n140), .B2(n427), .C1(n5660), .C2(n142), .A(n428), .ZN(
        n3166) );
  AOI22_X1 U515 ( .A1(n144), .A2(n426), .B1(\UUT/Mpath/the_mult/Mad_out [17]), 
        .B2(n145), .ZN(n428) );
  INV_X1 U516 ( .A(n5661), .ZN(n426) );
  OAI22_X1 U517 ( .A1(net54905), .A2(n429), .B1(n5661), .B2(net54873), .ZN(
        n3167) );
  OAI221_X1 U518 ( .B1(n422), .B2(n310), .C1(n147), .C2(n429), .A(n430), .ZN(
        n3168) );
  AOI22_X1 U519 ( .A1(n312), .A2(n431), .B1(n314), .B2(n432), .ZN(n430) );
  INV_X1 U520 ( .A(\UUT/Mpath/the_mult/x_operand1[17] ), .ZN(n429) );
  OAI221_X1 U521 ( .B1(n422), .B2(n316), .C1(\UUT/Mpath/the_alu/N49 ), .C2(
        net54885), .A(n433), .ZN(n3169) );
  AOI22_X1 U522 ( .A1(n318), .A2(n431), .B1(n319), .B2(n432), .ZN(n433) );
  OAI22_X1 U523 ( .A1(n5404), .A2(n6407), .B1(n423), .B2(n219), .ZN(n3170) );
  OAI22_X1 U524 ( .A1(n5372), .A2(n6410), .B1(n423), .B2(n221), .ZN(n3171) );
  OAI22_X1 U525 ( .A1(n5340), .A2(n6401), .B1(n423), .B2(n223), .ZN(n3172) );
  OAI22_X1 U526 ( .A1(n5308), .A2(n6406), .B1(n423), .B2(n225), .ZN(n3173) );
  OAI22_X1 U527 ( .A1(n5276), .A2(n6399), .B1(n423), .B2(n227), .ZN(n3174) );
  OAI22_X1 U528 ( .A1(n5244), .A2(n6404), .B1(n423), .B2(n229), .ZN(n3175) );
  OAI22_X1 U529 ( .A1(n5212), .A2(n6398), .B1(n423), .B2(n231), .ZN(n3176) );
  OAI22_X1 U530 ( .A1(n5180), .A2(n6396), .B1(n423), .B2(n233), .ZN(n3177) );
  OAI22_X1 U531 ( .A1(n5148), .A2(n6393), .B1(n423), .B2(n235), .ZN(n3178) );
  OAI22_X1 U532 ( .A1(n5116), .A2(n6391), .B1(n423), .B2(n237), .ZN(n3179) );
  OAI22_X1 U533 ( .A1(n5084), .A2(n6390), .B1(n423), .B2(n239), .ZN(n3180) );
  OAI22_X1 U534 ( .A1(n5052), .A2(n6388), .B1(n423), .B2(n241), .ZN(n3181) );
  OAI22_X1 U535 ( .A1(n5020), .A2(n6385), .B1(n423), .B2(n243), .ZN(n3182) );
  OAI22_X1 U536 ( .A1(n4988), .A2(n6383), .B1(n423), .B2(n245), .ZN(n3183) );
  OAI22_X1 U537 ( .A1(n4956), .A2(n6382), .B1(n423), .B2(n247), .ZN(n3184) );
  OAI22_X1 U538 ( .A1(n4924), .A2(n6380), .B1(n423), .B2(n249), .ZN(n3185) );
  OAI22_X1 U539 ( .A1(n4892), .A2(n6384), .B1(n423), .B2(n251), .ZN(n3186) );
  OAI22_X1 U540 ( .A1(n4860), .A2(n6381), .B1(n423), .B2(n253), .ZN(n3187) );
  OAI22_X1 U541 ( .A1(n4828), .A2(n6387), .B1(n423), .B2(n255), .ZN(n3188) );
  OAI22_X1 U542 ( .A1(n4796), .A2(n6386), .B1(n423), .B2(n257), .ZN(n3189) );
  OAI22_X1 U543 ( .A1(n4764), .A2(n6392), .B1(n423), .B2(n259), .ZN(n3190) );
  OAI22_X1 U544 ( .A1(n4732), .A2(n6394), .B1(n423), .B2(n261), .ZN(n3191) );
  OAI22_X1 U545 ( .A1(n4700), .A2(n6389), .B1(n423), .B2(n263), .ZN(n3192) );
  OAI22_X1 U546 ( .A1(n4668), .A2(n6395), .B1(n423), .B2(n265), .ZN(n3193) );
  OAI22_X1 U547 ( .A1(n4636), .A2(n6400), .B1(n423), .B2(n267), .ZN(n3194) );
  OAI22_X1 U548 ( .A1(n4604), .A2(n6402), .B1(n423), .B2(n269), .ZN(n3195) );
  OAI22_X1 U549 ( .A1(n4572), .A2(n6397), .B1(n423), .B2(n271), .ZN(n3196) );
  OAI22_X1 U550 ( .A1(n4540), .A2(n6403), .B1(n423), .B2(n273), .ZN(n3197) );
  OAI22_X1 U551 ( .A1(n4508), .A2(n6408), .B1(n423), .B2(n275), .ZN(n3198) );
  OAI22_X1 U552 ( .A1(n4476), .A2(n6405), .B1(n423), .B2(n277), .ZN(n3199) );
  OAI22_X1 U553 ( .A1(n4444), .A2(n6411), .B1(n423), .B2(n279), .ZN(n3200) );
  OAI221_X1 U555 ( .B1(n5919), .B2(n281), .C1(n5710), .C2(n5503), .A(n282), 
        .ZN(n432) );
  OAI22_X1 U556 ( .A1(n5503), .A2(net54881), .B1(net54923), .B2(n422), .ZN(
        n3201) );
  INV_X1 U557 ( .A(n434), .ZN(n422) );
  OAI211_X1 U558 ( .C1(n5660), .C2(n321), .A(n435), .B(n436), .ZN(n434) );
  AOI222_X1 U559 ( .A1(n285), .A2(n437), .B1(\UUT/Mpath/out_jar[17] ), .B2(
        n325), .C1(n284), .C2(n438), .ZN(n436) );
  INV_X1 U560 ( .A(n5701), .ZN(n438) );
  AOI22_X1 U561 ( .A1(n6379), .A2(n6152), .B1(
        \UUT/Mpath/the_mult/x_mult_out[17] ), .B2(n291), .ZN(n435) );
  OAI221_X1 U562 ( .B1(n439), .B2(n69), .C1(n97), .C2(n71), .A(n440), .ZN(
        n3202) );
  NAND2_X1 U563 ( .A1(\UUT/Mpath/the_mult/x_operand2 [16]), .A2(n6409), .ZN(
        n440) );
  INV_X1 U564 ( .A(n441), .ZN(n97) );
  INV_X1 U567 ( .A(\UUT/break_code[16] ), .ZN(n439) );
  OAI211_X1 U568 ( .C1(\UUT/Mpath/the_alu/N52 ), .C2(net54895), .A(n373), .B(
        n443), .ZN(n3204) );
  AOI222_X1 U569 ( .A1(n375), .A2(n441), .B1(n376), .B2(
        \UUT/Mcontrol/d_sampled_finstr [0]), .C1(n6162), .C2(n377), .ZN(n443)
         );
  AND2_X1 U570 ( .A1(n444), .A2(n445), .ZN(n377) );
  AND2_X1 U571 ( .A1(n125), .A2(net54895), .ZN(n376) );
  OAI222_X1 U572 ( .A1(n446), .A2(n129), .B1(n447), .B2(n131), .C1(n5505), 
        .C2(n132), .ZN(n441) );
  INV_X1 U573 ( .A(n123), .ZN(n375) );
  AOI22_X1 U574 ( .A1(n448), .A2(n449), .B1(n6127), .B2(n444), .ZN(n373) );
  NOR3_X1 U575 ( .A1(net54953), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .A3(n450), .ZN(n444) );
  OAI221_X1 U576 ( .B1(n133), .B2(n451), .C1(n5702), .C2(n135), .A(n452), .ZN(
        n3205) );
  AOI22_X1 U577 ( .A1(n137), .A2(n453), .B1(\UUT/Mpath/the_mult/Mad_out [48]), 
        .B2(n139), .ZN(n452) );
  OAI221_X1 U578 ( .B1(n140), .B2(n454), .C1(n5662), .C2(n142), .A(n455), .ZN(
        n3206) );
  AOI22_X1 U579 ( .A1(n144), .A2(n453), .B1(\UUT/Mpath/the_mult/Mad_out [16]), 
        .B2(n145), .ZN(n455) );
  INV_X1 U580 ( .A(n5663), .ZN(n453) );
  OAI22_X1 U581 ( .A1(net54905), .A2(n456), .B1(n5663), .B2(net54873), .ZN(
        n3207) );
  OAI221_X1 U582 ( .B1(n446), .B2(n310), .C1(n147), .C2(n456), .A(n457), .ZN(
        n3208) );
  AOI22_X1 U583 ( .A1(n312), .A2(n458), .B1(n314), .B2(n459), .ZN(n457) );
  INV_X1 U584 ( .A(\UUT/Mpath/the_mult/x_operand1[16] ), .ZN(n456) );
  OAI221_X1 U585 ( .B1(n446), .B2(n316), .C1(\UUT/Mpath/the_alu/N51 ), .C2(
        net54885), .A(n460), .ZN(n3209) );
  AOI22_X1 U586 ( .A1(n318), .A2(n458), .B1(n319), .B2(n459), .ZN(n460) );
  OAI22_X1 U587 ( .A1(n5405), .A2(n6407), .B1(n447), .B2(n219), .ZN(n3210) );
  OAI22_X1 U588 ( .A1(n5373), .A2(n6410), .B1(n447), .B2(n221), .ZN(n3211) );
  OAI22_X1 U589 ( .A1(n5341), .A2(n6401), .B1(n447), .B2(n223), .ZN(n3212) );
  OAI22_X1 U590 ( .A1(n5309), .A2(n6406), .B1(n447), .B2(n225), .ZN(n3213) );
  OAI22_X1 U591 ( .A1(n5277), .A2(n6399), .B1(n447), .B2(n227), .ZN(n3214) );
  OAI22_X1 U592 ( .A1(n5245), .A2(n6404), .B1(n447), .B2(n229), .ZN(n3215) );
  OAI22_X1 U593 ( .A1(n5213), .A2(n6398), .B1(n447), .B2(n231), .ZN(n3216) );
  OAI22_X1 U594 ( .A1(n5181), .A2(n6396), .B1(n447), .B2(n233), .ZN(n3217) );
  OAI22_X1 U595 ( .A1(n5149), .A2(n6393), .B1(n447), .B2(n235), .ZN(n3218) );
  OAI22_X1 U596 ( .A1(n5117), .A2(n6391), .B1(n447), .B2(n237), .ZN(n3219) );
  OAI22_X1 U597 ( .A1(n5085), .A2(n6390), .B1(n447), .B2(n239), .ZN(n3220) );
  OAI22_X1 U598 ( .A1(n5053), .A2(n6388), .B1(n447), .B2(n241), .ZN(n3221) );
  OAI22_X1 U599 ( .A1(n5021), .A2(n6385), .B1(n447), .B2(n243), .ZN(n3222) );
  OAI22_X1 U600 ( .A1(n4989), .A2(n6383), .B1(n447), .B2(n245), .ZN(n3223) );
  OAI22_X1 U601 ( .A1(n4957), .A2(n6382), .B1(n447), .B2(n247), .ZN(n3224) );
  OAI22_X1 U602 ( .A1(n4925), .A2(n6380), .B1(n447), .B2(n249), .ZN(n3225) );
  OAI22_X1 U603 ( .A1(n4893), .A2(n6384), .B1(n447), .B2(n251), .ZN(n3226) );
  OAI22_X1 U604 ( .A1(n4861), .A2(n6381), .B1(n447), .B2(n253), .ZN(n3227) );
  OAI22_X1 U605 ( .A1(n4829), .A2(n6387), .B1(n447), .B2(n255), .ZN(n3228) );
  OAI22_X1 U606 ( .A1(n4797), .A2(n6386), .B1(n447), .B2(n257), .ZN(n3229) );
  OAI22_X1 U607 ( .A1(n4765), .A2(n6392), .B1(n447), .B2(n259), .ZN(n3230) );
  OAI22_X1 U608 ( .A1(n4733), .A2(n6394), .B1(n447), .B2(n261), .ZN(n3231) );
  OAI22_X1 U609 ( .A1(n4701), .A2(n6389), .B1(n447), .B2(n263), .ZN(n3232) );
  OAI22_X1 U610 ( .A1(n4669), .A2(n6395), .B1(n447), .B2(n265), .ZN(n3233) );
  OAI22_X1 U611 ( .A1(n4637), .A2(n6400), .B1(n447), .B2(n267), .ZN(n3234) );
  OAI22_X1 U612 ( .A1(n4605), .A2(n6402), .B1(n447), .B2(n269), .ZN(n3235) );
  OAI22_X1 U613 ( .A1(n4573), .A2(n6397), .B1(n447), .B2(n271), .ZN(n3236) );
  OAI22_X1 U614 ( .A1(n4541), .A2(n6403), .B1(n447), .B2(n273), .ZN(n3237) );
  OAI22_X1 U615 ( .A1(n4509), .A2(n6408), .B1(n447), .B2(n275), .ZN(n3238) );
  OAI22_X1 U616 ( .A1(n4477), .A2(n6405), .B1(n447), .B2(n277), .ZN(n3239) );
  OAI22_X1 U617 ( .A1(n4445), .A2(n6411), .B1(n447), .B2(n279), .ZN(n3240) );
  OAI221_X1 U619 ( .B1(n5944), .B2(n281), .C1(n5710), .C2(n5506), .A(n282), 
        .ZN(n459) );
  OAI22_X1 U620 ( .A1(n5506), .A2(net54885), .B1(net54923), .B2(n446), .ZN(
        n3241) );
  INV_X1 U621 ( .A(n461), .ZN(n446) );
  OAI211_X1 U622 ( .C1(n5662), .C2(n321), .A(n462), .B(n463), .ZN(n461) );
  AOI222_X1 U623 ( .A1(n285), .A2(n464), .B1(\UUT/Mpath/out_jar[16] ), .B2(
        n325), .C1(n284), .C2(n465), .ZN(n463) );
  INV_X1 U624 ( .A(n5702), .ZN(n465) );
  AOI22_X1 U625 ( .A1(n6379), .A2(n6161), .B1(
        \UUT/Mpath/the_mult/x_mult_out[16] ), .B2(n291), .ZN(n462) );
  OAI221_X1 U626 ( .B1(n69), .B2(n466), .C1(n96), .C2(n71), .A(n467), .ZN(
        n3242) );
  NAND2_X1 U627 ( .A1(\UUT/Mpath/the_mult/x_operand2 [15]), .A2(n6409), .ZN(
        n467) );
  OAI222_X1 U630 ( .A1(n96), .A2(n123), .B1(n300), .B2(n466), .C1(
        \UUT/Mpath/the_alu/N54 ), .C2(net54891), .ZN(n3244) );
  INV_X1 U631 ( .A(n469), .ZN(n96) );
  OAI222_X1 U632 ( .A1(n470), .A2(n129), .B1(n471), .B2(n131), .C1(n5508), 
        .C2(n132), .ZN(n469) );
  OAI221_X1 U633 ( .B1(n133), .B2(n472), .C1(n5703), .C2(n135), .A(n473), .ZN(
        n3245) );
  AOI22_X1 U634 ( .A1(n137), .A2(n474), .B1(\UUT/Mpath/the_mult/Mad_out [47]), 
        .B2(n139), .ZN(n473) );
  OAI221_X1 U635 ( .B1(n140), .B2(n475), .C1(n5664), .C2(n142), .A(n476), .ZN(
        n3246) );
  AOI22_X1 U636 ( .A1(n144), .A2(n474), .B1(\UUT/Mpath/the_mult/Mad_out [15]), 
        .B2(n145), .ZN(n476) );
  INV_X1 U637 ( .A(n5665), .ZN(n474) );
  OAI22_X1 U638 ( .A1(net54905), .A2(n477), .B1(n5665), .B2(net54873), .ZN(
        n3247) );
  OAI221_X1 U639 ( .B1(n470), .B2(n310), .C1(n147), .C2(n477), .A(n478), .ZN(
        n3248) );
  AOI22_X1 U640 ( .A1(n312), .A2(n479), .B1(n314), .B2(n480), .ZN(n478) );
  INV_X1 U641 ( .A(\UUT/Mpath/the_mult/x_operand1[15] ), .ZN(n477) );
  OAI221_X1 U642 ( .B1(n470), .B2(n316), .C1(\UUT/Mpath/the_alu/N53 ), .C2(
        net54885), .A(n481), .ZN(n3249) );
  AOI22_X1 U643 ( .A1(n318), .A2(n479), .B1(n319), .B2(n480), .ZN(n481) );
  OAI22_X1 U644 ( .A1(n5406), .A2(n6407), .B1(n471), .B2(n219), .ZN(n3250) );
  OAI22_X1 U645 ( .A1(n5374), .A2(n6410), .B1(n471), .B2(n221), .ZN(n3251) );
  OAI22_X1 U646 ( .A1(n5342), .A2(n6401), .B1(n471), .B2(n223), .ZN(n3252) );
  OAI22_X1 U647 ( .A1(n5310), .A2(n6406), .B1(n471), .B2(n225), .ZN(n3253) );
  OAI22_X1 U648 ( .A1(n5278), .A2(n6399), .B1(n471), .B2(n227), .ZN(n3254) );
  OAI22_X1 U649 ( .A1(n5246), .A2(n6404), .B1(n471), .B2(n229), .ZN(n3255) );
  OAI22_X1 U650 ( .A1(n5214), .A2(n6398), .B1(n471), .B2(n231), .ZN(n3256) );
  OAI22_X1 U651 ( .A1(n5182), .A2(n6396), .B1(n471), .B2(n233), .ZN(n3257) );
  OAI22_X1 U652 ( .A1(n5150), .A2(n6393), .B1(n471), .B2(n235), .ZN(n3258) );
  OAI22_X1 U653 ( .A1(n5118), .A2(n6391), .B1(n471), .B2(n237), .ZN(n3259) );
  OAI22_X1 U654 ( .A1(n5086), .A2(n6390), .B1(n471), .B2(n239), .ZN(n3260) );
  OAI22_X1 U655 ( .A1(n5054), .A2(n6388), .B1(n471), .B2(n241), .ZN(n3261) );
  OAI22_X1 U656 ( .A1(n5022), .A2(n6385), .B1(n471), .B2(n243), .ZN(n3262) );
  OAI22_X1 U657 ( .A1(n4990), .A2(n6383), .B1(n471), .B2(n245), .ZN(n3263) );
  OAI22_X1 U658 ( .A1(n4958), .A2(n6382), .B1(n471), .B2(n247), .ZN(n3264) );
  OAI22_X1 U659 ( .A1(n4926), .A2(n6380), .B1(n471), .B2(n249), .ZN(n3265) );
  OAI22_X1 U660 ( .A1(n4894), .A2(n6384), .B1(n471), .B2(n251), .ZN(n3266) );
  OAI22_X1 U661 ( .A1(n4862), .A2(n6381), .B1(n471), .B2(n253), .ZN(n3267) );
  OAI22_X1 U662 ( .A1(n4830), .A2(n6387), .B1(n471), .B2(n255), .ZN(n3268) );
  OAI22_X1 U663 ( .A1(n4798), .A2(n6386), .B1(n471), .B2(n257), .ZN(n3269) );
  OAI22_X1 U664 ( .A1(n4766), .A2(n6392), .B1(n471), .B2(n259), .ZN(n3270) );
  OAI22_X1 U665 ( .A1(n4734), .A2(n6394), .B1(n471), .B2(n261), .ZN(n3271) );
  OAI22_X1 U666 ( .A1(n4702), .A2(n6389), .B1(n471), .B2(n263), .ZN(n3272) );
  OAI22_X1 U667 ( .A1(n4670), .A2(n6395), .B1(n471), .B2(n265), .ZN(n3273) );
  OAI22_X1 U668 ( .A1(n4638), .A2(n6400), .B1(n471), .B2(n267), .ZN(n3274) );
  OAI22_X1 U669 ( .A1(n4606), .A2(n6402), .B1(n471), .B2(n269), .ZN(n3275) );
  OAI22_X1 U670 ( .A1(n4574), .A2(n6397), .B1(n471), .B2(n271), .ZN(n3276) );
  OAI22_X1 U671 ( .A1(n4542), .A2(n6403), .B1(n471), .B2(n273), .ZN(n3277) );
  OAI22_X1 U672 ( .A1(n4510), .A2(n6408), .B1(n471), .B2(n275), .ZN(n3278) );
  OAI22_X1 U673 ( .A1(n4478), .A2(n6405), .B1(n471), .B2(n277), .ZN(n3279) );
  OAI22_X1 U674 ( .A1(n4446), .A2(n6411), .B1(n471), .B2(n279), .ZN(n3280) );
  OAI211_X1 U676 ( .C1(n482), .C2(n483), .A(n484), .B(n485), .ZN(n480) );
  AOI22_X1 U677 ( .A1(n486), .A2(n487), .B1(n488), .B2(n489), .ZN(n485) );
  INV_X1 U678 ( .A(n5509), .ZN(n488) );
  INV_X1 U679 ( .A(n5756), .ZN(n483) );
  OAI22_X1 U680 ( .A1(n5509), .A2(net54883), .B1(net54921), .B2(n470), .ZN(
        n3281) );
  INV_X1 U681 ( .A(n490), .ZN(n470) );
  OAI211_X1 U682 ( .C1(n5664), .C2(n321), .A(n491), .B(n492), .ZN(n490) );
  AOI222_X1 U683 ( .A1(n285), .A2(n493), .B1(\UUT/Mpath/out_jar[15] ), .B2(
        n325), .C1(n284), .C2(n494), .ZN(n492) );
  INV_X1 U684 ( .A(n5703), .ZN(n494) );
  AOI22_X1 U685 ( .A1(n6379), .A2(n6169), .B1(
        \UUT/Mpath/the_mult/x_mult_out[15] ), .B2(n291), .ZN(n491) );
  OAI221_X1 U686 ( .B1(n495), .B2(n69), .C1(n95), .C2(n71), .A(n496), .ZN(
        n3282) );
  NAND2_X1 U687 ( .A1(\UUT/Mpath/the_mult/x_operand2 [14]), .A2(n6409), .ZN(
        n496) );
  OAI222_X1 U690 ( .A1(n95), .A2(n123), .B1(n495), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N56 ), .C2(net54891), .ZN(n3284) );
  INV_X1 U691 ( .A(\UUT/break_code[14] ), .ZN(n495) );
  INV_X1 U692 ( .A(n498), .ZN(n95) );
  OAI222_X1 U693 ( .A1(n499), .A2(n129), .B1(n500), .B2(n131), .C1(n5511), 
        .C2(n132), .ZN(n498) );
  OAI221_X1 U694 ( .B1(n133), .B2(n501), .C1(n5704), .C2(n135), .A(n502), .ZN(
        n3285) );
  AOI22_X1 U695 ( .A1(n137), .A2(n503), .B1(\UUT/Mpath/the_mult/Mad_out [46]), 
        .B2(n139), .ZN(n502) );
  OAI221_X1 U696 ( .B1(n140), .B2(n504), .C1(n5666), .C2(n142), .A(n505), .ZN(
        n3286) );
  AOI22_X1 U697 ( .A1(n144), .A2(n503), .B1(\UUT/Mpath/the_mult/Mad_out [14]), 
        .B2(n145), .ZN(n505) );
  INV_X1 U698 ( .A(n5667), .ZN(n503) );
  OAI22_X1 U699 ( .A1(net54905), .A2(n506), .B1(n5667), .B2(net54873), .ZN(
        n3287) );
  OAI221_X1 U700 ( .B1(n499), .B2(n310), .C1(n147), .C2(n506), .A(n507), .ZN(
        n3288) );
  AOI22_X1 U701 ( .A1(n312), .A2(n508), .B1(n314), .B2(n509), .ZN(n507) );
  INV_X1 U702 ( .A(\UUT/Mpath/the_mult/x_operand1[14] ), .ZN(n506) );
  OAI221_X1 U703 ( .B1(n499), .B2(n316), .C1(\UUT/Mpath/the_alu/N55 ), .C2(
        net54885), .A(n510), .ZN(n3289) );
  AOI22_X1 U704 ( .A1(n318), .A2(n508), .B1(n319), .B2(n509), .ZN(n510) );
  OAI22_X1 U705 ( .A1(n5407), .A2(n6407), .B1(n500), .B2(n219), .ZN(n3290) );
  OAI22_X1 U706 ( .A1(n5375), .A2(n6410), .B1(n500), .B2(n221), .ZN(n3291) );
  OAI22_X1 U707 ( .A1(n5343), .A2(n6401), .B1(n500), .B2(n223), .ZN(n3292) );
  OAI22_X1 U708 ( .A1(n5311), .A2(n6406), .B1(n500), .B2(n225), .ZN(n3293) );
  OAI22_X1 U709 ( .A1(n5279), .A2(n6399), .B1(n500), .B2(n227), .ZN(n3294) );
  OAI22_X1 U710 ( .A1(n5247), .A2(n6404), .B1(n500), .B2(n229), .ZN(n3295) );
  OAI22_X1 U711 ( .A1(n5215), .A2(n6398), .B1(n500), .B2(n231), .ZN(n3296) );
  OAI22_X1 U712 ( .A1(n5183), .A2(n6396), .B1(n500), .B2(n233), .ZN(n3297) );
  OAI22_X1 U713 ( .A1(n5151), .A2(n6393), .B1(n500), .B2(n235), .ZN(n3298) );
  OAI22_X1 U714 ( .A1(n5119), .A2(n6391), .B1(n500), .B2(n237), .ZN(n3299) );
  OAI22_X1 U715 ( .A1(n5087), .A2(n6390), .B1(n500), .B2(n239), .ZN(n3300) );
  OAI22_X1 U716 ( .A1(n5055), .A2(n6388), .B1(n500), .B2(n241), .ZN(n3301) );
  OAI22_X1 U717 ( .A1(n5023), .A2(n6385), .B1(n500), .B2(n243), .ZN(n3302) );
  OAI22_X1 U718 ( .A1(n4991), .A2(n6383), .B1(n500), .B2(n245), .ZN(n3303) );
  OAI22_X1 U719 ( .A1(n4959), .A2(n6382), .B1(n500), .B2(n247), .ZN(n3304) );
  OAI22_X1 U720 ( .A1(n4927), .A2(n6380), .B1(n500), .B2(n249), .ZN(n3305) );
  OAI22_X1 U721 ( .A1(n4895), .A2(n6384), .B1(n500), .B2(n251), .ZN(n3306) );
  OAI22_X1 U722 ( .A1(n4863), .A2(n6381), .B1(n500), .B2(n253), .ZN(n3307) );
  OAI22_X1 U723 ( .A1(n4831), .A2(n6387), .B1(n500), .B2(n255), .ZN(n3308) );
  OAI22_X1 U724 ( .A1(n4799), .A2(n6386), .B1(n500), .B2(n257), .ZN(n3309) );
  OAI22_X1 U725 ( .A1(n4767), .A2(n6392), .B1(n500), .B2(n259), .ZN(n3310) );
  OAI22_X1 U726 ( .A1(n4735), .A2(n6394), .B1(n500), .B2(n261), .ZN(n3311) );
  OAI22_X1 U727 ( .A1(n4703), .A2(n6389), .B1(n500), .B2(n263), .ZN(n3312) );
  OAI22_X1 U728 ( .A1(n4671), .A2(n6395), .B1(n500), .B2(n265), .ZN(n3313) );
  OAI22_X1 U729 ( .A1(n4639), .A2(n6400), .B1(n500), .B2(n267), .ZN(n3314) );
  OAI22_X1 U730 ( .A1(n4607), .A2(n6402), .B1(n500), .B2(n269), .ZN(n3315) );
  OAI22_X1 U731 ( .A1(n4575), .A2(n6397), .B1(n500), .B2(n271), .ZN(n3316) );
  OAI22_X1 U732 ( .A1(n4543), .A2(n6403), .B1(n500), .B2(n273), .ZN(n3317) );
  OAI22_X1 U733 ( .A1(n4511), .A2(n6408), .B1(n500), .B2(n275), .ZN(n3318) );
  OAI22_X1 U734 ( .A1(n4479), .A2(n6405), .B1(n500), .B2(n277), .ZN(n3319) );
  OAI22_X1 U735 ( .A1(n4447), .A2(n6411), .B1(n500), .B2(n279), .ZN(n3320) );
  OAI211_X1 U737 ( .C1(n482), .C2(n511), .A(n484), .B(n512), .ZN(n509) );
  AOI22_X1 U738 ( .A1(n486), .A2(n513), .B1(n514), .B2(n489), .ZN(n512) );
  INV_X1 U739 ( .A(n5512), .ZN(n514) );
  INV_X1 U740 ( .A(n5769), .ZN(n511) );
  OAI22_X1 U741 ( .A1(n5512), .A2(net54881), .B1(net54921), .B2(n499), .ZN(
        n3321) );
  INV_X1 U742 ( .A(n515), .ZN(n499) );
  OAI211_X1 U743 ( .C1(n5666), .C2(n321), .A(n516), .B(n517), .ZN(n515) );
  AOI222_X1 U744 ( .A1(n285), .A2(n518), .B1(\UUT/Mpath/out_jar[14] ), .B2(
        n325), .C1(n284), .C2(n519), .ZN(n517) );
  INV_X1 U745 ( .A(n5704), .ZN(n519) );
  AOI22_X1 U746 ( .A1(n6379), .A2(n6180), .B1(
        \UUT/Mpath/the_mult/x_mult_out[14] ), .B2(n291), .ZN(n516) );
  OAI221_X1 U747 ( .B1(n520), .B2(n69), .C1(n94), .C2(n71), .A(n521), .ZN(
        n3322) );
  NAND2_X1 U748 ( .A1(\UUT/Mpath/the_mult/x_operand2 [13]), .A2(n6409), .ZN(
        n521) );
  OAI222_X1 U751 ( .A1(n94), .A2(n123), .B1(n520), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N58 ), .C2(net54893), .ZN(n3324) );
  INV_X1 U752 ( .A(\UUT/break_code[13] ), .ZN(n520) );
  INV_X1 U753 ( .A(n523), .ZN(n94) );
  OAI222_X1 U754 ( .A1(n524), .A2(n129), .B1(n525), .B2(n131), .C1(n5514), 
        .C2(n132), .ZN(n523) );
  OAI221_X1 U755 ( .B1(n133), .B2(n526), .C1(n5705), .C2(n135), .A(n527), .ZN(
        n3325) );
  AOI22_X1 U756 ( .A1(n137), .A2(n528), .B1(\UUT/Mpath/the_mult/Mad_out [45]), 
        .B2(n139), .ZN(n527) );
  OAI221_X1 U757 ( .B1(n140), .B2(n529), .C1(n5668), .C2(n142), .A(n530), .ZN(
        n3326) );
  AOI22_X1 U758 ( .A1(n144), .A2(n528), .B1(\UUT/Mpath/the_mult/Mad_out [13]), 
        .B2(n145), .ZN(n530) );
  INV_X1 U759 ( .A(n5669), .ZN(n528) );
  OAI22_X1 U760 ( .A1(net54905), .A2(n531), .B1(n5669), .B2(net54871), .ZN(
        n3327) );
  OAI221_X1 U761 ( .B1(n524), .B2(n310), .C1(n147), .C2(n531), .A(n532), .ZN(
        n3328) );
  AOI22_X1 U762 ( .A1(n312), .A2(n533), .B1(n314), .B2(n534), .ZN(n532) );
  INV_X1 U763 ( .A(\UUT/Mpath/the_mult/x_operand1[13] ), .ZN(n531) );
  OAI221_X1 U764 ( .B1(n524), .B2(n316), .C1(\UUT/Mpath/the_alu/N57 ), .C2(
        net54887), .A(n535), .ZN(n3329) );
  AOI22_X1 U765 ( .A1(n318), .A2(n533), .B1(n319), .B2(n534), .ZN(n535) );
  OAI22_X1 U766 ( .A1(n5408), .A2(n6407), .B1(n525), .B2(n219), .ZN(n3330) );
  OAI22_X1 U767 ( .A1(n5376), .A2(n6410), .B1(n525), .B2(n221), .ZN(n3331) );
  OAI22_X1 U768 ( .A1(n5344), .A2(n6401), .B1(n525), .B2(n223), .ZN(n3332) );
  OAI22_X1 U769 ( .A1(n5312), .A2(n6406), .B1(n525), .B2(n225), .ZN(n3333) );
  OAI22_X1 U770 ( .A1(n5280), .A2(n6399), .B1(n525), .B2(n227), .ZN(n3334) );
  OAI22_X1 U771 ( .A1(n5248), .A2(n6404), .B1(n525), .B2(n229), .ZN(n3335) );
  OAI22_X1 U772 ( .A1(n5216), .A2(n6398), .B1(n525), .B2(n231), .ZN(n3336) );
  OAI22_X1 U773 ( .A1(n5184), .A2(n6396), .B1(n525), .B2(n233), .ZN(n3337) );
  OAI22_X1 U774 ( .A1(n5152), .A2(n6393), .B1(n525), .B2(n235), .ZN(n3338) );
  OAI22_X1 U775 ( .A1(n5120), .A2(n6391), .B1(n525), .B2(n237), .ZN(n3339) );
  OAI22_X1 U776 ( .A1(n5088), .A2(n6390), .B1(n525), .B2(n239), .ZN(n3340) );
  OAI22_X1 U777 ( .A1(n5056), .A2(n6388), .B1(n525), .B2(n241), .ZN(n3341) );
  OAI22_X1 U778 ( .A1(n5024), .A2(n6385), .B1(n525), .B2(n243), .ZN(n3342) );
  OAI22_X1 U779 ( .A1(n4992), .A2(n6383), .B1(n525), .B2(n245), .ZN(n3343) );
  OAI22_X1 U780 ( .A1(n4960), .A2(n6382), .B1(n525), .B2(n247), .ZN(n3344) );
  OAI22_X1 U781 ( .A1(n4928), .A2(n6380), .B1(n525), .B2(n249), .ZN(n3345) );
  OAI22_X1 U782 ( .A1(n4896), .A2(n6384), .B1(n525), .B2(n251), .ZN(n3346) );
  OAI22_X1 U783 ( .A1(n4864), .A2(n6381), .B1(n525), .B2(n253), .ZN(n3347) );
  OAI22_X1 U784 ( .A1(n4832), .A2(n6387), .B1(n525), .B2(n255), .ZN(n3348) );
  OAI22_X1 U785 ( .A1(n4800), .A2(n6386), .B1(n525), .B2(n257), .ZN(n3349) );
  OAI22_X1 U786 ( .A1(n4768), .A2(n6392), .B1(n525), .B2(n259), .ZN(n3350) );
  OAI22_X1 U787 ( .A1(n4736), .A2(n6394), .B1(n525), .B2(n261), .ZN(n3351) );
  OAI22_X1 U788 ( .A1(n4704), .A2(n6389), .B1(n525), .B2(n263), .ZN(n3352) );
  OAI22_X1 U789 ( .A1(n4672), .A2(n6395), .B1(n525), .B2(n265), .ZN(n3353) );
  OAI22_X1 U790 ( .A1(n4640), .A2(n6400), .B1(n525), .B2(n267), .ZN(n3354) );
  OAI22_X1 U791 ( .A1(n4608), .A2(n6402), .B1(n525), .B2(n269), .ZN(n3355) );
  OAI22_X1 U792 ( .A1(n4576), .A2(n6397), .B1(n525), .B2(n271), .ZN(n3356) );
  OAI22_X1 U793 ( .A1(n4544), .A2(n6403), .B1(n525), .B2(n273), .ZN(n3357) );
  OAI22_X1 U794 ( .A1(n4512), .A2(n6408), .B1(n525), .B2(n275), .ZN(n3358) );
  OAI22_X1 U795 ( .A1(n4480), .A2(n6405), .B1(n525), .B2(n277), .ZN(n3359) );
  OAI22_X1 U796 ( .A1(n4448), .A2(n6411), .B1(n525), .B2(n279), .ZN(n3360) );
  OAI211_X1 U798 ( .C1(n482), .C2(n536), .A(n484), .B(n537), .ZN(n534) );
  AOI22_X1 U799 ( .A1(n486), .A2(n538), .B1(n539), .B2(n489), .ZN(n537) );
  INV_X1 U800 ( .A(n5515), .ZN(n539) );
  INV_X1 U801 ( .A(n5786), .ZN(n536) );
  OAI22_X1 U802 ( .A1(n5515), .A2(net54883), .B1(net54925), .B2(n524), .ZN(
        n3361) );
  INV_X1 U803 ( .A(n540), .ZN(n524) );
  OAI211_X1 U804 ( .C1(n5668), .C2(n321), .A(n541), .B(n542), .ZN(n540) );
  AOI222_X1 U805 ( .A1(n285), .A2(n543), .B1(\UUT/Mpath/out_jar[13] ), .B2(
        n325), .C1(n284), .C2(n544), .ZN(n542) );
  INV_X1 U806 ( .A(n5705), .ZN(n544) );
  AOI22_X1 U807 ( .A1(n6379), .A2(n6187), .B1(
        \UUT/Mpath/the_mult/x_mult_out[13] ), .B2(n291), .ZN(n541) );
  OAI22_X1 U808 ( .A1(n545), .A2(n546), .B1(n295), .B2(n2668), .ZN(n3362) );
  OAI221_X1 U809 ( .B1(n547), .B2(n69), .C1(n93), .C2(n71), .A(n548), .ZN(
        n3363) );
  NAND2_X1 U810 ( .A1(\UUT/Mpath/the_mult/x_operand2 [12]), .A2(n6409), .ZN(
        n548) );
  OAI222_X1 U811 ( .A1(n93), .A2(n123), .B1(n547), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N60 ), .C2(net54891), .ZN(n3364) );
  INV_X1 U812 ( .A(\UUT/break_code[12] ), .ZN(n547) );
  INV_X1 U813 ( .A(n549), .ZN(n93) );
  OAI222_X1 U814 ( .A1(n550), .A2(n129), .B1(n551), .B2(n131), .C1(n5517), 
        .C2(n132), .ZN(n549) );
  OAI221_X1 U815 ( .B1(n133), .B2(n552), .C1(n5706), .C2(n135), .A(n553), .ZN(
        n3365) );
  AOI22_X1 U816 ( .A1(n137), .A2(n554), .B1(\UUT/Mpath/the_mult/Mad_out [44]), 
        .B2(n139), .ZN(n553) );
  OAI221_X1 U817 ( .B1(n140), .B2(n555), .C1(n5670), .C2(n142), .A(n556), .ZN(
        n3366) );
  AOI22_X1 U818 ( .A1(n144), .A2(n554), .B1(\UUT/Mpath/the_mult/Mad_out [12]), 
        .B2(n145), .ZN(n556) );
  INV_X1 U819 ( .A(n5671), .ZN(n554) );
  OAI22_X1 U820 ( .A1(net54909), .A2(n557), .B1(n5671), .B2(net54871), .ZN(
        n3367) );
  OAI221_X1 U821 ( .B1(n550), .B2(n310), .C1(n147), .C2(n557), .A(n558), .ZN(
        n3368) );
  AOI22_X1 U822 ( .A1(n312), .A2(n559), .B1(n314), .B2(n560), .ZN(n558) );
  INV_X1 U823 ( .A(\UUT/Mpath/the_mult/x_operand1[12] ), .ZN(n557) );
  OAI221_X1 U824 ( .B1(n550), .B2(n316), .C1(\UUT/Mpath/the_alu/N59 ), .C2(
        net54887), .A(n561), .ZN(n3369) );
  AOI22_X1 U825 ( .A1(n318), .A2(n559), .B1(n319), .B2(n560), .ZN(n561) );
  OAI22_X1 U826 ( .A1(n5409), .A2(n6407), .B1(n551), .B2(n219), .ZN(n3370) );
  OAI22_X1 U827 ( .A1(n5377), .A2(n6410), .B1(n551), .B2(n221), .ZN(n3371) );
  OAI22_X1 U828 ( .A1(n5345), .A2(n6401), .B1(n551), .B2(n223), .ZN(n3372) );
  OAI22_X1 U829 ( .A1(n5313), .A2(n6406), .B1(n551), .B2(n225), .ZN(n3373) );
  OAI22_X1 U830 ( .A1(n5281), .A2(n6399), .B1(n551), .B2(n227), .ZN(n3374) );
  OAI22_X1 U831 ( .A1(n5249), .A2(n6404), .B1(n551), .B2(n229), .ZN(n3375) );
  OAI22_X1 U832 ( .A1(n5217), .A2(n6398), .B1(n551), .B2(n231), .ZN(n3376) );
  OAI22_X1 U833 ( .A1(n5185), .A2(n6396), .B1(n551), .B2(n233), .ZN(n3377) );
  OAI22_X1 U834 ( .A1(n5153), .A2(n6393), .B1(n551), .B2(n235), .ZN(n3378) );
  OAI22_X1 U835 ( .A1(n5121), .A2(n6391), .B1(n551), .B2(n237), .ZN(n3379) );
  OAI22_X1 U836 ( .A1(n5089), .A2(n6390), .B1(n551), .B2(n239), .ZN(n3380) );
  OAI22_X1 U837 ( .A1(n5057), .A2(n6388), .B1(n551), .B2(n241), .ZN(n3381) );
  OAI22_X1 U838 ( .A1(n5025), .A2(n6385), .B1(n551), .B2(n243), .ZN(n3382) );
  OAI22_X1 U839 ( .A1(n4993), .A2(n6383), .B1(n551), .B2(n245), .ZN(n3383) );
  OAI22_X1 U840 ( .A1(n4961), .A2(n6382), .B1(n551), .B2(n247), .ZN(n3384) );
  OAI22_X1 U841 ( .A1(n4929), .A2(n6380), .B1(n551), .B2(n249), .ZN(n3385) );
  OAI22_X1 U842 ( .A1(n4897), .A2(n6384), .B1(n551), .B2(n251), .ZN(n3386) );
  OAI22_X1 U843 ( .A1(n4865), .A2(n6381), .B1(n551), .B2(n253), .ZN(n3387) );
  OAI22_X1 U844 ( .A1(n4833), .A2(n6387), .B1(n551), .B2(n255), .ZN(n3388) );
  OAI22_X1 U845 ( .A1(n4801), .A2(n6386), .B1(n551), .B2(n257), .ZN(n3389) );
  OAI22_X1 U846 ( .A1(n4769), .A2(n6392), .B1(n551), .B2(n259), .ZN(n3390) );
  OAI22_X1 U847 ( .A1(n4737), .A2(n6394), .B1(n551), .B2(n261), .ZN(n3391) );
  OAI22_X1 U848 ( .A1(n4705), .A2(n6389), .B1(n551), .B2(n263), .ZN(n3392) );
  OAI22_X1 U849 ( .A1(n4673), .A2(n6395), .B1(n551), .B2(n265), .ZN(n3393) );
  OAI22_X1 U850 ( .A1(n4641), .A2(n6400), .B1(n551), .B2(n267), .ZN(n3394) );
  OAI22_X1 U851 ( .A1(n4609), .A2(n6402), .B1(n551), .B2(n269), .ZN(n3395) );
  OAI22_X1 U852 ( .A1(n4577), .A2(n6397), .B1(n551), .B2(n271), .ZN(n3396) );
  OAI22_X1 U853 ( .A1(n4545), .A2(n6403), .B1(n551), .B2(n273), .ZN(n3397) );
  OAI22_X1 U854 ( .A1(n4513), .A2(n6408), .B1(n551), .B2(n275), .ZN(n3398) );
  OAI22_X1 U855 ( .A1(n4481), .A2(n6405), .B1(n551), .B2(n277), .ZN(n3399) );
  OAI22_X1 U856 ( .A1(n4449), .A2(n6411), .B1(n551), .B2(n279), .ZN(n3400) );
  OAI211_X1 U858 ( .C1(n482), .C2(n562), .A(n484), .B(n563), .ZN(n560) );
  AOI22_X1 U859 ( .A1(n486), .A2(n564), .B1(n565), .B2(n489), .ZN(n563) );
  INV_X1 U860 ( .A(n5518), .ZN(n565) );
  INV_X1 U861 ( .A(n5799), .ZN(n562) );
  OAI22_X1 U862 ( .A1(n5518), .A2(net54883), .B1(net54921), .B2(n550), .ZN(
        n3401) );
  INV_X1 U863 ( .A(n566), .ZN(n550) );
  OAI211_X1 U864 ( .C1(n5670), .C2(n321), .A(n567), .B(n568), .ZN(n566) );
  AOI222_X1 U865 ( .A1(n285), .A2(n569), .B1(\UUT/Mpath/out_jar[12] ), .B2(
        n325), .C1(n284), .C2(n570), .ZN(n568) );
  INV_X1 U866 ( .A(n5706), .ZN(n570) );
  AOI22_X1 U867 ( .A1(n6379), .A2(n6203), .B1(
        \UUT/Mpath/the_mult/x_mult_out[12] ), .B2(n291), .ZN(n567) );
  OAI22_X1 U868 ( .A1(n571), .A2(n546), .B1(n295), .B2(n2671), .ZN(n3402) );
  OAI221_X1 U869 ( .B1(n572), .B2(n69), .C1(n92), .C2(n71), .A(n573), .ZN(
        n3403) );
  NAND2_X1 U870 ( .A1(\UUT/Mpath/the_mult/x_operand2 [11]), .A2(n6409), .ZN(
        n573) );
  OAI222_X1 U871 ( .A1(n92), .A2(n123), .B1(n572), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N62 ), .C2(net54891), .ZN(n3404) );
  INV_X1 U872 ( .A(\UUT/break_code[11] ), .ZN(n572) );
  INV_X1 U873 ( .A(n574), .ZN(n92) );
  OAI222_X1 U874 ( .A1(n575), .A2(n129), .B1(n576), .B2(n131), .C1(n5520), 
        .C2(n132), .ZN(n574) );
  OAI221_X1 U875 ( .B1(n133), .B2(n577), .C1(n5707), .C2(n135), .A(n578), .ZN(
        n3405) );
  AOI22_X1 U876 ( .A1(n137), .A2(n579), .B1(\UUT/Mpath/the_mult/Mad_out [43]), 
        .B2(n139), .ZN(n578) );
  OAI221_X1 U877 ( .B1(n140), .B2(n580), .C1(n5672), .C2(n142), .A(n581), .ZN(
        n3406) );
  AOI22_X1 U878 ( .A1(n144), .A2(n579), .B1(\UUT/Mpath/the_mult/Mad_out [11]), 
        .B2(n145), .ZN(n581) );
  INV_X1 U879 ( .A(n5673), .ZN(n579) );
  OAI22_X1 U880 ( .A1(net54907), .A2(n582), .B1(n5673), .B2(net54873), .ZN(
        n3407) );
  OAI221_X1 U881 ( .B1(n575), .B2(n310), .C1(n147), .C2(n582), .A(n583), .ZN(
        n3408) );
  AOI22_X1 U882 ( .A1(n312), .A2(n584), .B1(n314), .B2(n585), .ZN(n583) );
  INV_X1 U883 ( .A(\UUT/Mpath/the_mult/x_operand1[11] ), .ZN(n582) );
  OAI221_X1 U884 ( .B1(n575), .B2(n316), .C1(\UUT/Mpath/the_alu/N61 ), .C2(
        net54887), .A(n586), .ZN(n3409) );
  AOI22_X1 U885 ( .A1(n318), .A2(n584), .B1(n319), .B2(n585), .ZN(n586) );
  OAI22_X1 U886 ( .A1(n5410), .A2(n6407), .B1(n576), .B2(n219), .ZN(n3410) );
  OAI22_X1 U887 ( .A1(n5378), .A2(n6410), .B1(n576), .B2(n221), .ZN(n3411) );
  OAI22_X1 U888 ( .A1(n5346), .A2(n6401), .B1(n576), .B2(n223), .ZN(n3412) );
  OAI22_X1 U889 ( .A1(n5314), .A2(n6406), .B1(n576), .B2(n225), .ZN(n3413) );
  OAI22_X1 U890 ( .A1(n5282), .A2(n6399), .B1(n576), .B2(n227), .ZN(n3414) );
  OAI22_X1 U891 ( .A1(n5250), .A2(n6404), .B1(n576), .B2(n229), .ZN(n3415) );
  OAI22_X1 U892 ( .A1(n5218), .A2(n6398), .B1(n576), .B2(n231), .ZN(n3416) );
  OAI22_X1 U893 ( .A1(n5186), .A2(n6396), .B1(n576), .B2(n233), .ZN(n3417) );
  OAI22_X1 U894 ( .A1(n5154), .A2(n6393), .B1(n576), .B2(n235), .ZN(n3418) );
  OAI22_X1 U895 ( .A1(n5122), .A2(n6391), .B1(n576), .B2(n237), .ZN(n3419) );
  OAI22_X1 U896 ( .A1(n5090), .A2(n6390), .B1(n576), .B2(n239), .ZN(n3420) );
  OAI22_X1 U897 ( .A1(n5058), .A2(n6388), .B1(n576), .B2(n241), .ZN(n3421) );
  OAI22_X1 U898 ( .A1(n5026), .A2(n6385), .B1(n576), .B2(n243), .ZN(n3422) );
  OAI22_X1 U899 ( .A1(n4994), .A2(n6383), .B1(n576), .B2(n245), .ZN(n3423) );
  OAI22_X1 U900 ( .A1(n4962), .A2(n6382), .B1(n576), .B2(n247), .ZN(n3424) );
  OAI22_X1 U901 ( .A1(n4930), .A2(n6380), .B1(n576), .B2(n249), .ZN(n3425) );
  OAI22_X1 U902 ( .A1(n4898), .A2(n6384), .B1(n576), .B2(n251), .ZN(n3426) );
  OAI22_X1 U903 ( .A1(n4866), .A2(n6381), .B1(n576), .B2(n253), .ZN(n3427) );
  OAI22_X1 U904 ( .A1(n4834), .A2(n6387), .B1(n576), .B2(n255), .ZN(n3428) );
  OAI22_X1 U905 ( .A1(n4802), .A2(n6386), .B1(n576), .B2(n257), .ZN(n3429) );
  OAI22_X1 U906 ( .A1(n4770), .A2(n6392), .B1(n576), .B2(n259), .ZN(n3430) );
  OAI22_X1 U907 ( .A1(n4738), .A2(n6394), .B1(n576), .B2(n261), .ZN(n3431) );
  OAI22_X1 U908 ( .A1(n4706), .A2(n6389), .B1(n576), .B2(n263), .ZN(n3432) );
  OAI22_X1 U909 ( .A1(n4674), .A2(n6395), .B1(n576), .B2(n265), .ZN(n3433) );
  OAI22_X1 U910 ( .A1(n4642), .A2(n6400), .B1(n576), .B2(n267), .ZN(n3434) );
  OAI22_X1 U911 ( .A1(n4610), .A2(n6402), .B1(n576), .B2(n269), .ZN(n3435) );
  OAI22_X1 U912 ( .A1(n4578), .A2(n6397), .B1(n576), .B2(n271), .ZN(n3436) );
  OAI22_X1 U913 ( .A1(n4546), .A2(n6403), .B1(n576), .B2(n273), .ZN(n3437) );
  OAI22_X1 U914 ( .A1(n4514), .A2(n6408), .B1(n576), .B2(n275), .ZN(n3438) );
  OAI22_X1 U915 ( .A1(n4482), .A2(n6405), .B1(n576), .B2(n277), .ZN(n3439) );
  OAI22_X1 U916 ( .A1(n4450), .A2(n6411), .B1(n576), .B2(n279), .ZN(n3440) );
  OAI211_X1 U918 ( .C1(n482), .C2(n587), .A(n484), .B(n588), .ZN(n585) );
  AOI22_X1 U919 ( .A1(n486), .A2(n589), .B1(n590), .B2(n489), .ZN(n588) );
  INV_X1 U920 ( .A(n5521), .ZN(n590) );
  INV_X1 U921 ( .A(n5812), .ZN(n587) );
  OAI22_X1 U922 ( .A1(n5521), .A2(net54883), .B1(net54921), .B2(n575), .ZN(
        n3441) );
  INV_X1 U923 ( .A(n591), .ZN(n575) );
  OAI211_X1 U924 ( .C1(n5672), .C2(n321), .A(n592), .B(n593), .ZN(n591) );
  AOI222_X1 U925 ( .A1(n285), .A2(n594), .B1(\UUT/Mpath/out_jar[11] ), .B2(
        n325), .C1(n284), .C2(n595), .ZN(n593) );
  INV_X1 U926 ( .A(n5707), .ZN(n595) );
  AOI22_X1 U927 ( .A1(n6379), .A2(n6204), .B1(
        \UUT/Mpath/the_mult/x_mult_out[11] ), .B2(n291), .ZN(n592) );
  OAI221_X1 U928 ( .B1(n133), .B2(n596), .C1(n5708), .C2(n135), .A(n597), .ZN(
        n3442) );
  AOI22_X1 U929 ( .A1(n137), .A2(n598), .B1(\UUT/Mpath/the_mult/Mad_out [42]), 
        .B2(n139), .ZN(n597) );
  OAI221_X1 U930 ( .B1(n140), .B2(n599), .C1(n5674), .C2(n142), .A(n600), .ZN(
        n3443) );
  AOI22_X1 U931 ( .A1(n144), .A2(n598), .B1(\UUT/Mpath/the_mult/Mad_out [10]), 
        .B2(n145), .ZN(n600) );
  INV_X1 U932 ( .A(n5675), .ZN(n598) );
  OAI22_X1 U933 ( .A1(net54907), .A2(n601), .B1(n5675), .B2(net54871), .ZN(
        n3444) );
  OAI221_X1 U934 ( .B1(n602), .B2(n310), .C1(n147), .C2(n601), .A(n603), .ZN(
        n3445) );
  AOI22_X1 U935 ( .A1(n312), .A2(n604), .B1(n314), .B2(n605), .ZN(n603) );
  INV_X1 U936 ( .A(\UUT/Mpath/the_mult/x_operand1[10] ), .ZN(n601) );
  OAI221_X1 U937 ( .B1(n602), .B2(n316), .C1(\UUT/Mpath/the_alu/N63 ), .C2(
        net54887), .A(n606), .ZN(n3446) );
  AOI22_X1 U938 ( .A1(n318), .A2(n604), .B1(n319), .B2(n605), .ZN(n606) );
  OAI22_X1 U939 ( .A1(n5524), .A2(net54883), .B1(net54923), .B2(n602), .ZN(
        n3447) );
  OAI221_X1 U940 ( .B1(n607), .B2(n69), .C1(n91), .C2(n71), .A(n608), .ZN(
        n3448) );
  NAND2_X1 U941 ( .A1(\UUT/Mpath/the_mult/x_operand2 [9]), .A2(n6409), .ZN(
        n608) );
  OAI222_X1 U942 ( .A1(n91), .A2(n123), .B1(n607), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N66 ), .C2(net54893), .ZN(n3449) );
  INV_X1 U943 ( .A(\UUT/break_code[9] ), .ZN(n607) );
  INV_X1 U944 ( .A(n609), .ZN(n91) );
  OAI222_X1 U945 ( .A1(n610), .A2(n129), .B1(n611), .B2(n131), .C1(n5431), 
        .C2(n132), .ZN(n609) );
  OAI221_X1 U946 ( .B1(n133), .B2(n612), .C1(n5678), .C2(n135), .A(n613), .ZN(
        n3450) );
  AOI22_X1 U947 ( .A1(n137), .A2(n614), .B1(\UUT/Mpath/the_mult/Mad_out [41]), 
        .B2(n139), .ZN(n613) );
  OAI221_X1 U948 ( .B1(n140), .B2(n615), .C1(n5614), .C2(n142), .A(n616), .ZN(
        n3451) );
  AOI22_X1 U949 ( .A1(n144), .A2(n614), .B1(\UUT/Mpath/the_mult/Mad_out [9]), 
        .B2(n145), .ZN(n616) );
  INV_X1 U950 ( .A(n5615), .ZN(n614) );
  OAI22_X1 U951 ( .A1(net54907), .A2(n617), .B1(n5615), .B2(net54871), .ZN(
        n3452) );
  OAI221_X1 U952 ( .B1(n610), .B2(n310), .C1(n147), .C2(n617), .A(n618), .ZN(
        n3453) );
  AOI22_X1 U953 ( .A1(n312), .A2(n619), .B1(n314), .B2(n620), .ZN(n618) );
  INV_X1 U954 ( .A(\UUT/Mpath/the_mult/x_operand1[9] ), .ZN(n617) );
  OAI221_X1 U955 ( .B1(n610), .B2(n316), .C1(\UUT/Mpath/the_alu/N65 ), .C2(
        net54889), .A(n621), .ZN(n3454) );
  AOI22_X1 U956 ( .A1(n318), .A2(n619), .B1(n319), .B2(n620), .ZN(n621) );
  OAI22_X1 U957 ( .A1(n5381), .A2(n6407), .B1(n611), .B2(n219), .ZN(n3455) );
  OAI22_X1 U958 ( .A1(n5349), .A2(n6410), .B1(n611), .B2(n221), .ZN(n3456) );
  OAI22_X1 U959 ( .A1(n5317), .A2(n6401), .B1(n611), .B2(n223), .ZN(n3457) );
  OAI22_X1 U960 ( .A1(n5285), .A2(n6406), .B1(n611), .B2(n225), .ZN(n3458) );
  OAI22_X1 U961 ( .A1(n5253), .A2(n6399), .B1(n611), .B2(n227), .ZN(n3459) );
  OAI22_X1 U962 ( .A1(n5221), .A2(n6404), .B1(n611), .B2(n229), .ZN(n3460) );
  OAI22_X1 U963 ( .A1(n5189), .A2(n6398), .B1(n611), .B2(n231), .ZN(n3461) );
  OAI22_X1 U964 ( .A1(n5157), .A2(n6396), .B1(n611), .B2(n233), .ZN(n3462) );
  OAI22_X1 U965 ( .A1(n5125), .A2(n6393), .B1(n611), .B2(n235), .ZN(n3463) );
  OAI22_X1 U966 ( .A1(n5093), .A2(n6391), .B1(n611), .B2(n237), .ZN(n3464) );
  OAI22_X1 U967 ( .A1(n5061), .A2(n6390), .B1(n611), .B2(n239), .ZN(n3465) );
  OAI22_X1 U968 ( .A1(n5029), .A2(n6388), .B1(n611), .B2(n241), .ZN(n3466) );
  OAI22_X1 U969 ( .A1(n4997), .A2(n6385), .B1(n611), .B2(n243), .ZN(n3467) );
  OAI22_X1 U970 ( .A1(n4965), .A2(n6383), .B1(n611), .B2(n245), .ZN(n3468) );
  OAI22_X1 U971 ( .A1(n4933), .A2(n6382), .B1(n611), .B2(n247), .ZN(n3469) );
  OAI22_X1 U972 ( .A1(n4901), .A2(n6380), .B1(n611), .B2(n249), .ZN(n3470) );
  OAI22_X1 U973 ( .A1(n4869), .A2(n6384), .B1(n611), .B2(n251), .ZN(n3471) );
  OAI22_X1 U974 ( .A1(n4837), .A2(n6381), .B1(n611), .B2(n253), .ZN(n3472) );
  OAI22_X1 U975 ( .A1(n4805), .A2(n6387), .B1(n611), .B2(n255), .ZN(n3473) );
  OAI22_X1 U976 ( .A1(n4773), .A2(n6386), .B1(n611), .B2(n257), .ZN(n3474) );
  OAI22_X1 U977 ( .A1(n4741), .A2(n6392), .B1(n611), .B2(n259), .ZN(n3475) );
  OAI22_X1 U978 ( .A1(n4709), .A2(n6394), .B1(n611), .B2(n261), .ZN(n3476) );
  OAI22_X1 U979 ( .A1(n4677), .A2(n6389), .B1(n611), .B2(n263), .ZN(n3477) );
  OAI22_X1 U980 ( .A1(n4645), .A2(n6395), .B1(n611), .B2(n265), .ZN(n3478) );
  OAI22_X1 U981 ( .A1(n4613), .A2(n6400), .B1(n611), .B2(n267), .ZN(n3479) );
  OAI22_X1 U982 ( .A1(n4581), .A2(n6402), .B1(n611), .B2(n269), .ZN(n3480) );
  OAI22_X1 U983 ( .A1(n4549), .A2(n6397), .B1(n611), .B2(n271), .ZN(n3481) );
  OAI22_X1 U984 ( .A1(n4517), .A2(n6403), .B1(n611), .B2(n273), .ZN(n3482) );
  OAI22_X1 U985 ( .A1(n4485), .A2(n6408), .B1(n611), .B2(n275), .ZN(n3483) );
  OAI22_X1 U986 ( .A1(n4453), .A2(n6405), .B1(n611), .B2(n277), .ZN(n3484) );
  OAI22_X1 U987 ( .A1(n4421), .A2(n6411), .B1(n611), .B2(n279), .ZN(n3485) );
  OAI211_X1 U989 ( .C1(n482), .C2(n622), .A(n484), .B(n623), .ZN(n620) );
  AOI22_X1 U990 ( .A1(n486), .A2(n624), .B1(n625), .B2(n489), .ZN(n623) );
  INV_X1 U991 ( .A(n5433), .ZN(n625) );
  INV_X1 U992 ( .A(n5712), .ZN(n622) );
  OAI22_X1 U993 ( .A1(n5433), .A2(net54877), .B1(net54923), .B2(n610), .ZN(
        n3486) );
  INV_X1 U994 ( .A(n626), .ZN(n610) );
  OAI211_X1 U995 ( .C1(n5614), .C2(n321), .A(n627), .B(n628), .ZN(n626) );
  AOI222_X1 U996 ( .A1(n285), .A2(n629), .B1(\UUT/Mpath/out_jar[9] ), .B2(n325), .C1(n284), .C2(n630), .ZN(n628) );
  INV_X1 U997 ( .A(n5678), .ZN(n630) );
  AOI22_X1 U998 ( .A1(n6379), .A2(n6189), .B1(
        \UUT/Mpath/the_mult/x_mult_out[9] ), .B2(n291), .ZN(n627) );
  OAI22_X1 U999 ( .A1(n631), .A2(n546), .B1(n295), .B2(n2677), .ZN(n3487) );
  OAI221_X1 U1000 ( .B1(n133), .B2(n632), .C1(n5679), .C2(n135), .A(n633), 
        .ZN(n3488) );
  AOI22_X1 U1001 ( .A1(n137), .A2(n634), .B1(\UUT/Mpath/the_mult/Mad_out [40]), 
        .B2(n139), .ZN(n633) );
  OAI221_X1 U1002 ( .B1(n140), .B2(n635), .C1(n5616), .C2(n142), .A(n636), 
        .ZN(n3489) );
  AOI22_X1 U1003 ( .A1(n144), .A2(n634), .B1(\UUT/Mpath/the_mult/Mad_out [8]), 
        .B2(n145), .ZN(n636) );
  INV_X1 U1004 ( .A(n5617), .ZN(n634) );
  OAI22_X1 U1005 ( .A1(net54907), .A2(n637), .B1(n5617), .B2(net54875), .ZN(
        n3490) );
  OAI221_X1 U1006 ( .B1(n638), .B2(n310), .C1(n147), .C2(n637), .A(n639), .ZN(
        n3491) );
  AOI22_X1 U1007 ( .A1(n312), .A2(n640), .B1(n314), .B2(n641), .ZN(n639) );
  INV_X1 U1008 ( .A(\UUT/Mpath/the_mult/x_operand1[8] ), .ZN(n637) );
  OAI221_X1 U1009 ( .B1(n638), .B2(n316), .C1(\UUT/Mpath/the_alu/N67 ), .C2(
        net54889), .A(n642), .ZN(n3492) );
  AOI22_X1 U1010 ( .A1(n318), .A2(n640), .B1(n319), .B2(n641), .ZN(n642) );
  OAI22_X1 U1011 ( .A1(n5437), .A2(net54879), .B1(net54923), .B2(n638), .ZN(
        n3493) );
  OAI22_X1 U1012 ( .A1(n643), .A2(n546), .B1(n295), .B2(n2679), .ZN(n3494) );
  OAI221_X1 U1013 ( .B1(n644), .B2(n69), .C1(n90), .C2(n71), .A(n645), .ZN(
        n3495) );
  NAND2_X1 U1014 ( .A1(\UUT/Mpath/the_mult/x_operand2 [7]), .A2(n6409), .ZN(
        n645) );
  OAI222_X1 U1015 ( .A1(n90), .A2(n123), .B1(n644), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N70 ), .C2(net54893), .ZN(n3496) );
  INV_X1 U1016 ( .A(\UUT/break_code[7] ), .ZN(n644) );
  INV_X1 U1017 ( .A(n646), .ZN(n90) );
  OAI222_X1 U1018 ( .A1(n647), .A2(n129), .B1(n648), .B2(n131), .C1(n5439), 
        .C2(n132), .ZN(n646) );
  OAI221_X1 U1019 ( .B1(n133), .B2(n649), .C1(n5680), .C2(n135), .A(n650), 
        .ZN(n3497) );
  AOI22_X1 U1020 ( .A1(n137), .A2(n651), .B1(\UUT/Mpath/the_mult/Mad_out [39]), 
        .B2(n139), .ZN(n650) );
  OAI221_X1 U1021 ( .B1(n140), .B2(n652), .C1(n5618), .C2(n142), .A(n653), 
        .ZN(n3498) );
  AOI22_X1 U1022 ( .A1(n144), .A2(n651), .B1(\UUT/Mpath/the_mult/Mad_out [7]), 
        .B2(n145), .ZN(n653) );
  INV_X1 U1023 ( .A(n5619), .ZN(n651) );
  OAI22_X1 U1024 ( .A1(net54907), .A2(n654), .B1(n5619), .B2(net54871), .ZN(
        n3499) );
  OAI221_X1 U1025 ( .B1(n647), .B2(n310), .C1(n147), .C2(n654), .A(n655), .ZN(
        n3500) );
  AOI22_X1 U1026 ( .A1(n312), .A2(n656), .B1(n314), .B2(n657), .ZN(n655) );
  INV_X1 U1027 ( .A(\UUT/Mpath/the_mult/x_operand1[7] ), .ZN(n654) );
  OAI221_X1 U1028 ( .B1(n647), .B2(n316), .C1(\UUT/Mpath/the_alu/N69 ), .C2(
        net54887), .A(n658), .ZN(n3501) );
  AOI22_X1 U1029 ( .A1(n318), .A2(n656), .B1(n319), .B2(n657), .ZN(n658) );
  OAI22_X1 U1030 ( .A1(n5383), .A2(n6407), .B1(n648), .B2(n219), .ZN(n3502) );
  OAI22_X1 U1031 ( .A1(n5351), .A2(n6410), .B1(n648), .B2(n221), .ZN(n3503) );
  OAI22_X1 U1032 ( .A1(n5319), .A2(n6401), .B1(n648), .B2(n223), .ZN(n3504) );
  OAI22_X1 U1033 ( .A1(n5287), .A2(n6406), .B1(n648), .B2(n225), .ZN(n3505) );
  OAI22_X1 U1034 ( .A1(n5255), .A2(n6399), .B1(n648), .B2(n227), .ZN(n3506) );
  OAI22_X1 U1035 ( .A1(n5223), .A2(n6404), .B1(n648), .B2(n229), .ZN(n3507) );
  OAI22_X1 U1036 ( .A1(n5191), .A2(n6398), .B1(n648), .B2(n231), .ZN(n3508) );
  OAI22_X1 U1037 ( .A1(n5159), .A2(n6396), .B1(n648), .B2(n233), .ZN(n3509) );
  OAI22_X1 U1038 ( .A1(n5127), .A2(n6393), .B1(n648), .B2(n235), .ZN(n3510) );
  OAI22_X1 U1039 ( .A1(n5095), .A2(n6391), .B1(n648), .B2(n237), .ZN(n3511) );
  OAI22_X1 U1040 ( .A1(n5063), .A2(n6390), .B1(n648), .B2(n239), .ZN(n3512) );
  OAI22_X1 U1041 ( .A1(n5031), .A2(n6388), .B1(n648), .B2(n241), .ZN(n3513) );
  OAI22_X1 U1042 ( .A1(n4999), .A2(n6385), .B1(n648), .B2(n243), .ZN(n3514) );
  OAI22_X1 U1043 ( .A1(n4967), .A2(n6383), .B1(n648), .B2(n245), .ZN(n3515) );
  OAI22_X1 U1044 ( .A1(n4935), .A2(n6382), .B1(n648), .B2(n247), .ZN(n3516) );
  OAI22_X1 U1045 ( .A1(n4903), .A2(n6380), .B1(n648), .B2(n249), .ZN(n3517) );
  OAI22_X1 U1046 ( .A1(n4871), .A2(n6384), .B1(n648), .B2(n251), .ZN(n3518) );
  OAI22_X1 U1047 ( .A1(n4839), .A2(n6381), .B1(n648), .B2(n253), .ZN(n3519) );
  OAI22_X1 U1048 ( .A1(n4807), .A2(n6387), .B1(n648), .B2(n255), .ZN(n3520) );
  OAI22_X1 U1049 ( .A1(n4775), .A2(n6386), .B1(n648), .B2(n257), .ZN(n3521) );
  OAI22_X1 U1050 ( .A1(n4743), .A2(n6392), .B1(n648), .B2(n259), .ZN(n3522) );
  OAI22_X1 U1051 ( .A1(n4711), .A2(n6394), .B1(n648), .B2(n261), .ZN(n3523) );
  OAI22_X1 U1052 ( .A1(n4679), .A2(n6389), .B1(n648), .B2(n263), .ZN(n3524) );
  OAI22_X1 U1053 ( .A1(n4647), .A2(n6395), .B1(n648), .B2(n265), .ZN(n3525) );
  OAI22_X1 U1054 ( .A1(n4615), .A2(n6400), .B1(n648), .B2(n267), .ZN(n3526) );
  OAI22_X1 U1055 ( .A1(n4583), .A2(n6402), .B1(n648), .B2(n269), .ZN(n3527) );
  OAI22_X1 U1056 ( .A1(n4551), .A2(n6397), .B1(n648), .B2(n271), .ZN(n3528) );
  OAI22_X1 U1057 ( .A1(n4519), .A2(n6403), .B1(n648), .B2(n273), .ZN(n3529) );
  OAI22_X1 U1058 ( .A1(n4487), .A2(n6408), .B1(n648), .B2(n275), .ZN(n3530) );
  OAI22_X1 U1059 ( .A1(n4455), .A2(n6405), .B1(n648), .B2(n277), .ZN(n3531) );
  OAI22_X1 U1060 ( .A1(n4423), .A2(n6411), .B1(n648), .B2(n279), .ZN(n3532) );
  OAI222_X1 U1062 ( .A1(n5754), .A2(n489), .B1(n659), .B2(n660), .C1(n5710), 
        .C2(n5440), .ZN(n657) );
  AOI221_X1 U1063 ( .B1(n5757), .B2(n487), .C1(n5756), .C2(n5755), .A(n5759), 
        .ZN(n659) );
  INV_X1 U1064 ( .A(n5957), .ZN(n487) );
  OAI22_X1 U1065 ( .A1(n5440), .A2(net54881), .B1(net54923), .B2(n647), .ZN(
        n3533) );
  INV_X1 U1066 ( .A(n661), .ZN(n647) );
  OAI211_X1 U1067 ( .C1(n5618), .C2(n321), .A(n662), .B(n663), .ZN(n661) );
  AOI222_X1 U1068 ( .A1(n285), .A2(n664), .B1(\UUT/Mpath/out_jar[7] ), .B2(
        n325), .C1(n284), .C2(n665), .ZN(n663) );
  INV_X1 U1069 ( .A(n5680), .ZN(n665) );
  AOI22_X1 U1070 ( .A1(n6379), .A2(n6191), .B1(
        \UUT/Mpath/the_mult/x_mult_out[7] ), .B2(n291), .ZN(n662) );
  OAI22_X1 U1071 ( .A1(n666), .A2(n546), .B1(n295), .B2(n2682), .ZN(n3534) );
  OAI221_X1 U1072 ( .B1(n667), .B2(n69), .C1(n89), .C2(n71), .A(n668), .ZN(
        n3535) );
  NAND2_X1 U1073 ( .A1(\UUT/Mpath/the_mult/x_operand2 [6]), .A2(n6409), .ZN(
        n668) );
  OAI222_X1 U1074 ( .A1(n89), .A2(n123), .B1(n667), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N72 ), .C2(net54893), .ZN(n3536) );
  INV_X1 U1075 ( .A(\UUT/break_code[6] ), .ZN(n667) );
  INV_X1 U1076 ( .A(n669), .ZN(n89) );
  OAI222_X1 U1077 ( .A1(n670), .A2(n129), .B1(n671), .B2(n131), .C1(n5442), 
        .C2(n132), .ZN(n669) );
  OAI221_X1 U1078 ( .B1(n133), .B2(n672), .C1(n5681), .C2(n135), .A(n673), 
        .ZN(n3537) );
  AOI22_X1 U1079 ( .A1(n137), .A2(n674), .B1(\UUT/Mpath/the_mult/Mad_out [38]), 
        .B2(n139), .ZN(n673) );
  OAI221_X1 U1080 ( .B1(n140), .B2(n675), .C1(n5620), .C2(n142), .A(n676), 
        .ZN(n3538) );
  AOI22_X1 U1081 ( .A1(n144), .A2(n674), .B1(\UUT/Mpath/the_mult/Mad_out [6]), 
        .B2(n145), .ZN(n676) );
  INV_X1 U1082 ( .A(n5621), .ZN(n674) );
  OAI22_X1 U1083 ( .A1(net54907), .A2(n677), .B1(n5621), .B2(net54869), .ZN(
        n3539) );
  OAI221_X1 U1084 ( .B1(n670), .B2(n310), .C1(n147), .C2(n677), .A(n678), .ZN(
        n3540) );
  AOI22_X1 U1085 ( .A1(n312), .A2(n679), .B1(n314), .B2(n680), .ZN(n678) );
  INV_X1 U1086 ( .A(\UUT/Mpath/the_mult/x_operand1[6] ), .ZN(n677) );
  OAI221_X1 U1087 ( .B1(n670), .B2(n316), .C1(\UUT/Mpath/the_alu/N71 ), .C2(
        net54889), .A(n681), .ZN(n3541) );
  AOI22_X1 U1088 ( .A1(n318), .A2(n679), .B1(n319), .B2(n680), .ZN(n681) );
  OAI22_X1 U1089 ( .A1(n5384), .A2(n6407), .B1(n671), .B2(n219), .ZN(n3542) );
  OAI22_X1 U1090 ( .A1(n5352), .A2(n6410), .B1(n671), .B2(n221), .ZN(n3543) );
  OAI22_X1 U1091 ( .A1(n5320), .A2(n6401), .B1(n671), .B2(n223), .ZN(n3544) );
  OAI22_X1 U1092 ( .A1(n5288), .A2(n6406), .B1(n671), .B2(n225), .ZN(n3545) );
  OAI22_X1 U1093 ( .A1(n5256), .A2(n6399), .B1(n671), .B2(n227), .ZN(n3546) );
  OAI22_X1 U1094 ( .A1(n5224), .A2(n6404), .B1(n671), .B2(n229), .ZN(n3547) );
  OAI22_X1 U1095 ( .A1(n5192), .A2(n6398), .B1(n671), .B2(n231), .ZN(n3548) );
  OAI22_X1 U1096 ( .A1(n5160), .A2(n6396), .B1(n671), .B2(n233), .ZN(n3549) );
  OAI22_X1 U1097 ( .A1(n5128), .A2(n6393), .B1(n671), .B2(n235), .ZN(n3550) );
  OAI22_X1 U1098 ( .A1(n5096), .A2(n6391), .B1(n671), .B2(n237), .ZN(n3551) );
  OAI22_X1 U1099 ( .A1(n5064), .A2(n6390), .B1(n671), .B2(n239), .ZN(n3552) );
  OAI22_X1 U1100 ( .A1(n5032), .A2(n6388), .B1(n671), .B2(n241), .ZN(n3553) );
  OAI22_X1 U1101 ( .A1(n5000), .A2(n6385), .B1(n671), .B2(n243), .ZN(n3554) );
  OAI22_X1 U1102 ( .A1(n4968), .A2(n6383), .B1(n671), .B2(n245), .ZN(n3555) );
  OAI22_X1 U1103 ( .A1(n4936), .A2(n6382), .B1(n671), .B2(n247), .ZN(n3556) );
  OAI22_X1 U1104 ( .A1(n4904), .A2(n6380), .B1(n671), .B2(n249), .ZN(n3557) );
  OAI22_X1 U1105 ( .A1(n4872), .A2(n6384), .B1(n671), .B2(n251), .ZN(n3558) );
  OAI22_X1 U1106 ( .A1(n4840), .A2(n6381), .B1(n671), .B2(n253), .ZN(n3559) );
  OAI22_X1 U1107 ( .A1(n4808), .A2(n6387), .B1(n671), .B2(n255), .ZN(n3560) );
  OAI22_X1 U1108 ( .A1(n4776), .A2(n6386), .B1(n671), .B2(n257), .ZN(n3561) );
  OAI22_X1 U1109 ( .A1(n4744), .A2(n6392), .B1(n671), .B2(n259), .ZN(n3562) );
  OAI22_X1 U1110 ( .A1(n4712), .A2(n6394), .B1(n671), .B2(n261), .ZN(n3563) );
  OAI22_X1 U1111 ( .A1(n4680), .A2(n6389), .B1(n671), .B2(n263), .ZN(n3564) );
  OAI22_X1 U1112 ( .A1(n4648), .A2(n6395), .B1(n671), .B2(n265), .ZN(n3565) );
  OAI22_X1 U1113 ( .A1(n4616), .A2(n6400), .B1(n671), .B2(n267), .ZN(n3566) );
  OAI22_X1 U1114 ( .A1(n4584), .A2(n6402), .B1(n671), .B2(n269), .ZN(n3567) );
  OAI22_X1 U1115 ( .A1(n4552), .A2(n6397), .B1(n671), .B2(n271), .ZN(n3568) );
  OAI22_X1 U1116 ( .A1(n4520), .A2(n6403), .B1(n671), .B2(n273), .ZN(n3569) );
  OAI22_X1 U1117 ( .A1(n4488), .A2(n6408), .B1(n671), .B2(n275), .ZN(n3570) );
  OAI22_X1 U1118 ( .A1(n4456), .A2(n6405), .B1(n671), .B2(n277), .ZN(n3571) );
  OAI22_X1 U1119 ( .A1(n4424), .A2(n6411), .B1(n671), .B2(n279), .ZN(n3572) );
  OAI211_X1 U1121 ( .C1(n5710), .C2(n5443), .A(n682), .B(n683), .ZN(n680) );
  AOI222_X1 U1122 ( .A1(n5769), .A2(n684), .B1(n685), .B2(n513), .C1(n5774), 
        .C2(n686), .ZN(n683) );
  INV_X1 U1123 ( .A(n5776), .ZN(n513) );
  AOI22_X1 U1124 ( .A1(n5775), .A2(n687), .B1(n5771), .B2(n688), .ZN(n682) );
  OAI22_X1 U1125 ( .A1(n5443), .A2(net54881), .B1(net54923), .B2(n670), .ZN(
        n3573) );
  INV_X1 U1126 ( .A(n689), .ZN(n670) );
  OAI211_X1 U1127 ( .C1(n5620), .C2(n321), .A(n690), .B(n691), .ZN(n689) );
  AOI222_X1 U1128 ( .A1(n285), .A2(n692), .B1(\UUT/Mpath/out_jar[6] ), .B2(
        n325), .C1(n284), .C2(n693), .ZN(n691) );
  INV_X1 U1129 ( .A(n5681), .ZN(n693) );
  AOI22_X1 U1130 ( .A1(n6379), .A2(n6192), .B1(
        \UUT/Mpath/the_mult/x_mult_out[6] ), .B2(n291), .ZN(n690) );
  OAI22_X1 U1131 ( .A1(n694), .A2(n546), .B1(n295), .B2(n2685), .ZN(n3574) );
  OAI221_X1 U1132 ( .B1(n695), .B2(n69), .C1(n88), .C2(n71), .A(n696), .ZN(
        n3575) );
  NAND2_X1 U1133 ( .A1(\UUT/Mpath/the_mult/x_operand2 [5]), .A2(n6409), .ZN(
        n696) );
  OAI222_X1 U1134 ( .A1(n88), .A2(n123), .B1(n695), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N74 ), .C2(net54893), .ZN(n3576) );
  INV_X1 U1135 ( .A(\UUT/break_code[5] ), .ZN(n695) );
  INV_X1 U1136 ( .A(n697), .ZN(n88) );
  OAI222_X1 U1137 ( .A1(n698), .A2(n129), .B1(n699), .B2(n131), .C1(n5445), 
        .C2(n132), .ZN(n697) );
  OAI221_X1 U1138 ( .B1(n133), .B2(n700), .C1(n5682), .C2(n135), .A(n701), 
        .ZN(n3577) );
  AOI22_X1 U1139 ( .A1(n137), .A2(n702), .B1(\UUT/Mpath/the_mult/Mad_out [37]), 
        .B2(n139), .ZN(n701) );
  OAI221_X1 U1140 ( .B1(n140), .B2(n703), .C1(n5622), .C2(n142), .A(n704), 
        .ZN(n3578) );
  AOI22_X1 U1141 ( .A1(n144), .A2(n702), .B1(\UUT/Mpath/the_mult/Mad_out [5]), 
        .B2(n145), .ZN(n704) );
  INV_X1 U1142 ( .A(n5623), .ZN(n702) );
  OAI22_X1 U1143 ( .A1(net54909), .A2(n705), .B1(n5623), .B2(net54869), .ZN(
        n3579) );
  OAI221_X1 U1144 ( .B1(n698), .B2(n310), .C1(n147), .C2(n705), .A(n706), .ZN(
        n3580) );
  AOI22_X1 U1145 ( .A1(n312), .A2(n707), .B1(n314), .B2(n708), .ZN(n706) );
  INV_X1 U1146 ( .A(\UUT/Mpath/the_mult/x_operand1[5] ), .ZN(n705) );
  OAI221_X1 U1147 ( .B1(n698), .B2(n316), .C1(\UUT/Mpath/the_alu/N73 ), .C2(
        net54887), .A(n709), .ZN(n3581) );
  AOI22_X1 U1148 ( .A1(n318), .A2(n707), .B1(n319), .B2(n708), .ZN(n709) );
  OAI22_X1 U1149 ( .A1(n5385), .A2(n6407), .B1(n699), .B2(n219), .ZN(n3582) );
  OAI22_X1 U1150 ( .A1(n5353), .A2(n6410), .B1(n699), .B2(n221), .ZN(n3583) );
  OAI22_X1 U1151 ( .A1(n5321), .A2(n6401), .B1(n699), .B2(n223), .ZN(n3584) );
  OAI22_X1 U1152 ( .A1(n5289), .A2(n6406), .B1(n699), .B2(n225), .ZN(n3585) );
  OAI22_X1 U1153 ( .A1(n5257), .A2(n6399), .B1(n699), .B2(n227), .ZN(n3586) );
  OAI22_X1 U1154 ( .A1(n5225), .A2(n6404), .B1(n699), .B2(n229), .ZN(n3587) );
  OAI22_X1 U1155 ( .A1(n5193), .A2(n6398), .B1(n699), .B2(n231), .ZN(n3588) );
  OAI22_X1 U1156 ( .A1(n5161), .A2(n6396), .B1(n699), .B2(n233), .ZN(n3589) );
  OAI22_X1 U1157 ( .A1(n5129), .A2(n6393), .B1(n699), .B2(n235), .ZN(n3590) );
  OAI22_X1 U1158 ( .A1(n5097), .A2(n6391), .B1(n699), .B2(n237), .ZN(n3591) );
  OAI22_X1 U1159 ( .A1(n5065), .A2(n6390), .B1(n699), .B2(n239), .ZN(n3592) );
  OAI22_X1 U1160 ( .A1(n5033), .A2(n6388), .B1(n699), .B2(n241), .ZN(n3593) );
  OAI22_X1 U1161 ( .A1(n5001), .A2(n6385), .B1(n699), .B2(n243), .ZN(n3594) );
  OAI22_X1 U1162 ( .A1(n4969), .A2(n6383), .B1(n699), .B2(n245), .ZN(n3595) );
  OAI22_X1 U1163 ( .A1(n4937), .A2(n6382), .B1(n699), .B2(n247), .ZN(n3596) );
  OAI22_X1 U1164 ( .A1(n4905), .A2(n6380), .B1(n699), .B2(n249), .ZN(n3597) );
  OAI22_X1 U1165 ( .A1(n4873), .A2(n6384), .B1(n699), .B2(n251), .ZN(n3598) );
  OAI22_X1 U1166 ( .A1(n4841), .A2(n6381), .B1(n699), .B2(n253), .ZN(n3599) );
  OAI22_X1 U1167 ( .A1(n4809), .A2(n6387), .B1(n699), .B2(n255), .ZN(n3600) );
  OAI22_X1 U1168 ( .A1(n4777), .A2(n6386), .B1(n699), .B2(n257), .ZN(n3601) );
  OAI22_X1 U1169 ( .A1(n4745), .A2(n6392), .B1(n699), .B2(n259), .ZN(n3602) );
  OAI22_X1 U1170 ( .A1(n4713), .A2(n6394), .B1(n699), .B2(n261), .ZN(n3603) );
  OAI22_X1 U1171 ( .A1(n4681), .A2(n6389), .B1(n699), .B2(n263), .ZN(n3604) );
  OAI22_X1 U1172 ( .A1(n4649), .A2(n6395), .B1(n699), .B2(n265), .ZN(n3605) );
  OAI22_X1 U1173 ( .A1(n4617), .A2(n6400), .B1(n699), .B2(n267), .ZN(n3606) );
  OAI22_X1 U1174 ( .A1(n4585), .A2(n6402), .B1(n699), .B2(n269), .ZN(n3607) );
  OAI22_X1 U1175 ( .A1(n4553), .A2(n6397), .B1(n699), .B2(n271), .ZN(n3608) );
  OAI22_X1 U1176 ( .A1(n4521), .A2(n6403), .B1(n699), .B2(n273), .ZN(n3609) );
  OAI22_X1 U1177 ( .A1(n4489), .A2(n6408), .B1(n699), .B2(n275), .ZN(n3610) );
  OAI22_X1 U1178 ( .A1(n4457), .A2(n6405), .B1(n699), .B2(n277), .ZN(n3611) );
  OAI22_X1 U1179 ( .A1(n4425), .A2(n6411), .B1(n699), .B2(n279), .ZN(n3612) );
  OAI211_X1 U1181 ( .C1(n5710), .C2(n5446), .A(n710), .B(n711), .ZN(n708) );
  AOI222_X1 U1182 ( .A1(n5786), .A2(n684), .B1(n685), .B2(n538), .C1(n5791), 
        .C2(n686), .ZN(n711) );
  INV_X1 U1183 ( .A(n5793), .ZN(n538) );
  AOI22_X1 U1184 ( .A1(n5792), .A2(n687), .B1(n5788), .B2(n688), .ZN(n710) );
  OAI22_X1 U1185 ( .A1(n5446), .A2(net54883), .B1(net54923), .B2(n698), .ZN(
        n3613) );
  INV_X1 U1186 ( .A(n712), .ZN(n698) );
  OAI211_X1 U1187 ( .C1(n5622), .C2(n321), .A(n713), .B(n714), .ZN(n712) );
  AOI222_X1 U1188 ( .A1(n285), .A2(n715), .B1(\UUT/Mpath/out_jar[5] ), .B2(
        n325), .C1(n284), .C2(n716), .ZN(n714) );
  INV_X1 U1189 ( .A(n5682), .ZN(n716) );
  AOI22_X1 U1190 ( .A1(n6379), .A2(n6193), .B1(
        \UUT/Mpath/the_mult/x_mult_out[5] ), .B2(n291), .ZN(n713) );
  OAI22_X1 U1191 ( .A1(n6463), .A2(n546), .B1(n295), .B2(n2688), .ZN(n3614) );
  OAI221_X1 U1192 ( .B1(n718), .B2(n69), .C1(n87), .C2(n71), .A(n719), .ZN(
        n3615) );
  NAND2_X1 U1193 ( .A1(\UUT/Mpath/the_mult/x_operand2 [4]), .A2(n6409), .ZN(
        n719) );
  OAI222_X1 U1194 ( .A1(n87), .A2(n123), .B1(n718), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N76 ), .C2(net54891), .ZN(n3616) );
  INV_X1 U1195 ( .A(n720), .ZN(n87) );
  OAI222_X1 U1196 ( .A1(n721), .A2(n129), .B1(n722), .B2(n131), .C1(n5448), 
        .C2(n132), .ZN(n720) );
  OAI221_X1 U1197 ( .B1(n133), .B2(n723), .C1(n5683), .C2(n135), .A(n724), 
        .ZN(n3617) );
  AOI22_X1 U1198 ( .A1(n137), .A2(n725), .B1(\UUT/Mpath/the_mult/Mad_out [36]), 
        .B2(n139), .ZN(n724) );
  OAI221_X1 U1199 ( .B1(n140), .B2(n726), .C1(n5624), .C2(n142), .A(n727), 
        .ZN(n3618) );
  AOI22_X1 U1200 ( .A1(n144), .A2(n725), .B1(\UUT/Mpath/the_mult/Mad_out [4]), 
        .B2(n145), .ZN(n727) );
  INV_X1 U1201 ( .A(n5625), .ZN(n725) );
  OAI22_X1 U1202 ( .A1(net54907), .A2(n728), .B1(n5625), .B2(net54869), .ZN(
        n3619) );
  OAI221_X1 U1203 ( .B1(n721), .B2(n310), .C1(n147), .C2(n728), .A(n729), .ZN(
        n3620) );
  AOI22_X1 U1204 ( .A1(n312), .A2(n730), .B1(n314), .B2(n731), .ZN(n729) );
  INV_X1 U1205 ( .A(\UUT/Mpath/the_mult/x_operand1[4] ), .ZN(n728) );
  OAI221_X1 U1206 ( .B1(n721), .B2(n316), .C1(\UUT/Mpath/the_alu/N75 ), .C2(
        net54887), .A(n732), .ZN(n3621) );
  AOI22_X1 U1207 ( .A1(n318), .A2(n730), .B1(n319), .B2(n731), .ZN(n732) );
  OAI22_X1 U1208 ( .A1(n5386), .A2(n6407), .B1(n722), .B2(n219), .ZN(n3622) );
  OAI22_X1 U1209 ( .A1(n5354), .A2(n6410), .B1(n722), .B2(n221), .ZN(n3623) );
  OAI22_X1 U1210 ( .A1(n5322), .A2(n6401), .B1(n722), .B2(n223), .ZN(n3624) );
  OAI22_X1 U1211 ( .A1(n5290), .A2(n6406), .B1(n722), .B2(n225), .ZN(n3625) );
  OAI22_X1 U1212 ( .A1(n5258), .A2(n6399), .B1(n722), .B2(n227), .ZN(n3626) );
  OAI22_X1 U1213 ( .A1(n5226), .A2(n6404), .B1(n722), .B2(n229), .ZN(n3627) );
  OAI22_X1 U1214 ( .A1(n5194), .A2(n6398), .B1(n722), .B2(n231), .ZN(n3628) );
  OAI22_X1 U1215 ( .A1(n5162), .A2(n6396), .B1(n722), .B2(n233), .ZN(n3629) );
  OAI22_X1 U1216 ( .A1(n5130), .A2(n6393), .B1(n722), .B2(n235), .ZN(n3630) );
  OAI22_X1 U1217 ( .A1(n5098), .A2(n6391), .B1(n722), .B2(n237), .ZN(n3631) );
  OAI22_X1 U1218 ( .A1(n5066), .A2(n6390), .B1(n722), .B2(n239), .ZN(n3632) );
  OAI22_X1 U1219 ( .A1(n5034), .A2(n6388), .B1(n722), .B2(n241), .ZN(n3633) );
  OAI22_X1 U1220 ( .A1(n5002), .A2(n6385), .B1(n722), .B2(n243), .ZN(n3634) );
  OAI22_X1 U1221 ( .A1(n4970), .A2(n6383), .B1(n722), .B2(n245), .ZN(n3635) );
  OAI22_X1 U1222 ( .A1(n4938), .A2(n6382), .B1(n722), .B2(n247), .ZN(n3636) );
  OAI22_X1 U1223 ( .A1(n4906), .A2(n6380), .B1(n722), .B2(n249), .ZN(n3637) );
  OAI22_X1 U1224 ( .A1(n4874), .A2(n6384), .B1(n722), .B2(n251), .ZN(n3638) );
  OAI22_X1 U1225 ( .A1(n4842), .A2(n6381), .B1(n722), .B2(n253), .ZN(n3639) );
  OAI22_X1 U1226 ( .A1(n4810), .A2(n6387), .B1(n722), .B2(n255), .ZN(n3640) );
  OAI22_X1 U1227 ( .A1(n4778), .A2(n6386), .B1(n722), .B2(n257), .ZN(n3641) );
  OAI22_X1 U1228 ( .A1(n4746), .A2(n6392), .B1(n722), .B2(n259), .ZN(n3642) );
  OAI22_X1 U1229 ( .A1(n4714), .A2(n6394), .B1(n722), .B2(n261), .ZN(n3643) );
  OAI22_X1 U1230 ( .A1(n4682), .A2(n6389), .B1(n722), .B2(n263), .ZN(n3644) );
  OAI22_X1 U1231 ( .A1(n4650), .A2(n6395), .B1(n722), .B2(n265), .ZN(n3645) );
  OAI22_X1 U1232 ( .A1(n4618), .A2(n6400), .B1(n722), .B2(n267), .ZN(n3646) );
  OAI22_X1 U1233 ( .A1(n4586), .A2(n6402), .B1(n722), .B2(n269), .ZN(n3647) );
  OAI22_X1 U1234 ( .A1(n4554), .A2(n6397), .B1(n722), .B2(n271), .ZN(n3648) );
  OAI22_X1 U1235 ( .A1(n4522), .A2(n6403), .B1(n722), .B2(n273), .ZN(n3649) );
  OAI22_X1 U1236 ( .A1(n4490), .A2(n6408), .B1(n722), .B2(n275), .ZN(n3650) );
  OAI22_X1 U1237 ( .A1(n4458), .A2(n6405), .B1(n722), .B2(n277), .ZN(n3651) );
  OAI22_X1 U1238 ( .A1(n4426), .A2(n6411), .B1(n722), .B2(n279), .ZN(n3652) );
  OAI211_X1 U1240 ( .C1(n5710), .C2(n5449), .A(n733), .B(n734), .ZN(n731) );
  AOI222_X1 U1241 ( .A1(n5799), .A2(n684), .B1(n685), .B2(n564), .C1(n5804), 
        .C2(n686), .ZN(n734) );
  INV_X1 U1242 ( .A(n5806), .ZN(n564) );
  AOI22_X1 U1243 ( .A1(n5805), .A2(n687), .B1(n5801), .B2(n688), .ZN(n733) );
  OAI22_X1 U1244 ( .A1(n5449), .A2(net54881), .B1(net54923), .B2(n721), .ZN(
        n3653) );
  INV_X1 U1245 ( .A(n735), .ZN(n721) );
  OAI211_X1 U1246 ( .C1(n5624), .C2(n321), .A(n736), .B(n737), .ZN(n735) );
  AOI222_X1 U1247 ( .A1(n285), .A2(n738), .B1(\UUT/Mpath/out_jar[4] ), .B2(
        n325), .C1(n284), .C2(n739), .ZN(n737) );
  INV_X1 U1248 ( .A(n5683), .ZN(n739) );
  AOI22_X1 U1249 ( .A1(n6379), .A2(n6194), .B1(
        \UUT/Mpath/the_mult/x_mult_out[4] ), .B2(n291), .ZN(n736) );
  OAI22_X1 U1250 ( .A1(n740), .A2(n546), .B1(n295), .B2(n2691), .ZN(n3654) );
  OAI221_X1 U1251 ( .B1(n741), .B2(n69), .C1(n86), .C2(n71), .A(n742), .ZN(
        n3655) );
  NAND2_X1 U1252 ( .A1(\UUT/Mpath/the_mult/x_operand2 [3]), .A2(n6409), .ZN(
        n742) );
  OAI222_X1 U1253 ( .A1(n86), .A2(n123), .B1(n741), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N78 ), .C2(net54891), .ZN(n3656) );
  INV_X1 U1254 ( .A(n743), .ZN(n86) );
  OAI222_X1 U1255 ( .A1(n744), .A2(n129), .B1(n745), .B2(n131), .C1(n5451), 
        .C2(n132), .ZN(n743) );
  OAI221_X1 U1256 ( .B1(n133), .B2(n746), .C1(n5684), .C2(n135), .A(n747), 
        .ZN(n3657) );
  AOI22_X1 U1257 ( .A1(n137), .A2(n748), .B1(\UUT/Mpath/the_mult/Mad_out [35]), 
        .B2(n139), .ZN(n747) );
  OAI221_X1 U1258 ( .B1(n140), .B2(n749), .C1(n5626), .C2(n142), .A(n750), 
        .ZN(n3658) );
  AOI22_X1 U1259 ( .A1(n144), .A2(n748), .B1(\UUT/Mpath/the_mult/Mad_out [3]), 
        .B2(n145), .ZN(n750) );
  INV_X1 U1260 ( .A(n5627), .ZN(n748) );
  OAI22_X1 U1261 ( .A1(net54907), .A2(n751), .B1(n5627), .B2(net54871), .ZN(
        n3659) );
  OAI221_X1 U1262 ( .B1(n744), .B2(n310), .C1(n147), .C2(n751), .A(n752), .ZN(
        n3660) );
  AOI22_X1 U1263 ( .A1(n312), .A2(n753), .B1(n314), .B2(n754), .ZN(n752) );
  INV_X1 U1264 ( .A(\UUT/Mpath/the_mult/x_operand1[3] ), .ZN(n751) );
  OAI221_X1 U1265 ( .B1(n744), .B2(n316), .C1(\UUT/Mpath/the_alu/N77 ), .C2(
        net54887), .A(n755), .ZN(n3661) );
  AOI22_X1 U1266 ( .A1(n318), .A2(n753), .B1(n319), .B2(n754), .ZN(n755) );
  OAI22_X1 U1267 ( .A1(n5387), .A2(n6407), .B1(n745), .B2(n219), .ZN(n3662) );
  OAI22_X1 U1268 ( .A1(n5355), .A2(n6410), .B1(n745), .B2(n221), .ZN(n3663) );
  OAI22_X1 U1269 ( .A1(n5323), .A2(n6401), .B1(n745), .B2(n223), .ZN(n3664) );
  OAI22_X1 U1270 ( .A1(n5291), .A2(n6406), .B1(n745), .B2(n225), .ZN(n3665) );
  OAI22_X1 U1271 ( .A1(n5259), .A2(n6399), .B1(n745), .B2(n227), .ZN(n3666) );
  OAI22_X1 U1272 ( .A1(n5227), .A2(n6404), .B1(n745), .B2(n229), .ZN(n3667) );
  OAI22_X1 U1273 ( .A1(n5195), .A2(n6398), .B1(n745), .B2(n231), .ZN(n3668) );
  OAI22_X1 U1274 ( .A1(n5163), .A2(n6396), .B1(n745), .B2(n233), .ZN(n3669) );
  OAI22_X1 U1275 ( .A1(n5131), .A2(n6393), .B1(n745), .B2(n235), .ZN(n3670) );
  OAI22_X1 U1276 ( .A1(n5099), .A2(n6391), .B1(n745), .B2(n237), .ZN(n3671) );
  OAI22_X1 U1277 ( .A1(n5067), .A2(n6390), .B1(n745), .B2(n239), .ZN(n3672) );
  OAI22_X1 U1278 ( .A1(n5035), .A2(n6388), .B1(n745), .B2(n241), .ZN(n3673) );
  OAI22_X1 U1279 ( .A1(n5003), .A2(n6385), .B1(n745), .B2(n243), .ZN(n3674) );
  OAI22_X1 U1280 ( .A1(n4971), .A2(n6383), .B1(n745), .B2(n245), .ZN(n3675) );
  OAI22_X1 U1281 ( .A1(n4939), .A2(n6382), .B1(n745), .B2(n247), .ZN(n3676) );
  OAI22_X1 U1282 ( .A1(n4907), .A2(n6380), .B1(n745), .B2(n249), .ZN(n3677) );
  OAI22_X1 U1283 ( .A1(n4875), .A2(n6384), .B1(n745), .B2(n251), .ZN(n3678) );
  OAI22_X1 U1284 ( .A1(n4843), .A2(n6381), .B1(n745), .B2(n253), .ZN(n3679) );
  OAI22_X1 U1285 ( .A1(n4811), .A2(n6387), .B1(n745), .B2(n255), .ZN(n3680) );
  OAI22_X1 U1286 ( .A1(n4779), .A2(n6386), .B1(n745), .B2(n257), .ZN(n3681) );
  OAI22_X1 U1287 ( .A1(n4747), .A2(n6392), .B1(n745), .B2(n259), .ZN(n3682) );
  OAI22_X1 U1288 ( .A1(n4715), .A2(n6394), .B1(n745), .B2(n261), .ZN(n3683) );
  OAI22_X1 U1289 ( .A1(n4683), .A2(n6389), .B1(n745), .B2(n263), .ZN(n3684) );
  OAI22_X1 U1290 ( .A1(n4651), .A2(n6395), .B1(n745), .B2(n265), .ZN(n3685) );
  OAI22_X1 U1291 ( .A1(n4619), .A2(n6400), .B1(n745), .B2(n267), .ZN(n3686) );
  OAI22_X1 U1292 ( .A1(n4587), .A2(n6402), .B1(n745), .B2(n269), .ZN(n3687) );
  OAI22_X1 U1293 ( .A1(n4555), .A2(n6397), .B1(n745), .B2(n271), .ZN(n3688) );
  OAI22_X1 U1294 ( .A1(n4523), .A2(n6403), .B1(n745), .B2(n273), .ZN(n3689) );
  OAI22_X1 U1295 ( .A1(n4491), .A2(n6408), .B1(n745), .B2(n275), .ZN(n3690) );
  OAI22_X1 U1296 ( .A1(n4459), .A2(n6405), .B1(n745), .B2(n277), .ZN(n3691) );
  OAI22_X1 U1297 ( .A1(n4427), .A2(n6411), .B1(n745), .B2(n279), .ZN(n3692) );
  OAI211_X1 U1299 ( .C1(n5710), .C2(n5452), .A(n756), .B(n757), .ZN(n754) );
  AOI222_X1 U1300 ( .A1(n5812), .A2(n684), .B1(n685), .B2(n589), .C1(n5817), 
        .C2(n686), .ZN(n757) );
  INV_X1 U1301 ( .A(n5819), .ZN(n589) );
  AOI22_X1 U1302 ( .A1(n5818), .A2(n687), .B1(n5814), .B2(n688), .ZN(n756) );
  OAI22_X1 U1303 ( .A1(n5452), .A2(net54883), .B1(net54923), .B2(n744), .ZN(
        n3693) );
  INV_X1 U1304 ( .A(n758), .ZN(n744) );
  OAI211_X1 U1305 ( .C1(n5626), .C2(n321), .A(n759), .B(n760), .ZN(n758) );
  AOI222_X1 U1306 ( .A1(n285), .A2(n761), .B1(\UUT/Mpath/out_jar[3] ), .B2(
        n325), .C1(n284), .C2(n762), .ZN(n760) );
  INV_X1 U1307 ( .A(n5684), .ZN(n762) );
  AOI22_X1 U1308 ( .A1(n6379), .A2(n6195), .B1(
        \UUT/Mpath/the_mult/x_mult_out[3] ), .B2(n291), .ZN(n759) );
  OAI22_X1 U1309 ( .A1(n763), .A2(n546), .B1(n295), .B2(n2694), .ZN(n3694) );
  OAI221_X1 U1310 ( .B1(n764), .B2(n69), .C1(n85), .C2(n71), .A(n765), .ZN(
        n3695) );
  NAND2_X1 U1311 ( .A1(\UUT/Mpath/the_mult/x_operand2 [2]), .A2(n6409), .ZN(
        n765) );
  OAI222_X1 U1312 ( .A1(n85), .A2(n123), .B1(n764), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N80 ), .C2(net54891), .ZN(n3696) );
  INV_X1 U1313 ( .A(n766), .ZN(n85) );
  OAI222_X1 U1314 ( .A1(n767), .A2(n129), .B1(n768), .B2(n131), .C1(n5460), 
        .C2(n132), .ZN(n766) );
  OAI221_X1 U1315 ( .B1(n133), .B2(n769), .C1(n5687), .C2(n135), .A(n770), 
        .ZN(n3697) );
  AOI22_X1 U1316 ( .A1(n137), .A2(n771), .B1(\UUT/Mpath/the_mult/Mad_out [34]), 
        .B2(n139), .ZN(n770) );
  OAI221_X1 U1317 ( .B1(n140), .B2(n772), .C1(n5632), .C2(n142), .A(n773), 
        .ZN(n3698) );
  AOI22_X1 U1318 ( .A1(n144), .A2(n771), .B1(\UUT/Mpath/the_mult/Mad_out [2]), 
        .B2(n145), .ZN(n773) );
  INV_X1 U1319 ( .A(n5633), .ZN(n771) );
  OAI22_X1 U1320 ( .A1(net54907), .A2(n774), .B1(n5633), .B2(net54871), .ZN(
        n3699) );
  OAI221_X1 U1321 ( .B1(n767), .B2(n310), .C1(n147), .C2(n774), .A(n775), .ZN(
        n3700) );
  AOI22_X1 U1322 ( .A1(n312), .A2(n776), .B1(n314), .B2(n777), .ZN(n775) );
  INV_X1 U1323 ( .A(\UUT/Mpath/the_mult/x_operand1[2] ), .ZN(n774) );
  OAI221_X1 U1324 ( .B1(n767), .B2(n316), .C1(\UUT/Mpath/the_alu/N79 ), .C2(
        net54887), .A(n778), .ZN(n3701) );
  AOI22_X1 U1325 ( .A1(n318), .A2(n776), .B1(n319), .B2(n777), .ZN(n778) );
  OAI22_X1 U1326 ( .A1(n5390), .A2(n6407), .B1(n768), .B2(n219), .ZN(n3702) );
  OAI22_X1 U1327 ( .A1(n5358), .A2(n6410), .B1(n768), .B2(n221), .ZN(n3703) );
  OAI22_X1 U1328 ( .A1(n5326), .A2(n6401), .B1(n768), .B2(n223), .ZN(n3704) );
  OAI22_X1 U1329 ( .A1(n5294), .A2(n6406), .B1(n768), .B2(n225), .ZN(n3705) );
  OAI22_X1 U1330 ( .A1(n5262), .A2(n6399), .B1(n768), .B2(n227), .ZN(n3706) );
  OAI22_X1 U1331 ( .A1(n5230), .A2(n6404), .B1(n768), .B2(n229), .ZN(n3707) );
  OAI22_X1 U1332 ( .A1(n5198), .A2(n6398), .B1(n768), .B2(n231), .ZN(n3708) );
  OAI22_X1 U1333 ( .A1(n5166), .A2(n6396), .B1(n768), .B2(n233), .ZN(n3709) );
  OAI22_X1 U1334 ( .A1(n5134), .A2(n6393), .B1(n768), .B2(n235), .ZN(n3710) );
  OAI22_X1 U1335 ( .A1(n5102), .A2(n6391), .B1(n768), .B2(n237), .ZN(n3711) );
  OAI22_X1 U1336 ( .A1(n5070), .A2(n6390), .B1(n768), .B2(n239), .ZN(n3712) );
  OAI22_X1 U1337 ( .A1(n5038), .A2(n6388), .B1(n768), .B2(n241), .ZN(n3713) );
  OAI22_X1 U1338 ( .A1(n5006), .A2(n6385), .B1(n768), .B2(n243), .ZN(n3714) );
  OAI22_X1 U1339 ( .A1(n4974), .A2(n6383), .B1(n768), .B2(n245), .ZN(n3715) );
  OAI22_X1 U1340 ( .A1(n4942), .A2(n6382), .B1(n768), .B2(n247), .ZN(n3716) );
  OAI22_X1 U1341 ( .A1(n4910), .A2(n6380), .B1(n768), .B2(n249), .ZN(n3717) );
  OAI22_X1 U1342 ( .A1(n4878), .A2(n6384), .B1(n768), .B2(n251), .ZN(n3718) );
  OAI22_X1 U1343 ( .A1(n4846), .A2(n6381), .B1(n768), .B2(n253), .ZN(n3719) );
  OAI22_X1 U1344 ( .A1(n4814), .A2(n6387), .B1(n768), .B2(n255), .ZN(n3720) );
  OAI22_X1 U1345 ( .A1(n4782), .A2(n6386), .B1(n768), .B2(n257), .ZN(n3721) );
  OAI22_X1 U1346 ( .A1(n4750), .A2(n6392), .B1(n768), .B2(n259), .ZN(n3722) );
  OAI22_X1 U1347 ( .A1(n4718), .A2(n6394), .B1(n768), .B2(n261), .ZN(n3723) );
  OAI22_X1 U1348 ( .A1(n4686), .A2(n6389), .B1(n768), .B2(n263), .ZN(n3724) );
  OAI22_X1 U1349 ( .A1(n4654), .A2(n6395), .B1(n768), .B2(n265), .ZN(n3725) );
  OAI22_X1 U1350 ( .A1(n4622), .A2(n6400), .B1(n768), .B2(n267), .ZN(n3726) );
  OAI22_X1 U1351 ( .A1(n4590), .A2(n6402), .B1(n768), .B2(n269), .ZN(n3727) );
  OAI22_X1 U1352 ( .A1(n4558), .A2(n6397), .B1(n768), .B2(n271), .ZN(n3728) );
  OAI22_X1 U1353 ( .A1(n4526), .A2(n6403), .B1(n768), .B2(n273), .ZN(n3729) );
  OAI22_X1 U1354 ( .A1(n4494), .A2(n6408), .B1(n768), .B2(n275), .ZN(n3730) );
  OAI22_X1 U1355 ( .A1(n4462), .A2(n6405), .B1(n768), .B2(n277), .ZN(n3731) );
  OAI22_X1 U1356 ( .A1(n4430), .A2(n6411), .B1(n768), .B2(n279), .ZN(n3732) );
  OAI211_X1 U1358 ( .C1(n5710), .C2(n5461), .A(n779), .B(n780), .ZN(n777) );
  AOI222_X1 U1359 ( .A1(n5838), .A2(n684), .B1(n685), .B2(n781), .C1(n5843), 
        .C2(n686), .ZN(n780) );
  AOI22_X1 U1360 ( .A1(n5844), .A2(n687), .B1(n5840), .B2(n688), .ZN(n779) );
  OAI22_X1 U1361 ( .A1(n5461), .A2(net54885), .B1(net54923), .B2(n767), .ZN(
        n3733) );
  INV_X1 U1362 ( .A(n782), .ZN(n767) );
  OAI211_X1 U1363 ( .C1(n5632), .C2(n321), .A(n783), .B(n784), .ZN(n782) );
  AOI222_X1 U1364 ( .A1(n285), .A2(n785), .B1(\UUT/Mpath/out_jar[2] ), .B2(
        n325), .C1(n284), .C2(n786), .ZN(n784) );
  INV_X1 U1365 ( .A(n5687), .ZN(n786) );
  AOI22_X1 U1366 ( .A1(n6379), .A2(n6202), .B1(
        \UUT/Mpath/the_mult/x_mult_out[2] ), .B2(n291), .ZN(n783) );
  OAI221_X1 U1367 ( .B1(n787), .B2(n69), .C1(n84), .C2(n71), .A(n788), .ZN(
        n3734) );
  NAND2_X1 U1368 ( .A1(\UUT/Mpath/the_mult/x_operand2 [1]), .A2(n6409), .ZN(
        n788) );
  NAND2_X1 U1370 ( .A1(n147), .A2(n789), .ZN(n69) );
  OAI221_X1 U1373 ( .B1(n133), .B2(n791), .C1(n5698), .C2(n135), .A(n792), 
        .ZN(n3736) );
  AOI22_X1 U1374 ( .A1(n137), .A2(n793), .B1(\UUT/Mpath/the_mult/Mad_out [33]), 
        .B2(n139), .ZN(n792) );
  OAI221_X1 U1375 ( .B1(n140), .B2(n794), .C1(n5654), .C2(n142), .A(n795), 
        .ZN(n3737) );
  AOI22_X1 U1376 ( .A1(n144), .A2(n793), .B1(\UUT/Mpath/the_mult/Mad_out [1]), 
        .B2(n145), .ZN(n795) );
  INV_X1 U1377 ( .A(n5655), .ZN(n793) );
  OAI22_X1 U1378 ( .A1(net54907), .A2(n796), .B1(n5655), .B2(net54871), .ZN(
        n3738) );
  OAI221_X1 U1379 ( .B1(n797), .B2(n310), .C1(n147), .C2(n796), .A(n798), .ZN(
        n3739) );
  AOI22_X1 U1380 ( .A1(n312), .A2(n799), .B1(n314), .B2(n800), .ZN(n798) );
  INV_X1 U1381 ( .A(\UUT/Mpath/the_mult/x_operand1[1] ), .ZN(n796) );
  OAI221_X1 U1382 ( .B1(n797), .B2(n316), .C1(\UUT/Mpath/the_alu/N81 ), .C2(
        net54885), .A(n801), .ZN(n3740) );
  AOI22_X1 U1383 ( .A1(n318), .A2(n799), .B1(n319), .B2(n800), .ZN(n801) );
  OAI22_X1 U1384 ( .A1(n5401), .A2(n6407), .B1(n802), .B2(n219), .ZN(n3741) );
  OAI22_X1 U1385 ( .A1(n5369), .A2(n6410), .B1(n802), .B2(n221), .ZN(n3742) );
  OAI22_X1 U1386 ( .A1(n5337), .A2(n6401), .B1(n802), .B2(n223), .ZN(n3743) );
  OAI22_X1 U1387 ( .A1(n5305), .A2(n6406), .B1(n802), .B2(n225), .ZN(n3744) );
  OAI22_X1 U1388 ( .A1(n5273), .A2(n6399), .B1(n802), .B2(n227), .ZN(n3745) );
  OAI22_X1 U1389 ( .A1(n5241), .A2(n6404), .B1(n802), .B2(n229), .ZN(n3746) );
  OAI22_X1 U1390 ( .A1(n5209), .A2(n6398), .B1(n802), .B2(n231), .ZN(n3747) );
  OAI22_X1 U1391 ( .A1(n5177), .A2(n6396), .B1(n802), .B2(n233), .ZN(n3748) );
  OAI22_X1 U1392 ( .A1(n5145), .A2(n6393), .B1(n802), .B2(n235), .ZN(n3749) );
  OAI22_X1 U1393 ( .A1(n5113), .A2(n6391), .B1(n802), .B2(n237), .ZN(n3750) );
  OAI22_X1 U1394 ( .A1(n5081), .A2(n6390), .B1(n802), .B2(n239), .ZN(n3751) );
  OAI22_X1 U1395 ( .A1(n5049), .A2(n6388), .B1(n802), .B2(n241), .ZN(n3752) );
  OAI22_X1 U1396 ( .A1(n5017), .A2(n6385), .B1(n802), .B2(n243), .ZN(n3753) );
  OAI22_X1 U1397 ( .A1(n4985), .A2(n6383), .B1(n802), .B2(n245), .ZN(n3754) );
  OAI22_X1 U1398 ( .A1(n4953), .A2(n6382), .B1(n802), .B2(n247), .ZN(n3755) );
  OAI22_X1 U1399 ( .A1(n4921), .A2(n6380), .B1(n802), .B2(n249), .ZN(n3756) );
  OAI22_X1 U1400 ( .A1(n4889), .A2(n6384), .B1(n802), .B2(n251), .ZN(n3757) );
  OAI22_X1 U1401 ( .A1(n4857), .A2(n6381), .B1(n802), .B2(n253), .ZN(n3758) );
  OAI22_X1 U1402 ( .A1(n4825), .A2(n6387), .B1(n802), .B2(n255), .ZN(n3759) );
  OAI22_X1 U1403 ( .A1(n4793), .A2(n6386), .B1(n802), .B2(n257), .ZN(n3760) );
  OAI22_X1 U1404 ( .A1(n4761), .A2(n6392), .B1(n802), .B2(n259), .ZN(n3761) );
  OAI22_X1 U1405 ( .A1(n4729), .A2(n6394), .B1(n802), .B2(n261), .ZN(n3762) );
  OAI22_X1 U1406 ( .A1(n4697), .A2(n6389), .B1(n802), .B2(n263), .ZN(n3763) );
  OAI22_X1 U1407 ( .A1(n4665), .A2(n6395), .B1(n802), .B2(n265), .ZN(n3764) );
  OAI22_X1 U1408 ( .A1(n4633), .A2(n6400), .B1(n802), .B2(n267), .ZN(n3765) );
  OAI22_X1 U1409 ( .A1(n4601), .A2(n6402), .B1(n802), .B2(n269), .ZN(n3766) );
  OAI22_X1 U1410 ( .A1(n4569), .A2(n6397), .B1(n802), .B2(n271), .ZN(n3767) );
  OAI22_X1 U1411 ( .A1(n4537), .A2(n6403), .B1(n802), .B2(n273), .ZN(n3768) );
  OAI22_X1 U1412 ( .A1(n4505), .A2(n6408), .B1(n802), .B2(n275), .ZN(n3769) );
  OAI22_X1 U1413 ( .A1(n4473), .A2(n6405), .B1(n802), .B2(n277), .ZN(n3770) );
  OAI22_X1 U1414 ( .A1(n4441), .A2(n6411), .B1(n802), .B2(n279), .ZN(n3771) );
  OAI221_X1 U1415 ( .B1(n133), .B2(n803), .C1(n5694), .C2(n135), .A(n804), 
        .ZN(n3772) );
  AOI22_X1 U1416 ( .A1(n137), .A2(n805), .B1(\UUT/Mpath/the_mult/Mad_out [55]), 
        .B2(n139), .ZN(n804) );
  OAI221_X1 U1417 ( .B1(n140), .B2(n806), .C1(n5646), .C2(n142), .A(n807), 
        .ZN(n3773) );
  AOI22_X1 U1418 ( .A1(n144), .A2(n805), .B1(\UUT/Mpath/the_mult/Mad_out [23]), 
        .B2(n145), .ZN(n807) );
  INV_X1 U1419 ( .A(n5647), .ZN(n805) );
  OAI22_X1 U1420 ( .A1(net54911), .A2(n808), .B1(n5647), .B2(net54871), .ZN(
        n3774) );
  OAI221_X1 U1421 ( .B1(n809), .B2(n310), .C1(n147), .C2(n808), .A(n810), .ZN(
        n3775) );
  AOI22_X1 U1422 ( .A1(n312), .A2(n811), .B1(n314), .B2(n812), .ZN(n810) );
  INV_X1 U1423 ( .A(\UUT/Mpath/the_mult/x_operand1[23] ), .ZN(n808) );
  OAI221_X1 U1424 ( .B1(n809), .B2(n316), .C1(\UUT/Mpath/the_alu/N37 ), .C2(
        net54887), .A(n813), .ZN(n3776) );
  AOI22_X1 U1425 ( .A1(n318), .A2(n811), .B1(n319), .B2(n812), .ZN(n813) );
  OAI22_X1 U1426 ( .A1(n5397), .A2(n6407), .B1(n814), .B2(n219), .ZN(n3777) );
  OAI22_X1 U1427 ( .A1(n5365), .A2(n6410), .B1(n814), .B2(n221), .ZN(n3778) );
  OAI22_X1 U1428 ( .A1(n5333), .A2(n6401), .B1(n814), .B2(n223), .ZN(n3779) );
  OAI22_X1 U1429 ( .A1(n5301), .A2(n6406), .B1(n814), .B2(n225), .ZN(n3780) );
  OAI22_X1 U1430 ( .A1(n5269), .A2(n6399), .B1(n814), .B2(n227), .ZN(n3781) );
  OAI22_X1 U1431 ( .A1(n5237), .A2(n6404), .B1(n814), .B2(n229), .ZN(n3782) );
  OAI22_X1 U1432 ( .A1(n5205), .A2(n6398), .B1(n814), .B2(n231), .ZN(n3783) );
  OAI22_X1 U1433 ( .A1(n5173), .A2(n6396), .B1(n814), .B2(n233), .ZN(n3784) );
  OAI22_X1 U1434 ( .A1(n5141), .A2(n6393), .B1(n814), .B2(n235), .ZN(n3785) );
  OAI22_X1 U1435 ( .A1(n5109), .A2(n6391), .B1(n814), .B2(n237), .ZN(n3786) );
  OAI22_X1 U1436 ( .A1(n5077), .A2(n6390), .B1(n814), .B2(n239), .ZN(n3787) );
  OAI22_X1 U1437 ( .A1(n5045), .A2(n6388), .B1(n814), .B2(n241), .ZN(n3788) );
  OAI22_X1 U1438 ( .A1(n5013), .A2(n6385), .B1(n814), .B2(n243), .ZN(n3789) );
  OAI22_X1 U1439 ( .A1(n4981), .A2(n6383), .B1(n814), .B2(n245), .ZN(n3790) );
  OAI22_X1 U1440 ( .A1(n4949), .A2(n6382), .B1(n814), .B2(n247), .ZN(n3791) );
  OAI22_X1 U1441 ( .A1(n4917), .A2(n6380), .B1(n814), .B2(n249), .ZN(n3792) );
  OAI22_X1 U1442 ( .A1(n4885), .A2(n6384), .B1(n814), .B2(n251), .ZN(n3793) );
  OAI22_X1 U1443 ( .A1(n4853), .A2(n6381), .B1(n814), .B2(n253), .ZN(n3794) );
  OAI22_X1 U1444 ( .A1(n4821), .A2(n6387), .B1(n814), .B2(n255), .ZN(n3795) );
  OAI22_X1 U1445 ( .A1(n4789), .A2(n6386), .B1(n814), .B2(n257), .ZN(n3796) );
  OAI22_X1 U1446 ( .A1(n4757), .A2(n6392), .B1(n814), .B2(n259), .ZN(n3797) );
  OAI22_X1 U1447 ( .A1(n4725), .A2(n6394), .B1(n814), .B2(n261), .ZN(n3798) );
  OAI22_X1 U1448 ( .A1(n4693), .A2(n6389), .B1(n814), .B2(n263), .ZN(n3799) );
  OAI22_X1 U1449 ( .A1(n4661), .A2(n6395), .B1(n814), .B2(n265), .ZN(n3800) );
  OAI22_X1 U1450 ( .A1(n4629), .A2(n6400), .B1(n814), .B2(n267), .ZN(n3801) );
  OAI22_X1 U1451 ( .A1(n4597), .A2(n6402), .B1(n814), .B2(n269), .ZN(n3802) );
  OAI22_X1 U1452 ( .A1(n4565), .A2(n6397), .B1(n814), .B2(n271), .ZN(n3803) );
  OAI22_X1 U1453 ( .A1(n4533), .A2(n6403), .B1(n814), .B2(n273), .ZN(n3804) );
  OAI22_X1 U1454 ( .A1(n4501), .A2(n6408), .B1(n814), .B2(n275), .ZN(n3805) );
  OAI22_X1 U1455 ( .A1(n4469), .A2(n6405), .B1(n814), .B2(n277), .ZN(n3806) );
  OAI22_X1 U1456 ( .A1(n4437), .A2(n6411), .B1(n814), .B2(n279), .ZN(n3807) );
  OAI22_X1 U1457 ( .A1(net54909), .A2(n815), .B1(net54867), .B2(
        \UUT/Mpath/the_memhandle/N239 ), .ZN(n3808) );
  INV_X1 U1458 ( .A(\UUT/daddr_out [1]), .ZN(n815) );
  OAI222_X1 U1459 ( .A1(n84), .A2(n123), .B1(n787), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N82 ), .C2(net54895), .ZN(n3809) );
  INV_X1 U1460 ( .A(\UUT/break_code[1] ), .ZN(n787) );
  INV_X1 U1461 ( .A(n816), .ZN(n84) );
  OAI222_X1 U1462 ( .A1(n797), .A2(n129), .B1(n802), .B2(n131), .C1(n5493), 
        .C2(n132), .ZN(n816) );
  OAI211_X1 U1464 ( .C1(n5710), .C2(n5494), .A(n817), .B(n818), .ZN(n800) );
  AOI222_X1 U1465 ( .A1(n5712), .A2(n684), .B1(n685), .B2(n624), .C1(n5922), 
        .C2(n686), .ZN(n818) );
  INV_X1 U1466 ( .A(n5921), .ZN(n624) );
  AOI22_X1 U1467 ( .A1(n5923), .A2(n687), .B1(n5918), .B2(n688), .ZN(n817) );
  OAI22_X1 U1468 ( .A1(n5494), .A2(net54877), .B1(net54925), .B2(n797), .ZN(
        n3810) );
  INV_X1 U1469 ( .A(n819), .ZN(n797) );
  OAI211_X1 U1470 ( .C1(n5654), .C2(n321), .A(n820), .B(n821), .ZN(n819) );
  AOI222_X1 U1471 ( .A1(n285), .A2(n822), .B1(\UUT/Mpath/out_jar[1] ), .B2(
        n325), .C1(n284), .C2(n823), .ZN(n821) );
  INV_X1 U1472 ( .A(n5698), .ZN(n823) );
  AOI22_X1 U1473 ( .A1(n6379), .A2(\UUT/daddr_out [1]), .B1(
        \UUT/Mpath/the_mult/x_mult_out[1] ), .B2(n291), .ZN(n820) );
  OAI22_X1 U1474 ( .A1(\UUT/Mpath/the_alu/N33 ), .A2(net54877), .B1(net54925), 
        .B2(n201), .ZN(n3811) );
  INV_X1 U1475 ( .A(n824), .ZN(n201) );
  OAI222_X1 U1476 ( .A1(n5530), .A2(n194), .B1(n5528), .B2(n193), .C1(n6364), 
        .C2(n5420), .ZN(n824) );
  OAI22_X1 U1477 ( .A1(n5395), .A2(n6407), .B1(n194), .B2(n219), .ZN(n3812) );
  OAI22_X1 U1478 ( .A1(n5363), .A2(n6410), .B1(n194), .B2(n221), .ZN(n3813) );
  OAI22_X1 U1479 ( .A1(n5331), .A2(n6401), .B1(n194), .B2(n223), .ZN(n3814) );
  OAI22_X1 U1480 ( .A1(n5299), .A2(n6406), .B1(n194), .B2(n225), .ZN(n3815) );
  OAI22_X1 U1481 ( .A1(n5267), .A2(n6399), .B1(n194), .B2(n227), .ZN(n3816) );
  OAI22_X1 U1482 ( .A1(n5235), .A2(n6404), .B1(n194), .B2(n229), .ZN(n3817) );
  OAI22_X1 U1483 ( .A1(n5203), .A2(n6398), .B1(n194), .B2(n231), .ZN(n3818) );
  OAI22_X1 U1484 ( .A1(n5171), .A2(n6396), .B1(n194), .B2(n233), .ZN(n3819) );
  OAI22_X1 U1485 ( .A1(n5139), .A2(n6393), .B1(n194), .B2(n235), .ZN(n3820) );
  OAI22_X1 U1486 ( .A1(n5107), .A2(n6391), .B1(n194), .B2(n237), .ZN(n3821) );
  OAI22_X1 U1487 ( .A1(n5075), .A2(n6390), .B1(n194), .B2(n239), .ZN(n3822) );
  OAI22_X1 U1488 ( .A1(n5043), .A2(n6388), .B1(n194), .B2(n241), .ZN(n3823) );
  OAI22_X1 U1489 ( .A1(n5011), .A2(n6385), .B1(n194), .B2(n243), .ZN(n3824) );
  OAI22_X1 U1490 ( .A1(n4979), .A2(n6383), .B1(n194), .B2(n245), .ZN(n3825) );
  OAI22_X1 U1491 ( .A1(n4947), .A2(n6382), .B1(n194), .B2(n247), .ZN(n3826) );
  OAI22_X1 U1492 ( .A1(n4915), .A2(n6380), .B1(n194), .B2(n249), .ZN(n3827) );
  OAI22_X1 U1493 ( .A1(n4883), .A2(n6384), .B1(n194), .B2(n251), .ZN(n3828) );
  OAI22_X1 U1494 ( .A1(n4851), .A2(n6381), .B1(n194), .B2(n253), .ZN(n3829) );
  OAI22_X1 U1495 ( .A1(n4819), .A2(n6387), .B1(n194), .B2(n255), .ZN(n3830) );
  OAI22_X1 U1496 ( .A1(n4787), .A2(n6386), .B1(n194), .B2(n257), .ZN(n3831) );
  OAI22_X1 U1497 ( .A1(n4755), .A2(n6392), .B1(n194), .B2(n259), .ZN(n3832) );
  OAI22_X1 U1498 ( .A1(n4723), .A2(n6394), .B1(n194), .B2(n261), .ZN(n3833) );
  OAI22_X1 U1499 ( .A1(n4691), .A2(n6389), .B1(n194), .B2(n263), .ZN(n3834) );
  OAI22_X1 U1500 ( .A1(n4659), .A2(n6395), .B1(n194), .B2(n265), .ZN(n3835) );
  OAI22_X1 U1501 ( .A1(n4627), .A2(n6400), .B1(n194), .B2(n267), .ZN(n3836) );
  OAI22_X1 U1502 ( .A1(n4595), .A2(n6402), .B1(n194), .B2(n269), .ZN(n3837) );
  OAI22_X1 U1503 ( .A1(n4563), .A2(n6397), .B1(n194), .B2(n271), .ZN(n3838) );
  OAI22_X1 U1504 ( .A1(n4531), .A2(n6403), .B1(n194), .B2(n273), .ZN(n3839) );
  OAI22_X1 U1505 ( .A1(n4499), .A2(n6408), .B1(n194), .B2(n275), .ZN(n3840) );
  OAI22_X1 U1506 ( .A1(n4467), .A2(n6405), .B1(n194), .B2(n277), .ZN(n3841) );
  OAI22_X1 U1507 ( .A1(n4435), .A2(n6411), .B1(n194), .B2(n279), .ZN(n3842) );
  OAI22_X1 U1510 ( .A1(n5476), .A2(net54877), .B1(net54925), .B2(n193), .ZN(
        n3843) );
  AOI221_X1 U1511 ( .B1(n826), .B2(n284), .C1(n5598), .C2(n285), .A(n827), 
        .ZN(n193) );
  INV_X1 U1512 ( .A(n828), .ZN(n827) );
  AOI222_X1 U1513 ( .A1(n288), .A2(n829), .B1(n6379), .B2(n5599), .C1(
        \UUT/Mpath/the_mult/x_mult_out[25] ), .C2(n291), .ZN(n828) );
  INV_X1 U1514 ( .A(n5642), .ZN(n829) );
  INV_X1 U1515 ( .A(n5692), .ZN(n826) );
  OAI22_X1 U1516 ( .A1(\UUT/Mpath/the_alu/N31 ), .A2(net54879), .B1(net54925), 
        .B2(n188), .ZN(n3844) );
  INV_X1 U1517 ( .A(n830), .ZN(n188) );
  OAI222_X1 U1518 ( .A1(n5530), .A2(n181), .B1(n5528), .B2(n180), .C1(n6364), 
        .C2(n5419), .ZN(n830) );
  OAI22_X1 U1519 ( .A1(n5394), .A2(n6407), .B1(n181), .B2(n219), .ZN(n3845) );
  OAI22_X1 U1520 ( .A1(n5362), .A2(n6410), .B1(n181), .B2(n221), .ZN(n3846) );
  OAI22_X1 U1521 ( .A1(n5330), .A2(n6401), .B1(n181), .B2(n223), .ZN(n3847) );
  OAI22_X1 U1522 ( .A1(n5298), .A2(n6406), .B1(n181), .B2(n225), .ZN(n3848) );
  OAI22_X1 U1523 ( .A1(n5266), .A2(n6399), .B1(n181), .B2(n227), .ZN(n3849) );
  OAI22_X1 U1524 ( .A1(n5234), .A2(n6404), .B1(n181), .B2(n229), .ZN(n3850) );
  OAI22_X1 U1525 ( .A1(n5202), .A2(n6398), .B1(n181), .B2(n231), .ZN(n3851) );
  OAI22_X1 U1526 ( .A1(n5170), .A2(n6396), .B1(n181), .B2(n233), .ZN(n3852) );
  OAI22_X1 U1527 ( .A1(n5138), .A2(n6393), .B1(n181), .B2(n235), .ZN(n3853) );
  OAI22_X1 U1528 ( .A1(n5106), .A2(n6391), .B1(n181), .B2(n237), .ZN(n3854) );
  OAI22_X1 U1529 ( .A1(n5074), .A2(n6390), .B1(n181), .B2(n239), .ZN(n3855) );
  OAI22_X1 U1530 ( .A1(n5042), .A2(n6388), .B1(n181), .B2(n241), .ZN(n3856) );
  OAI22_X1 U1531 ( .A1(n5010), .A2(n6385), .B1(n181), .B2(n243), .ZN(n3857) );
  OAI22_X1 U1532 ( .A1(n4978), .A2(n6383), .B1(n181), .B2(n245), .ZN(n3858) );
  OAI22_X1 U1533 ( .A1(n4946), .A2(n6382), .B1(n181), .B2(n247), .ZN(n3859) );
  OAI22_X1 U1534 ( .A1(n4914), .A2(n6380), .B1(n181), .B2(n249), .ZN(n3860) );
  OAI22_X1 U1535 ( .A1(n4882), .A2(n6384), .B1(n181), .B2(n251), .ZN(n3861) );
  OAI22_X1 U1536 ( .A1(n4850), .A2(n6381), .B1(n181), .B2(n253), .ZN(n3862) );
  OAI22_X1 U1537 ( .A1(n4818), .A2(n6387), .B1(n181), .B2(n255), .ZN(n3863) );
  OAI22_X1 U1538 ( .A1(n4786), .A2(n6386), .B1(n181), .B2(n257), .ZN(n3864) );
  OAI22_X1 U1539 ( .A1(n4754), .A2(n6392), .B1(n181), .B2(n259), .ZN(n3865) );
  OAI22_X1 U1540 ( .A1(n4722), .A2(n6394), .B1(n181), .B2(n261), .ZN(n3866) );
  OAI22_X1 U1541 ( .A1(n4690), .A2(n6389), .B1(n181), .B2(n263), .ZN(n3867) );
  OAI22_X1 U1542 ( .A1(n4658), .A2(n6395), .B1(n181), .B2(n265), .ZN(n3868) );
  OAI22_X1 U1543 ( .A1(n4626), .A2(n6400), .B1(n181), .B2(n267), .ZN(n3869) );
  OAI22_X1 U1544 ( .A1(n4594), .A2(n6402), .B1(n181), .B2(n269), .ZN(n3870) );
  OAI22_X1 U1545 ( .A1(n4562), .A2(n6397), .B1(n181), .B2(n271), .ZN(n3871) );
  OAI22_X1 U1546 ( .A1(n4530), .A2(n6403), .B1(n181), .B2(n273), .ZN(n3872) );
  OAI22_X1 U1547 ( .A1(n4498), .A2(n6408), .B1(n181), .B2(n275), .ZN(n3873) );
  OAI22_X1 U1548 ( .A1(n4466), .A2(n6405), .B1(n181), .B2(n277), .ZN(n3874) );
  OAI22_X1 U1549 ( .A1(n4434), .A2(n6411), .B1(n181), .B2(n279), .ZN(n3875) );
  OAI22_X1 U1552 ( .A1(n5473), .A2(net54879), .B1(net54927), .B2(n180), .ZN(
        n3876) );
  AOI221_X1 U1553 ( .B1(n832), .B2(n284), .C1(n5591), .C2(n285), .A(n833), 
        .ZN(n180) );
  INV_X1 U1554 ( .A(n834), .ZN(n833) );
  AOI222_X1 U1555 ( .A1(n288), .A2(n835), .B1(n6379), .B2(n5592), .C1(
        \UUT/Mpath/the_mult/x_mult_out[26] ), .C2(n291), .ZN(n834) );
  INV_X1 U1556 ( .A(n5640), .ZN(n835) );
  INV_X1 U1557 ( .A(n5691), .ZN(n832) );
  OAI22_X1 U1558 ( .A1(\UUT/Mpath/the_alu/N29 ), .A2(net54879), .B1(net54927), 
        .B2(n172), .ZN(n3877) );
  INV_X1 U1559 ( .A(n836), .ZN(n172) );
  OAI222_X1 U1560 ( .A1(n5530), .A2(n165), .B1(n5528), .B2(n164), .C1(n6364), 
        .C2(n5418), .ZN(n836) );
  OAI22_X1 U1561 ( .A1(n5393), .A2(n6407), .B1(n165), .B2(n219), .ZN(n3878) );
  OAI22_X1 U1562 ( .A1(n5361), .A2(n6410), .B1(n165), .B2(n221), .ZN(n3879) );
  OAI22_X1 U1563 ( .A1(n5329), .A2(n6401), .B1(n165), .B2(n223), .ZN(n3880) );
  OAI22_X1 U1564 ( .A1(n5297), .A2(n6406), .B1(n165), .B2(n225), .ZN(n3881) );
  OAI22_X1 U1565 ( .A1(n5265), .A2(n6399), .B1(n165), .B2(n227), .ZN(n3882) );
  OAI22_X1 U1566 ( .A1(n5233), .A2(n6404), .B1(n165), .B2(n229), .ZN(n3883) );
  OAI22_X1 U1567 ( .A1(n5201), .A2(n6398), .B1(n165), .B2(n231), .ZN(n3884) );
  OAI22_X1 U1568 ( .A1(n5169), .A2(n6396), .B1(n165), .B2(n233), .ZN(n3885) );
  OAI22_X1 U1569 ( .A1(n5137), .A2(n6393), .B1(n165), .B2(n235), .ZN(n3886) );
  OAI22_X1 U1570 ( .A1(n5105), .A2(n6391), .B1(n165), .B2(n237), .ZN(n3887) );
  OAI22_X1 U1571 ( .A1(n5073), .A2(n6390), .B1(n165), .B2(n239), .ZN(n3888) );
  OAI22_X1 U1572 ( .A1(n5041), .A2(n6388), .B1(n165), .B2(n241), .ZN(n3889) );
  OAI22_X1 U1573 ( .A1(n5009), .A2(n6385), .B1(n165), .B2(n243), .ZN(n3890) );
  OAI22_X1 U1574 ( .A1(n4977), .A2(n6383), .B1(n165), .B2(n245), .ZN(n3891) );
  OAI22_X1 U1575 ( .A1(n4945), .A2(n6382), .B1(n165), .B2(n247), .ZN(n3892) );
  OAI22_X1 U1576 ( .A1(n4913), .A2(n6380), .B1(n165), .B2(n249), .ZN(n3893) );
  OAI22_X1 U1577 ( .A1(n4881), .A2(n6384), .B1(n165), .B2(n251), .ZN(n3894) );
  OAI22_X1 U1578 ( .A1(n4849), .A2(n6381), .B1(n165), .B2(n253), .ZN(n3895) );
  OAI22_X1 U1579 ( .A1(n4817), .A2(n6387), .B1(n165), .B2(n255), .ZN(n3896) );
  OAI22_X1 U1580 ( .A1(n4785), .A2(n6386), .B1(n165), .B2(n257), .ZN(n3897) );
  OAI22_X1 U1581 ( .A1(n4753), .A2(n6392), .B1(n165), .B2(n259), .ZN(n3898) );
  OAI22_X1 U1582 ( .A1(n4721), .A2(n6394), .B1(n165), .B2(n261), .ZN(n3899) );
  OAI22_X1 U1583 ( .A1(n4689), .A2(n6389), .B1(n165), .B2(n263), .ZN(n3900) );
  OAI22_X1 U1584 ( .A1(n4657), .A2(n6395), .B1(n165), .B2(n265), .ZN(n3901) );
  OAI22_X1 U1585 ( .A1(n4625), .A2(n6400), .B1(n165), .B2(n267), .ZN(n3902) );
  OAI22_X1 U1586 ( .A1(n4593), .A2(n6402), .B1(n165), .B2(n269), .ZN(n3903) );
  OAI22_X1 U1587 ( .A1(n4561), .A2(n6397), .B1(n165), .B2(n271), .ZN(n3904) );
  OAI22_X1 U1588 ( .A1(n4529), .A2(n6403), .B1(n165), .B2(n273), .ZN(n3905) );
  OAI22_X1 U1589 ( .A1(n4497), .A2(n6408), .B1(n165), .B2(n275), .ZN(n3906) );
  OAI22_X1 U1590 ( .A1(n4465), .A2(n6405), .B1(n165), .B2(n277), .ZN(n3907) );
  OAI22_X1 U1591 ( .A1(n4433), .A2(n6411), .B1(n165), .B2(n279), .ZN(n3908) );
  OAI22_X1 U1594 ( .A1(n5470), .A2(net54879), .B1(net54927), .B2(n164), .ZN(
        n3909) );
  AOI221_X1 U1595 ( .B1(n838), .B2(n284), .C1(n5584), .C2(n285), .A(n839), 
        .ZN(n164) );
  INV_X1 U1596 ( .A(n840), .ZN(n839) );
  AOI222_X1 U1597 ( .A1(n288), .A2(n841), .B1(n6379), .B2(n5585), .C1(
        \UUT/Mpath/the_mult/x_mult_out[27] ), .C2(n291), .ZN(n840) );
  INV_X1 U1598 ( .A(n5638), .ZN(n841) );
  INV_X1 U1599 ( .A(n5690), .ZN(n838) );
  OAI22_X1 U1600 ( .A1(\UUT/Mpath/the_alu/N27 ), .A2(net54879), .B1(net54927), 
        .B2(n160), .ZN(n3910) );
  INV_X1 U1601 ( .A(n842), .ZN(n160) );
  OAI222_X1 U1602 ( .A1(n5530), .A2(n153), .B1(n5528), .B2(n152), .C1(n6364), 
        .C2(n5417), .ZN(n842) );
  OAI22_X1 U1603 ( .A1(n5392), .A2(n6407), .B1(n153), .B2(n219), .ZN(n3911) );
  OAI22_X1 U1604 ( .A1(n5360), .A2(n6410), .B1(n153), .B2(n221), .ZN(n3912) );
  OAI22_X1 U1605 ( .A1(n5328), .A2(n6401), .B1(n153), .B2(n223), .ZN(n3913) );
  OAI22_X1 U1606 ( .A1(n5296), .A2(n6406), .B1(n153), .B2(n225), .ZN(n3914) );
  OAI22_X1 U1607 ( .A1(n5264), .A2(n6399), .B1(n153), .B2(n227), .ZN(n3915) );
  OAI22_X1 U1608 ( .A1(n5232), .A2(n6404), .B1(n153), .B2(n229), .ZN(n3916) );
  OAI22_X1 U1609 ( .A1(n5200), .A2(n6398), .B1(n153), .B2(n231), .ZN(n3917) );
  OAI22_X1 U1610 ( .A1(n5168), .A2(n6396), .B1(n153), .B2(n233), .ZN(n3918) );
  OAI22_X1 U1611 ( .A1(n5136), .A2(n6393), .B1(n153), .B2(n235), .ZN(n3919) );
  OAI22_X1 U1612 ( .A1(n5104), .A2(n6391), .B1(n153), .B2(n237), .ZN(n3920) );
  OAI22_X1 U1613 ( .A1(n5072), .A2(n6390), .B1(n153), .B2(n239), .ZN(n3921) );
  OAI22_X1 U1614 ( .A1(n5040), .A2(n6388), .B1(n153), .B2(n241), .ZN(n3922) );
  OAI22_X1 U1615 ( .A1(n5008), .A2(n6385), .B1(n153), .B2(n243), .ZN(n3923) );
  OAI22_X1 U1616 ( .A1(n4976), .A2(n6383), .B1(n153), .B2(n245), .ZN(n3924) );
  OAI22_X1 U1617 ( .A1(n4944), .A2(n6382), .B1(n153), .B2(n247), .ZN(n3925) );
  OAI22_X1 U1618 ( .A1(n4912), .A2(n6380), .B1(n153), .B2(n249), .ZN(n3926) );
  OAI22_X1 U1619 ( .A1(n4880), .A2(n6384), .B1(n153), .B2(n251), .ZN(n3927) );
  OAI22_X1 U1620 ( .A1(n4848), .A2(n6381), .B1(n153), .B2(n253), .ZN(n3928) );
  OAI22_X1 U1621 ( .A1(n4816), .A2(n6387), .B1(n153), .B2(n255), .ZN(n3929) );
  OAI22_X1 U1622 ( .A1(n4784), .A2(n6386), .B1(n153), .B2(n257), .ZN(n3930) );
  OAI22_X1 U1623 ( .A1(n4752), .A2(n6392), .B1(n153), .B2(n259), .ZN(n3931) );
  OAI22_X1 U1624 ( .A1(n4720), .A2(n6394), .B1(n153), .B2(n261), .ZN(n3932) );
  OAI22_X1 U1625 ( .A1(n4688), .A2(n6389), .B1(n153), .B2(n263), .ZN(n3933) );
  OAI22_X1 U1626 ( .A1(n4656), .A2(n6395), .B1(n153), .B2(n265), .ZN(n3934) );
  OAI22_X1 U1627 ( .A1(n4624), .A2(n6400), .B1(n153), .B2(n267), .ZN(n3935) );
  OAI22_X1 U1628 ( .A1(n4592), .A2(n6402), .B1(n153), .B2(n269), .ZN(n3936) );
  OAI22_X1 U1629 ( .A1(n4560), .A2(n6397), .B1(n153), .B2(n271), .ZN(n3937) );
  OAI22_X1 U1630 ( .A1(n4528), .A2(n6403), .B1(n153), .B2(n273), .ZN(n3938) );
  OAI22_X1 U1631 ( .A1(n4496), .A2(n6408), .B1(n153), .B2(n275), .ZN(n3939) );
  OAI22_X1 U1632 ( .A1(n4464), .A2(n6405), .B1(n153), .B2(n277), .ZN(n3940) );
  OAI22_X1 U1633 ( .A1(n4432), .A2(n6411), .B1(n153), .B2(n279), .ZN(n3941) );
  OAI22_X1 U1636 ( .A1(n5467), .A2(net54881), .B1(net54925), .B2(n152), .ZN(
        n3942) );
  AOI221_X1 U1637 ( .B1(n844), .B2(n284), .C1(n5577), .C2(n285), .A(n845), 
        .ZN(n152) );
  INV_X1 U1638 ( .A(n846), .ZN(n845) );
  AOI222_X1 U1639 ( .A1(n288), .A2(n847), .B1(n6379), .B2(n6452), .C1(
        \UUT/Mpath/the_mult/x_mult_out[28] ), .C2(n291), .ZN(n846) );
  INV_X1 U1640 ( .A(n5636), .ZN(n847) );
  INV_X1 U1641 ( .A(n5689), .ZN(n844) );
  OAI22_X1 U1642 ( .A1(\UUT/Mpath/the_alu/N25 ), .A2(net54881), .B1(net54925), 
        .B2(n148), .ZN(n3943) );
  INV_X1 U1643 ( .A(n848), .ZN(n148) );
  OAI222_X1 U1644 ( .A1(n5530), .A2(n130), .B1(n5528), .B2(n128), .C1(n6364), 
        .C2(n5416), .ZN(n848) );
  OAI22_X1 U1645 ( .A1(n5391), .A2(n6407), .B1(n130), .B2(n219), .ZN(n3944) );
  OAI22_X1 U1646 ( .A1(n5359), .A2(n6410), .B1(n130), .B2(n221), .ZN(n3945) );
  OAI22_X1 U1647 ( .A1(n5327), .A2(n6401), .B1(n130), .B2(n223), .ZN(n3946) );
  OAI22_X1 U1648 ( .A1(n5295), .A2(n6406), .B1(n130), .B2(n225), .ZN(n3947) );
  OAI22_X1 U1649 ( .A1(n5263), .A2(n6399), .B1(n130), .B2(n227), .ZN(n3948) );
  OAI22_X1 U1650 ( .A1(n5231), .A2(n6404), .B1(n130), .B2(n229), .ZN(n3949) );
  OAI22_X1 U1651 ( .A1(n5199), .A2(n6398), .B1(n130), .B2(n231), .ZN(n3950) );
  OAI22_X1 U1652 ( .A1(n5167), .A2(n6396), .B1(n130), .B2(n233), .ZN(n3951) );
  OAI22_X1 U1653 ( .A1(n5135), .A2(n6393), .B1(n130), .B2(n235), .ZN(n3952) );
  OAI22_X1 U1654 ( .A1(n5103), .A2(n6391), .B1(n130), .B2(n237), .ZN(n3953) );
  OAI22_X1 U1655 ( .A1(n5071), .A2(n6390), .B1(n130), .B2(n239), .ZN(n3954) );
  OAI22_X1 U1656 ( .A1(n5039), .A2(n6388), .B1(n130), .B2(n241), .ZN(n3955) );
  OAI22_X1 U1657 ( .A1(n5007), .A2(n6385), .B1(n130), .B2(n243), .ZN(n3956) );
  OAI22_X1 U1658 ( .A1(n4975), .A2(n6383), .B1(n130), .B2(n245), .ZN(n3957) );
  OAI22_X1 U1659 ( .A1(n4943), .A2(n6382), .B1(n130), .B2(n247), .ZN(n3958) );
  OAI22_X1 U1660 ( .A1(n4911), .A2(n6380), .B1(n130), .B2(n249), .ZN(n3959) );
  OAI22_X1 U1661 ( .A1(n4879), .A2(n6384), .B1(n130), .B2(n251), .ZN(n3960) );
  OAI22_X1 U1662 ( .A1(n4847), .A2(n6381), .B1(n130), .B2(n253), .ZN(n3961) );
  OAI22_X1 U1663 ( .A1(n4815), .A2(n6387), .B1(n130), .B2(n255), .ZN(n3962) );
  OAI22_X1 U1664 ( .A1(n4783), .A2(n6386), .B1(n130), .B2(n257), .ZN(n3963) );
  OAI22_X1 U1665 ( .A1(n4751), .A2(n6392), .B1(n130), .B2(n259), .ZN(n3964) );
  OAI22_X1 U1666 ( .A1(n4719), .A2(n6394), .B1(n130), .B2(n261), .ZN(n3965) );
  OAI22_X1 U1667 ( .A1(n4687), .A2(n6389), .B1(n130), .B2(n263), .ZN(n3966) );
  OAI22_X1 U1668 ( .A1(n4655), .A2(n6395), .B1(n130), .B2(n265), .ZN(n3967) );
  OAI22_X1 U1669 ( .A1(n4623), .A2(n6400), .B1(n130), .B2(n267), .ZN(n3968) );
  OAI22_X1 U1670 ( .A1(n4591), .A2(n6402), .B1(n130), .B2(n269), .ZN(n3969) );
  OAI22_X1 U1671 ( .A1(n4559), .A2(n6397), .B1(n130), .B2(n271), .ZN(n3970) );
  OAI22_X1 U1672 ( .A1(n4527), .A2(n6403), .B1(n130), .B2(n273), .ZN(n3971) );
  OAI22_X1 U1673 ( .A1(n4495), .A2(n6408), .B1(n130), .B2(n275), .ZN(n3972) );
  OAI22_X1 U1674 ( .A1(n4463), .A2(n6405), .B1(n130), .B2(n277), .ZN(n3973) );
  OAI22_X1 U1675 ( .A1(n4431), .A2(n6411), .B1(n130), .B2(n279), .ZN(n3974) );
  OAI22_X1 U1678 ( .A1(n5464), .A2(net54881), .B1(net54925), .B2(n128), .ZN(
        n3975) );
  AOI221_X1 U1679 ( .B1(n850), .B2(n284), .C1(n5570), .C2(n285), .A(n851), 
        .ZN(n128) );
  INV_X1 U1680 ( .A(n852), .ZN(n851) );
  AOI222_X1 U1681 ( .A1(n288), .A2(n853), .B1(n6379), .B2(n5571), .C1(
        \UUT/Mpath/the_mult/x_mult_out[29] ), .C2(n291), .ZN(n852) );
  INV_X1 U1682 ( .A(n5634), .ZN(n853) );
  INV_X1 U1683 ( .A(n5688), .ZN(n850) );
  OAI222_X1 U1684 ( .A1(n114), .A2(n123), .B1(net54933), .B2(n119), .C1(
        \UUT/Mpath/the_alu/N24 ), .C2(net54891), .ZN(n3976) );
  AOI21_X1 U1685 ( .B1(\UUT/Mcontrol/d_sampled_finstr [14]), .B2(n125), .A(
        n126), .ZN(n119) );
  OR2_X1 U1686 ( .A1(n176), .A2(n854), .ZN(n126) );
  OAI21_X1 U1687 ( .B1(n450), .B2(n855), .A(n856), .ZN(n176) );
  NOR2_X1 U1688 ( .A1(n857), .A2(n450), .ZN(n125) );
  INV_X1 U1689 ( .A(n858), .ZN(n114) );
  OAI222_X1 U1690 ( .A1(n859), .A2(n129), .B1(n860), .B2(n131), .C1(n5457), 
        .C2(n132), .ZN(n858) );
  OAI221_X1 U1693 ( .B1(n140), .B2(n864), .C1(n5630), .C2(n142), .A(n865), 
        .ZN(n3978) );
  AOI22_X1 U1694 ( .A1(n144), .A2(n863), .B1(\UUT/Mpath/the_mult/Mad_out [30]), 
        .B2(n145), .ZN(n865) );
  INV_X1 U1695 ( .A(n5631), .ZN(n863) );
  OAI22_X1 U1696 ( .A1(net54909), .A2(n866), .B1(n5631), .B2(net54873), .ZN(
        n3979) );
  OAI22_X1 U1697 ( .A1(n147), .A2(n866), .B1(n867), .B2(n6409), .ZN(n3980) );
  INV_X1 U1698 ( .A(\UUT/Mpath/the_mult/x_operand1[30] ), .ZN(n866) );
  OAI22_X1 U1699 ( .A1(\UUT/Mpath/the_alu/N23 ), .A2(net54883), .B1(net54925), 
        .B2(n867), .ZN(n3981) );
  INV_X1 U1700 ( .A(n868), .ZN(n867) );
  OAI222_X1 U1701 ( .A1(n5530), .A2(n860), .B1(n5528), .B2(n859), .C1(n6364), 
        .C2(n5415), .ZN(n868) );
  OAI22_X1 U1702 ( .A1(n5389), .A2(n6407), .B1(n860), .B2(n219), .ZN(n3982) );
  OAI22_X1 U1703 ( .A1(n5357), .A2(n6410), .B1(n860), .B2(n221), .ZN(n3983) );
  OAI22_X1 U1704 ( .A1(n5325), .A2(n6401), .B1(n860), .B2(n223), .ZN(n3984) );
  OAI22_X1 U1705 ( .A1(n5293), .A2(n6406), .B1(n860), .B2(n225), .ZN(n3985) );
  OAI22_X1 U1706 ( .A1(n5261), .A2(n6399), .B1(n860), .B2(n227), .ZN(n3986) );
  OAI22_X1 U1707 ( .A1(n5229), .A2(n6404), .B1(n860), .B2(n229), .ZN(n3987) );
  OAI22_X1 U1708 ( .A1(n5197), .A2(n6398), .B1(n860), .B2(n231), .ZN(n3988) );
  OAI22_X1 U1709 ( .A1(n5165), .A2(n6396), .B1(n860), .B2(n233), .ZN(n3989) );
  OAI22_X1 U1710 ( .A1(n5133), .A2(n6393), .B1(n860), .B2(n235), .ZN(n3990) );
  OAI22_X1 U1711 ( .A1(n5101), .A2(n6391), .B1(n860), .B2(n237), .ZN(n3991) );
  OAI22_X1 U1712 ( .A1(n5069), .A2(n6390), .B1(n860), .B2(n239), .ZN(n3992) );
  OAI22_X1 U1713 ( .A1(n5037), .A2(n6388), .B1(n860), .B2(n241), .ZN(n3993) );
  OAI22_X1 U1714 ( .A1(n5005), .A2(n6385), .B1(n860), .B2(n243), .ZN(n3994) );
  OAI22_X1 U1715 ( .A1(n4973), .A2(n6383), .B1(n860), .B2(n245), .ZN(n3995) );
  OAI22_X1 U1716 ( .A1(n4941), .A2(n6382), .B1(n860), .B2(n247), .ZN(n3996) );
  OAI22_X1 U1717 ( .A1(n4909), .A2(n6380), .B1(n860), .B2(n249), .ZN(n3997) );
  OAI22_X1 U1718 ( .A1(n4877), .A2(n6384), .B1(n860), .B2(n251), .ZN(n3998) );
  OAI22_X1 U1719 ( .A1(n4845), .A2(n6381), .B1(n860), .B2(n253), .ZN(n3999) );
  OAI22_X1 U1720 ( .A1(n4813), .A2(n6387), .B1(n860), .B2(n255), .ZN(n4000) );
  OAI22_X1 U1721 ( .A1(n4781), .A2(n6386), .B1(n860), .B2(n257), .ZN(n4001) );
  OAI22_X1 U1722 ( .A1(n4749), .A2(n6392), .B1(n860), .B2(n259), .ZN(n4002) );
  OAI22_X1 U1723 ( .A1(n4717), .A2(n6394), .B1(n860), .B2(n261), .ZN(n4003) );
  OAI22_X1 U1724 ( .A1(n4685), .A2(n6389), .B1(n860), .B2(n263), .ZN(n4004) );
  OAI22_X1 U1725 ( .A1(n4653), .A2(n6395), .B1(n860), .B2(n265), .ZN(n4005) );
  OAI22_X1 U1726 ( .A1(n4621), .A2(n6400), .B1(n860), .B2(n267), .ZN(n4006) );
  OAI22_X1 U1727 ( .A1(n4589), .A2(n6402), .B1(n860), .B2(n269), .ZN(n4007) );
  OAI22_X1 U1728 ( .A1(n4557), .A2(n6397), .B1(n860), .B2(n271), .ZN(n4008) );
  OAI22_X1 U1729 ( .A1(n4525), .A2(n6403), .B1(n860), .B2(n273), .ZN(n4009) );
  OAI22_X1 U1730 ( .A1(n4493), .A2(n6408), .B1(n860), .B2(n275), .ZN(n4010) );
  OAI22_X1 U1731 ( .A1(n4461), .A2(n6405), .B1(n860), .B2(n277), .ZN(n4011) );
  OAI22_X1 U1732 ( .A1(n4429), .A2(n6411), .B1(n860), .B2(n279), .ZN(n4012) );
  OAI22_X1 U1735 ( .A1(n5458), .A2(net54883), .B1(net54925), .B2(n859), .ZN(
        n4013) );
  AOI221_X1 U1736 ( .B1(n870), .B2(n284), .C1(n5562), .C2(n285), .A(n871), 
        .ZN(n859) );
  INV_X1 U1737 ( .A(n872), .ZN(n871) );
  AOI222_X1 U1738 ( .A1(n288), .A2(n873), .B1(n6379), .B2(n6542), .C1(
        \UUT/Mpath/the_mult/x_mult_out[30] ), .C2(n291), .ZN(n872) );
  INV_X1 U1739 ( .A(n5630), .ZN(n873) );
  INV_X1 U1740 ( .A(n5686), .ZN(n870) );
  OAI222_X1 U1741 ( .A1(n104), .A2(n123), .B1(n117), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N38 ), .C2(net54891), .ZN(n4014) );
  INV_X1 U1742 ( .A(n874), .ZN(n104) );
  OAI222_X1 U1743 ( .A1(n809), .A2(n129), .B1(n814), .B2(n131), .C1(n5481), 
        .C2(n132), .ZN(n874) );
  OAI221_X1 U1745 ( .B1(n5760), .B2(n281), .C1(n5710), .C2(n5482), .A(n282), 
        .ZN(n812) );
  OAI22_X1 U1746 ( .A1(n5482), .A2(net54885), .B1(net54925), .B2(n809), .ZN(
        n4015) );
  INV_X1 U1747 ( .A(n875), .ZN(n809) );
  OAI211_X1 U1748 ( .C1(n5646), .C2(n321), .A(n876), .B(n877), .ZN(n875) );
  AOI222_X1 U1749 ( .A1(n285), .A2(n878), .B1(\UUT/Mpath/out_jar[23] ), .B2(
        n325), .C1(n284), .C2(n879), .ZN(n877) );
  INV_X1 U1750 ( .A(n5694), .ZN(n879) );
  AOI22_X1 U1751 ( .A1(n6379), .A2(n6092), .B1(
        \UUT/Mpath/the_mult/x_mult_out[23] ), .B2(n291), .ZN(n876) );
  INV_X1 U1752 ( .A(n880), .ZN(n4016) );
  AOI22_X1 U1753 ( .A1(net54847), .A2(\UUT/jar_in [23]), .B1(net54933), .B2(
        \UUT/Mpath/out_jar[23] ), .ZN(n880) );
  INV_X1 U1754 ( .A(n881), .ZN(n4017) );
  AOI22_X1 U1755 ( .A1(net54843), .A2(\UUT/jar_in [22]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[22] ), .ZN(n881) );
  INV_X1 U1756 ( .A(n882), .ZN(n4018) );
  AOI22_X1 U1757 ( .A1(net54843), .A2(\UUT/jar_in [21]), .B1(net54933), .B2(
        \UUT/Mpath/out_jar[21] ), .ZN(n882) );
  INV_X1 U1758 ( .A(n883), .ZN(n4019) );
  AOI22_X1 U1759 ( .A1(net54843), .A2(\UUT/jar_in [20]), .B1(net54933), .B2(
        \UUT/Mpath/out_jar[20] ), .ZN(n883) );
  INV_X1 U1760 ( .A(n884), .ZN(n4020) );
  AOI22_X1 U1761 ( .A1(net54843), .A2(\UUT/jar_in [19]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[19] ), .ZN(n884) );
  INV_X1 U1762 ( .A(n885), .ZN(n4021) );
  AOI22_X1 U1763 ( .A1(net54843), .A2(\UUT/jar_in [18]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[18] ), .ZN(n885) );
  INV_X1 U1764 ( .A(n886), .ZN(n4022) );
  AOI22_X1 U1765 ( .A1(net54843), .A2(\UUT/jar_in [17]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[17] ), .ZN(n886) );
  INV_X1 U1766 ( .A(n887), .ZN(n4023) );
  AOI22_X1 U1767 ( .A1(net54843), .A2(\UUT/jar_in [16]), .B1(net54933), .B2(
        \UUT/Mpath/out_jar[16] ), .ZN(n887) );
  INV_X1 U1768 ( .A(n888), .ZN(n4024) );
  AOI22_X1 U1769 ( .A1(net54843), .A2(\UUT/jar_in [15]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[15] ), .ZN(n888) );
  INV_X1 U1770 ( .A(n889), .ZN(n4025) );
  AOI22_X1 U1771 ( .A1(net54843), .A2(\UUT/jar_in [14]), .B1(net54933), .B2(
        \UUT/Mpath/out_jar[14] ), .ZN(n889) );
  INV_X1 U1772 ( .A(n890), .ZN(n4026) );
  AOI22_X1 U1773 ( .A1(net54843), .A2(\UUT/jar_in [13]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[13] ), .ZN(n890) );
  INV_X1 U1774 ( .A(n891), .ZN(n4027) );
  AOI22_X1 U1775 ( .A1(net54843), .A2(\UUT/jar_in [12]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[12] ), .ZN(n891) );
  INV_X1 U1776 ( .A(n892), .ZN(n4028) );
  AOI22_X1 U1777 ( .A1(net54845), .A2(\UUT/jar_in [11]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[11] ), .ZN(n892) );
  INV_X1 U1778 ( .A(n893), .ZN(n4029) );
  AOI22_X1 U1779 ( .A1(net54845), .A2(\UUT/jar_in [10]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[10] ), .ZN(n893) );
  INV_X1 U1780 ( .A(n894), .ZN(n4030) );
  AOI22_X1 U1781 ( .A1(net54845), .A2(\UUT/jar_in [9]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[9] ), .ZN(n894) );
  INV_X1 U1782 ( .A(n895), .ZN(n4031) );
  AOI22_X1 U1783 ( .A1(net54845), .A2(\UUT/jar_in [8]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[8] ), .ZN(n895) );
  INV_X1 U1784 ( .A(n896), .ZN(n4032) );
  AOI22_X1 U1785 ( .A1(net54845), .A2(\UUT/jar_in [7]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[7] ), .ZN(n896) );
  INV_X1 U1786 ( .A(n897), .ZN(n4033) );
  AOI22_X1 U1787 ( .A1(net54845), .A2(\UUT/jar_in [6]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[6] ), .ZN(n897) );
  INV_X1 U1788 ( .A(n898), .ZN(n4034) );
  AOI22_X1 U1789 ( .A1(net54845), .A2(\UUT/jar_in [5]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[5] ), .ZN(n898) );
  INV_X1 U1790 ( .A(n899), .ZN(n4035) );
  AOI22_X1 U1791 ( .A1(net54845), .A2(\UUT/jar_in [4]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[4] ), .ZN(n899) );
  INV_X1 U1792 ( .A(n900), .ZN(n4036) );
  AOI22_X1 U1793 ( .A1(net54845), .A2(\UUT/jar_in [3]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[3] ), .ZN(n900) );
  INV_X1 U1794 ( .A(n901), .ZN(n4037) );
  AOI22_X1 U1795 ( .A1(net54845), .A2(\UUT/jar_in [2]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[2] ), .ZN(n901) );
  INV_X1 U1796 ( .A(n902), .ZN(n4038) );
  AOI22_X1 U1797 ( .A1(net54845), .A2(\UUT/jar_in [1]), .B1(net54937), .B2(
        \UUT/Mpath/out_jar[1] ), .ZN(n902) );
  OAI221_X1 U1798 ( .B1(n68), .B2(n294), .C1(n295), .C2(n2725), .A(n903), .ZN(
        n4039) );
  AOI22_X1 U1799 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [0]), .A2(n6511), 
        .B1(\UUT/jar_in [0]), .B2(n6711), .ZN(n903) );
  INV_X1 U1800 ( .A(n904), .ZN(n4040) );
  AOI22_X1 U1801 ( .A1(net54845), .A2(\UUT/jar_in [0]), .B1(net54935), .B2(
        \UUT/Mpath/out_jar[0] ), .ZN(n904) );
  NOR2_X1 U1805 ( .A1(n546), .A2(\UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(
        n298) );
  NAND2_X1 U1807 ( .A1(n908), .A2(n295), .ZN(n294) );
  OAI22_X1 U1808 ( .A1(n6642), .A2(n546), .B1(n295), .B2(n2728), .ZN(n4042) );
  OAI221_X1 U1809 ( .B1(n5428), .B2(n910), .C1(\UUT/Mpath/the_alu/N468 ), .C2(
        net54889), .A(n911), .ZN(n4043) );
  NAND3_X1 U1810 ( .A1(n912), .A2(net54869), .A3(n913), .ZN(n911) );
  NAND3_X1 U1811 ( .A1(n914), .A2(n915), .A3(n916), .ZN(n912) );
  OAI21_X1 U1812 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2071 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A(n917), .ZN(n916) );
  OAI21_X1 U1813 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2054 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N2061 ), .A(
        \UUT/Mcontrol/Operation_decoding32/N2066 ), .ZN(n917) );
  NAND3_X1 U1814 ( .A1(n918), .A2(\UUT/Mcontrol/Operation_decoding32/N2060 ), 
        .A3(n6077), .ZN(n914) );
  INV_X1 U1815 ( .A(n919), .ZN(n918) );
  AOI21_X1 U1816 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2047 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N2071 ), .A(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .ZN(n919) );
  OAI221_X1 U1817 ( .B1(n5427), .B2(n910), .C1(\UUT/Mpath/the_alu/N467 ), .C2(
        net54889), .A(n920), .ZN(n4044) );
  NAND4_X1 U1818 ( .A1(n921), .A2(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
        .A3(n922), .A4(net54859), .ZN(n920) );
  NAND2_X1 U1819 ( .A1(n923), .A2(n924), .ZN(n922) );
  OAI221_X1 U1820 ( .B1(n5426), .B2(n910), .C1(net54889), .C2(n2729), .A(n925), 
        .ZN(n4045) );
  OAI221_X1 U1821 ( .B1(n5425), .B2(n910), .C1(net54891), .C2(n2730), .A(n925), 
        .ZN(n4046) );
  NAND3_X1 U1822 ( .A1(net54875), .A2(n926), .A3(n927), .ZN(n925) );
  OAI221_X1 U1823 ( .B1(n5424), .B2(n910), .C1(\UUT/Mpath/the_alu/N453 ), .C2(
        net54887), .A(n928), .ZN(n4047) );
  NAND4_X1 U1824 ( .A1(n929), .A2(n930), .A3(net54859), .A4(n6030), .ZN(n928)
         );
  NAND3_X1 U1825 ( .A1(n6074), .A2(n931), .A3(n932), .ZN(n930) );
  NAND2_X1 U1826 ( .A1(net54877), .A2(n933), .ZN(n910) );
  OAI22_X1 U1827 ( .A1(\UUT/Mpath/the_alu/N466 ), .A2(net54881), .B1(net54925), 
        .B2(n934), .ZN(n4048) );
  AOI22_X1 U1828 ( .A1(n935), .A2(n936), .B1(
        \UUT/Mcontrol/d_sampled_finstr [5]), .B2(n933), .ZN(n934) );
  NAND2_X1 U1829 ( .A1(n923), .A2(n937), .ZN(n936) );
  INV_X1 U1830 ( .A(n926), .ZN(n923) );
  OAI21_X1 U1831 ( .B1(n6076), .B2(n6074), .A(n931), .ZN(n926) );
  NOR2_X1 U1832 ( .A1(n938), .A2(n939), .ZN(n4049) );
  AOI22_X1 U1833 ( .A1(\UUT/shift_op [0]), .A2(net54903), .B1(net54877), .B2(
        \UUT/Mcontrol/d_sampled_finstr [0]), .ZN(n939) );
  NOR2_X1 U1834 ( .A1(n938), .A2(n940), .ZN(n4050) );
  AOI22_X1 U1835 ( .A1(\UUT/shift_op [1]), .A2(net54903), .B1(net54877), .B2(
        \UUT/Mcontrol/d_sampled_finstr [1]), .ZN(n940) );
  NOR2_X1 U1836 ( .A1(n938), .A2(n941), .ZN(n4051) );
  AOI22_X1 U1837 ( .A1(\UUT/shift_op [2]), .A2(net54903), .B1(net54877), .B2(
        \UUT/Mcontrol/d_sampled_finstr [2]), .ZN(n941) );
  AND2_X1 U1838 ( .A1(n942), .A2(net54895), .ZN(n938) );
  OAI211_X1 U1839 ( .C1(\UUT/Mcontrol/Operation_decoding32/N2037 ), .C2(n943), 
        .A(n6028), .B(n927), .ZN(n942) );
  OAI22_X1 U1840 ( .A1(net54847), .A2(n944), .B1(n6071), .B2(n945), .ZN(n4052)
         );
  INV_X1 U1841 ( .A(\UUT/exe_outsel [0]), .ZN(n944) );
  OAI22_X1 U1842 ( .A1(net54847), .A2(\UUT/Mpath/N116 ), .B1(n6070), .B2(n945), 
        .ZN(n4053) );
  OAI221_X1 U1843 ( .B1(n140), .B2(n946), .C1(n5628), .C2(n142), .A(n947), 
        .ZN(n4054) );
  AOI22_X1 U1844 ( .A1(n144), .A2(n948), .B1(\UUT/Mpath/the_mult/Mad_out [31]), 
        .B2(n145), .ZN(n947) );
  OAI22_X1 U1845 ( .A1(net54909), .A2(n949), .B1(n5629), .B2(net54871), .ZN(
        n4055) );
  OAI22_X1 U1846 ( .A1(n147), .A2(n949), .B1(n950), .B2(n6409), .ZN(n4056) );
  INV_X1 U1847 ( .A(\UUT/Mpath/the_mult/x_operand1[31] ), .ZN(n949) );
  OAI22_X1 U1848 ( .A1(\UUT/Mpath/the_alu/N21 ), .A2(net54879), .B1(net54921), 
        .B2(n950), .ZN(n4057) );
  INV_X1 U1849 ( .A(n951), .ZN(n950) );
  OAI222_X1 U1850 ( .A1(n5530), .A2(n952), .B1(n5528), .B2(n953), .C1(n6364), 
        .C2(n5414), .ZN(n951) );
  OAI22_X1 U1851 ( .A1(net54909), .A2(n954), .B1(net54865), .B2(
        \UUT/Mpath/the_memhandle/N236 ), .ZN(n4058) );
  INV_X1 U1852 ( .A(dmem_isbyte), .ZN(n954) );
  OAI22_X1 U1853 ( .A1(net54909), .A2(n955), .B1(net54865), .B2(
        \UUT/Mpath/the_memhandle/N238 ), .ZN(n4059) );
  INV_X1 U1854 ( .A(dmem_ishalf), .ZN(n955) );
  OAI22_X1 U1855 ( .A1(net54909), .A2(n956), .B1(n5710), .B2(net54871), .ZN(
        n4060) );
  INV_X1 U1856 ( .A(dmem_read), .ZN(n956) );
  OAI21_X1 U1857 ( .B1(net54847), .B2(\UUT/Mpath/the_memhandle/N235 ), .A(n957), .ZN(n4063) );
  OAI21_X1 U1858 ( .B1(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), .B2(
        \UUT/x_we ), .A(net54859), .ZN(n957) );
  OAI22_X1 U1859 ( .A1(n4678), .A2(n6389), .B1(n958), .B2(n263), .ZN(n4064) );
  OAI22_X1 U1860 ( .A1(n4684), .A2(n6389), .B1(n952), .B2(n263), .ZN(n4065) );
  OAI22_X1 U1861 ( .A1(n4707), .A2(n6389), .B1(n959), .B2(n263), .ZN(n4066) );
  OAI22_X1 U1862 ( .A1(n4708), .A2(n262), .B1(n960), .B2(n263), .ZN(n4067) );
  NOR3_X1 U1864 ( .A1(\UUT/regfile/N451 ), .A2(net54927), .A3(n961), .ZN(n262)
         );
  OAI22_X1 U1865 ( .A1(n4774), .A2(n6386), .B1(n958), .B2(n257), .ZN(n4068) );
  OAI22_X1 U1866 ( .A1(n4780), .A2(n6386), .B1(n952), .B2(n257), .ZN(n4069) );
  OAI22_X1 U1867 ( .A1(n4803), .A2(n6386), .B1(n959), .B2(n257), .ZN(n4070) );
  OAI22_X1 U1868 ( .A1(n4804), .A2(n256), .B1(n960), .B2(n257), .ZN(n4071) );
  NOR3_X1 U1870 ( .A1(\UUT/regfile/N439 ), .A2(net54927), .A3(n962), .ZN(n256)
         );
  OAI22_X1 U1871 ( .A1(n4838), .A2(n6381), .B1(n958), .B2(n253), .ZN(n4072) );
  OAI22_X1 U1872 ( .A1(n4844), .A2(n6381), .B1(n952), .B2(n253), .ZN(n4073) );
  OAI22_X1 U1873 ( .A1(n4867), .A2(n6381), .B1(n959), .B2(n253), .ZN(n4074) );
  OAI22_X1 U1874 ( .A1(n4868), .A2(n252), .B1(n960), .B2(n253), .ZN(n4075) );
  NOR3_X1 U1876 ( .A1(\UUT/regfile/N427 ), .A2(net54929), .A3(n961), .ZN(n252)
         );
  OAI22_X1 U1877 ( .A1(n4902), .A2(n6380), .B1(n958), .B2(n249), .ZN(n4076) );
  OAI22_X1 U1878 ( .A1(n4908), .A2(n6380), .B1(n952), .B2(n249), .ZN(n4077) );
  OAI22_X1 U1879 ( .A1(n4931), .A2(n6380), .B1(n959), .B2(n249), .ZN(n4078) );
  OAI22_X1 U1880 ( .A1(n4932), .A2(n248), .B1(n960), .B2(n249), .ZN(n4079) );
  NOR3_X1 U1882 ( .A1(\UUT/regfile/N415 ), .A2(net54929), .A3(n962), .ZN(n248)
         );
  OAI22_X1 U1883 ( .A1(n4966), .A2(n6383), .B1(n958), .B2(n245), .ZN(n4080) );
  OAI22_X1 U1884 ( .A1(n4972), .A2(n6383), .B1(n952), .B2(n245), .ZN(n4081) );
  OAI22_X1 U1885 ( .A1(n4995), .A2(n6383), .B1(n959), .B2(n245), .ZN(n4082) );
  OAI22_X1 U1886 ( .A1(n4996), .A2(n244), .B1(n960), .B2(n245), .ZN(n4083) );
  NOR3_X1 U1888 ( .A1(\UUT/regfile/N403 ), .A2(net54929), .A3(n961), .ZN(n244)
         );
  OAI22_X1 U1889 ( .A1(n5030), .A2(n6388), .B1(n958), .B2(n241), .ZN(n4084) );
  OAI22_X1 U1890 ( .A1(n5036), .A2(n6388), .B1(n952), .B2(n241), .ZN(n4085) );
  OAI22_X1 U1891 ( .A1(n5059), .A2(n6388), .B1(n959), .B2(n241), .ZN(n4086) );
  OAI22_X1 U1892 ( .A1(n5060), .A2(n240), .B1(n960), .B2(n241), .ZN(n4087) );
  NOR3_X1 U1894 ( .A1(\UUT/regfile/N391 ), .A2(net54931), .A3(n962), .ZN(n240)
         );
  OAI22_X1 U1895 ( .A1(n5126), .A2(n6393), .B1(n958), .B2(n235), .ZN(n4088) );
  OAI22_X1 U1896 ( .A1(n5132), .A2(n6393), .B1(n952), .B2(n235), .ZN(n4089) );
  OAI22_X1 U1897 ( .A1(n5155), .A2(n6393), .B1(n959), .B2(n235), .ZN(n4090) );
  OAI22_X1 U1898 ( .A1(n5156), .A2(n234), .B1(n960), .B2(n235), .ZN(n4091) );
  NOR3_X1 U1900 ( .A1(\UUT/regfile/N379 ), .A2(net54927), .A3(n961), .ZN(n234)
         );
  OAI22_X1 U1901 ( .A1(n5190), .A2(n6398), .B1(n958), .B2(n231), .ZN(n4092) );
  OAI22_X1 U1902 ( .A1(n5196), .A2(n6398), .B1(n952), .B2(n231), .ZN(n4093) );
  OAI22_X1 U1903 ( .A1(n5219), .A2(n6398), .B1(n959), .B2(n231), .ZN(n4094) );
  OAI22_X1 U1904 ( .A1(n5220), .A2(n230), .B1(n960), .B2(n231), .ZN(n4095) );
  NOR3_X1 U1906 ( .A1(\UUT/regfile/N367 ), .A2(net54927), .A3(n962), .ZN(n230)
         );
  OAI22_X1 U1907 ( .A1(n5254), .A2(n6399), .B1(n958), .B2(n227), .ZN(n4096) );
  OAI22_X1 U1908 ( .A1(n5260), .A2(n6399), .B1(n952), .B2(n227), .ZN(n4097) );
  OAI22_X1 U1909 ( .A1(n5283), .A2(n6399), .B1(n959), .B2(n227), .ZN(n4098) );
  OAI22_X1 U1910 ( .A1(n5284), .A2(n226), .B1(n960), .B2(n227), .ZN(n4099) );
  NOR3_X1 U1912 ( .A1(\UUT/regfile/N354 ), .A2(net54927), .A3(n961), .ZN(n226)
         );
  OAI22_X1 U1913 ( .A1(n5318), .A2(n6401), .B1(n958), .B2(n223), .ZN(n4100) );
  OAI22_X1 U1914 ( .A1(n5324), .A2(n6401), .B1(n952), .B2(n223), .ZN(n4101) );
  OAI22_X1 U1915 ( .A1(n5347), .A2(n6401), .B1(n959), .B2(n223), .ZN(n4102) );
  OAI22_X1 U1916 ( .A1(n5348), .A2(n222), .B1(n960), .B2(n223), .ZN(n4103) );
  NOR3_X1 U1918 ( .A1(\UUT/regfile/N342 ), .A2(net54931), .A3(n962), .ZN(n222)
         );
  OAI22_X1 U1919 ( .A1(n5382), .A2(n6407), .B1(n958), .B2(n219), .ZN(n4104) );
  OAI22_X1 U1920 ( .A1(n5388), .A2(n6407), .B1(n952), .B2(n219), .ZN(n4105) );
  OAI22_X1 U1921 ( .A1(n5411), .A2(n6407), .B1(n959), .B2(n219), .ZN(n4106) );
  OAI22_X1 U1922 ( .A1(n5412), .A2(n218), .B1(n960), .B2(n219), .ZN(n4107) );
  NOR3_X1 U1924 ( .A1(\UUT/regfile/N330 ), .A2(net54929), .A3(n961), .ZN(n218)
         );
  OAI22_X1 U1925 ( .A1(n4454), .A2(n6405), .B1(n958), .B2(n277), .ZN(n4108) );
  OAI22_X1 U1926 ( .A1(n4460), .A2(n6405), .B1(n952), .B2(n277), .ZN(n4109) );
  OAI22_X1 U1927 ( .A1(n4483), .A2(n6405), .B1(n959), .B2(n277), .ZN(n4110) );
  OAI22_X1 U1928 ( .A1(n4484), .A2(n276), .B1(n960), .B2(n277), .ZN(n4111) );
  NOR3_X1 U1930 ( .A1(\UUT/regfile/N318 ), .A2(net54929), .A3(n962), .ZN(n276)
         );
  OAI22_X1 U1931 ( .A1(n4518), .A2(n6403), .B1(n958), .B2(n273), .ZN(n4112) );
  OAI22_X1 U1932 ( .A1(n4524), .A2(n6403), .B1(n952), .B2(n273), .ZN(n4113) );
  OAI22_X1 U1933 ( .A1(n4547), .A2(n6403), .B1(n959), .B2(n273), .ZN(n4114) );
  OAI22_X1 U1934 ( .A1(n4548), .A2(n272), .B1(n960), .B2(n273), .ZN(n4115) );
  NOR3_X1 U1936 ( .A1(\UUT/regfile/N305 ), .A2(net54927), .A3(n961), .ZN(n272)
         );
  OAI22_X1 U1937 ( .A1(n4582), .A2(n6402), .B1(n958), .B2(n269), .ZN(n4116) );
  OAI22_X1 U1938 ( .A1(n4588), .A2(n6402), .B1(n952), .B2(n269), .ZN(n4117) );
  OAI22_X1 U1939 ( .A1(n4611), .A2(n6402), .B1(n959), .B2(n269), .ZN(n4118) );
  OAI22_X1 U1940 ( .A1(n4612), .A2(n268), .B1(n960), .B2(n269), .ZN(n4119) );
  NOR3_X1 U1942 ( .A1(\UUT/regfile/N293 ), .A2(net54931), .A3(n962), .ZN(n268)
         );
  NAND2_X1 U1943 ( .A1(n963), .A2(n964), .ZN(n962) );
  OAI22_X1 U1944 ( .A1(n4710), .A2(n6394), .B1(n958), .B2(n261), .ZN(n4120) );
  OAI22_X1 U1945 ( .A1(n4716), .A2(n6394), .B1(n952), .B2(n261), .ZN(n4121) );
  OAI22_X1 U1946 ( .A1(n4739), .A2(n6394), .B1(n959), .B2(n261), .ZN(n4122) );
  OAI22_X1 U1947 ( .A1(n4740), .A2(n260), .B1(n960), .B2(n261), .ZN(n4123) );
  NOR3_X1 U1949 ( .A1(\UUT/regfile/N280 ), .A2(net54929), .A3(n961), .ZN(n260)
         );
  NAND2_X1 U1950 ( .A1(\UUT/rd_addr [1]), .A2(n964), .ZN(n961) );
  OAI22_X1 U1951 ( .A1(n4646), .A2(n6395), .B1(n958), .B2(n265), .ZN(n4124) );
  OAI22_X1 U1952 ( .A1(n4652), .A2(n6395), .B1(n952), .B2(n265), .ZN(n4125) );
  OAI22_X1 U1953 ( .A1(n4675), .A2(n6395), .B1(n959), .B2(n265), .ZN(n4126) );
  OAI22_X1 U1954 ( .A1(n4676), .A2(n264), .B1(n960), .B2(n265), .ZN(n4127) );
  NOR3_X1 U1956 ( .A1(\UUT/regfile/N457 ), .A2(net54931), .A3(n965), .ZN(n264)
         );
  OAI22_X1 U1957 ( .A1(n4742), .A2(n6392), .B1(n958), .B2(n259), .ZN(n4128) );
  OAI22_X1 U1958 ( .A1(n4748), .A2(n6392), .B1(n952), .B2(n259), .ZN(n4129) );
  OAI22_X1 U1959 ( .A1(n4771), .A2(n6392), .B1(n959), .B2(n259), .ZN(n4130) );
  OAI22_X1 U1960 ( .A1(n4772), .A2(n258), .B1(n960), .B2(n259), .ZN(n4131) );
  NOR3_X1 U1962 ( .A1(\UUT/regfile/N445 ), .A2(net54927), .A3(n966), .ZN(n258)
         );
  OAI22_X1 U1963 ( .A1(n4806), .A2(n6387), .B1(n958), .B2(n255), .ZN(n4132) );
  OAI22_X1 U1964 ( .A1(n4812), .A2(n6387), .B1(n952), .B2(n255), .ZN(n4133) );
  OAI22_X1 U1965 ( .A1(n4835), .A2(n6387), .B1(n959), .B2(n255), .ZN(n4134) );
  OAI22_X1 U1966 ( .A1(n4836), .A2(n254), .B1(n960), .B2(n255), .ZN(n4135) );
  NOR3_X1 U1968 ( .A1(\UUT/regfile/N433 ), .A2(net54931), .A3(n965), .ZN(n254)
         );
  OAI22_X1 U1969 ( .A1(n4870), .A2(n6384), .B1(n958), .B2(n251), .ZN(n4136) );
  OAI22_X1 U1970 ( .A1(n4876), .A2(n6384), .B1(n952), .B2(n251), .ZN(n4137) );
  OAI22_X1 U1971 ( .A1(n4899), .A2(n6384), .B1(n959), .B2(n251), .ZN(n4138) );
  OAI22_X1 U1972 ( .A1(n4900), .A2(n250), .B1(n960), .B2(n251), .ZN(n4139) );
  NOR3_X1 U1974 ( .A1(\UUT/regfile/N421 ), .A2(net54929), .A3(n966), .ZN(n250)
         );
  OAI22_X1 U1975 ( .A1(n4934), .A2(n6382), .B1(n958), .B2(n247), .ZN(n4140) );
  OAI22_X1 U1976 ( .A1(n4940), .A2(n6382), .B1(n952), .B2(n247), .ZN(n4141) );
  OAI22_X1 U1977 ( .A1(n4963), .A2(n6382), .B1(n959), .B2(n247), .ZN(n4142) );
  OAI22_X1 U1978 ( .A1(n4964), .A2(n246), .B1(n960), .B2(n247), .ZN(n4143) );
  NOR3_X1 U1980 ( .A1(\UUT/regfile/N409 ), .A2(net54931), .A3(n965), .ZN(n246)
         );
  OAI22_X1 U1981 ( .A1(n4998), .A2(n6385), .B1(n958), .B2(n243), .ZN(n4144) );
  OAI22_X1 U1982 ( .A1(n5004), .A2(n6385), .B1(n952), .B2(n243), .ZN(n4145) );
  OAI22_X1 U1983 ( .A1(n5027), .A2(n6385), .B1(n959), .B2(n243), .ZN(n4146) );
  OAI22_X1 U1984 ( .A1(n5028), .A2(n242), .B1(n960), .B2(n243), .ZN(n4147) );
  NOR3_X1 U1986 ( .A1(\UUT/regfile/N397 ), .A2(net54929), .A3(n966), .ZN(n242)
         );
  OAI22_X1 U1987 ( .A1(n5094), .A2(n6391), .B1(n958), .B2(n237), .ZN(n4148) );
  OAI22_X1 U1988 ( .A1(n5100), .A2(n6391), .B1(n952), .B2(n237), .ZN(n4149) );
  OAI22_X1 U1989 ( .A1(n5123), .A2(n6391), .B1(n959), .B2(n237), .ZN(n4150) );
  OAI22_X1 U1990 ( .A1(n5124), .A2(n236), .B1(n960), .B2(n237), .ZN(n4151) );
  NOR3_X1 U1992 ( .A1(\UUT/regfile/N385 ), .A2(net54929), .A3(n965), .ZN(n236)
         );
  OAI22_X1 U1993 ( .A1(n5158), .A2(n6396), .B1(n958), .B2(n233), .ZN(n4152) );
  OAI22_X1 U1994 ( .A1(n5164), .A2(n6396), .B1(n952), .B2(n233), .ZN(n4153) );
  OAI22_X1 U1995 ( .A1(n5187), .A2(n6396), .B1(n959), .B2(n233), .ZN(n4154) );
  OAI22_X1 U1996 ( .A1(n5188), .A2(n232), .B1(n960), .B2(n233), .ZN(n4155) );
  NOR3_X1 U1998 ( .A1(\UUT/regfile/N373 ), .A2(net54929), .A3(n966), .ZN(n232)
         );
  OAI22_X1 U1999 ( .A1(n5222), .A2(n6404), .B1(n958), .B2(n229), .ZN(n4156) );
  OAI22_X1 U2000 ( .A1(n5228), .A2(n6404), .B1(n952), .B2(n229), .ZN(n4157) );
  OAI22_X1 U2001 ( .A1(n5251), .A2(n6404), .B1(n959), .B2(n229), .ZN(n4158) );
  OAI22_X1 U2002 ( .A1(n5252), .A2(n228), .B1(n960), .B2(n229), .ZN(n4159) );
  NOR3_X1 U2004 ( .A1(\UUT/regfile/N360 ), .A2(net54931), .A3(n965), .ZN(n228)
         );
  OAI22_X1 U2005 ( .A1(n5286), .A2(n6406), .B1(n958), .B2(n225), .ZN(n4160) );
  OAI22_X1 U2006 ( .A1(n5292), .A2(n6406), .B1(n952), .B2(n225), .ZN(n4161) );
  OAI22_X1 U2007 ( .A1(n5315), .A2(n6406), .B1(n959), .B2(n225), .ZN(n4162) );
  OAI22_X1 U2008 ( .A1(n5316), .A2(n224), .B1(n960), .B2(n225), .ZN(n4163) );
  NOR3_X1 U2010 ( .A1(\UUT/regfile/N348 ), .A2(net54927), .A3(n966), .ZN(n224)
         );
  OAI22_X1 U2011 ( .A1(n5350), .A2(n6410), .B1(n958), .B2(n221), .ZN(n4164) );
  OAI22_X1 U2012 ( .A1(n5356), .A2(n6410), .B1(n952), .B2(n221), .ZN(n4165) );
  OAI22_X1 U2013 ( .A1(n5379), .A2(n6410), .B1(n959), .B2(n221), .ZN(n4166) );
  OAI22_X1 U2014 ( .A1(n5380), .A2(n220), .B1(n960), .B2(n221), .ZN(n4167) );
  NOR3_X1 U2016 ( .A1(\UUT/regfile/N336 ), .A2(net54931), .A3(n965), .ZN(n220)
         );
  OAI22_X1 U2017 ( .A1(n4422), .A2(n6411), .B1(n958), .B2(n279), .ZN(n4168) );
  OAI22_X1 U2018 ( .A1(n4428), .A2(n6411), .B1(n952), .B2(n279), .ZN(n4169) );
  OAI22_X1 U2019 ( .A1(n4451), .A2(n6411), .B1(n959), .B2(n279), .ZN(n4170) );
  OAI22_X1 U2020 ( .A1(n4452), .A2(n278), .B1(n960), .B2(n279), .ZN(n4171) );
  NOR3_X1 U2022 ( .A1(\UUT/regfile/N324 ), .A2(net54929), .A3(n966), .ZN(n278)
         );
  OAI22_X1 U2023 ( .A1(n4486), .A2(n6408), .B1(n958), .B2(n275), .ZN(n4172) );
  OAI22_X1 U2024 ( .A1(n4492), .A2(n6408), .B1(n952), .B2(n275), .ZN(n4173) );
  OAI22_X1 U2025 ( .A1(n4515), .A2(n6408), .B1(n959), .B2(n275), .ZN(n4174) );
  OAI22_X1 U2026 ( .A1(n4516), .A2(n274), .B1(n960), .B2(n275), .ZN(n4175) );
  NOR3_X1 U2028 ( .A1(\UUT/regfile/N311 ), .A2(net54929), .A3(n965), .ZN(n274)
         );
  OAI22_X1 U2029 ( .A1(n4550), .A2(n6397), .B1(n958), .B2(n271), .ZN(n4176) );
  OAI22_X1 U2030 ( .A1(n4556), .A2(n6397), .B1(n952), .B2(n271), .ZN(n4177) );
  OAI22_X1 U2031 ( .A1(n4579), .A2(n6397), .B1(n959), .B2(n271), .ZN(n4178) );
  OAI22_X1 U2032 ( .A1(n4580), .A2(n270), .B1(n960), .B2(n271), .ZN(n4179) );
  NOR3_X1 U2034 ( .A1(\UUT/regfile/N299 ), .A2(net54931), .A3(n966), .ZN(n270)
         );
  OAI22_X1 U2035 ( .A1(n4614), .A2(n6400), .B1(n958), .B2(n267), .ZN(n4180) );
  OAI22_X1 U2036 ( .A1(n4620), .A2(n6400), .B1(n952), .B2(n267), .ZN(n4181) );
  OAI22_X1 U2037 ( .A1(n4643), .A2(n6400), .B1(n959), .B2(n267), .ZN(n4182) );
  OAI22_X1 U2038 ( .A1(n4644), .A2(n266), .B1(n960), .B2(n267), .ZN(n4183) );
  NOR3_X1 U2040 ( .A1(\UUT/regfile/N286 ), .A2(net54931), .A3(n965), .ZN(n266)
         );
  NAND2_X1 U2041 ( .A1(n967), .A2(\UUT/rd_addr [1]), .ZN(n965) );
  OAI22_X1 U2042 ( .A1(n5062), .A2(n6390), .B1(n958), .B2(n239), .ZN(n4184) );
  OAI22_X1 U2043 ( .A1(n5068), .A2(n6390), .B1(n952), .B2(n239), .ZN(n4185) );
  OAI22_X1 U2044 ( .A1(n5091), .A2(n6390), .B1(n959), .B2(n239), .ZN(n4186) );
  OAI22_X1 U2045 ( .A1(n5092), .A2(n238), .B1(n960), .B2(n239), .ZN(n4187) );
  NOR3_X1 U2047 ( .A1(\UUT/regfile/N273 ), .A2(net54931), .A3(n966), .ZN(n238)
         );
  NAND2_X1 U2048 ( .A1(n967), .A2(n963), .ZN(n966) );
  INV_X1 U2049 ( .A(\UUT/rd_addr [1]), .ZN(n963) );
  INV_X1 U2050 ( .A(n964), .ZN(n967) );
  NAND2_X1 U2051 ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), .A2(n5413), .ZN(n964)
         );
  OAI221_X1 U2052 ( .B1(n140), .B2(n968), .C1(n5676), .C2(n142), .A(n969), 
        .ZN(n4188) );
  AOI22_X1 U2053 ( .A1(n144), .A2(n970), .B1(\UUT/Mpath/the_mult/Mad_out [0]), 
        .B2(n145), .ZN(n969) );
  NOR2_X1 U2055 ( .A1(n973), .A2(n974), .ZN(n972) );
  INV_X1 U2057 ( .A(\UUT/Mpath/the_mult/N255 ), .ZN(n973) );
  NAND3_X1 U2059 ( .A1(n971), .A2(n974), .A3(\UUT/Mpath/the_mult/N255 ), .ZN(
        n976) );
  INV_X1 U2060 ( .A(\UUT/Mpath/the_mult/N312 ), .ZN(n974) );
  INV_X1 U2061 ( .A(\UUT/Mpath/the_mult/N311 ), .ZN(n971) );
  OAI22_X1 U2063 ( .A1(net54909), .A2(n977), .B1(n5413), .B2(net54871), .ZN(
        n4189) );
  OAI22_X1 U2064 ( .A1(net54909), .A2(n978), .B1(net54863), .B2(n977), .ZN(
        n4190) );
  OAI22_X1 U2065 ( .A1(n6643), .A2(n546), .B1(n295), .B2(n2732), .ZN(n4191) );
  OAI22_X1 U2066 ( .A1(net54909), .A2(n980), .B1(net54863), .B2(n981), .ZN(
        n4192) );
  INV_X1 U2067 ( .A(\UUT/Mcontrol/m_sampled_xrd[0] ), .ZN(n981) );
  OAI221_X1 U2068 ( .B1(n6037), .B2(n982), .C1(net54889), .C2(n980), .A(n983), 
        .ZN(n4193) );
  AOI221_X1 U2069 ( .B1(n984), .B2(\UUT/Mcontrol/d_sampled_finstr [11]), .C1(
        n985), .C2(\UUT/Mcontrol/d_sampled_finstr [16]), .A(n986), .ZN(n983)
         );
  INV_X1 U2070 ( .A(\UUT/Mcontrol/x_rd[0] ), .ZN(n980) );
  OAI22_X1 U2071 ( .A1(net54909), .A2(n987), .B1(net54863), .B2(n2735), .ZN(
        n4194) );
  OAI221_X1 U2072 ( .B1(n5896), .B2(n982), .C1(net54891), .C2(n987), .A(n988), 
        .ZN(n4195) );
  AOI221_X1 U2073 ( .B1(n984), .B2(\UUT/Mcontrol/d_sampled_finstr [12]), .C1(
        n985), .C2(\UUT/Mcontrol/d_sampled_finstr [17]), .A(n986), .ZN(n988)
         );
  INV_X1 U2074 ( .A(\UUT/Mcontrol/x_rd[1] ), .ZN(n987) );
  OAI22_X1 U2075 ( .A1(net54911), .A2(n989), .B1(net54863), .B2(n2737), .ZN(
        n4196) );
  OAI221_X1 U2076 ( .B1(n5888), .B2(n982), .C1(net54889), .C2(n989), .A(n990), 
        .ZN(n4197) );
  AOI221_X1 U2077 ( .B1(n984), .B2(\UUT/Mcontrol/d_sampled_finstr [13]), .C1(
        n985), .C2(\UUT/Mcontrol/d_sampled_finstr [18]), .A(n986), .ZN(n990)
         );
  INV_X1 U2078 ( .A(\UUT/Mcontrol/x_rd[2] ), .ZN(n989) );
  OAI22_X1 U2079 ( .A1(net54911), .A2(n991), .B1(net54863), .B2(n2739), .ZN(
        n4198) );
  OAI221_X1 U2080 ( .B1(n5879), .B2(n982), .C1(net54889), .C2(n991), .A(n992), 
        .ZN(n4199) );
  AOI221_X1 U2081 ( .B1(n984), .B2(\UUT/Mcontrol/d_sampled_finstr [14]), .C1(
        n985), .C2(\UUT/Mcontrol/d_sampled_finstr [19]), .A(n986), .ZN(n992)
         );
  INV_X1 U2082 ( .A(\UUT/Mcontrol/x_rd[3] ), .ZN(n991) );
  OAI22_X1 U2083 ( .A1(net54911), .A2(n993), .B1(net54861), .B2(n2741), .ZN(
        n4200) );
  OAI221_X1 U2084 ( .B1(n5871), .B2(n982), .C1(net54889), .C2(n993), .A(n994), 
        .ZN(n4201) );
  AOI221_X1 U2085 ( .B1(n984), .B2(\UUT/Mcontrol/d_sampled_finstr [15]), .C1(
        n985), .C2(\UUT/Mcontrol/d_sampled_finstr [20]), .A(n986), .ZN(n994)
         );
  NOR4_X1 U2086 ( .A1(n995), .A2(n6039), .A3(n6038), .A4(
        \UUT/Mcontrol/Operation_decoding32/N1970 ), .ZN(n986) );
  AND2_X1 U2087 ( .A1(n996), .A2(net54895), .ZN(n985) );
  OAI21_X1 U2088 ( .B1(n997), .B2(n998), .A(n999), .ZN(n996) );
  INV_X1 U2089 ( .A(n1000), .ZN(n999) );
  AOI21_X1 U2090 ( .B1(n929), .B2(n6075), .A(n933), .ZN(n1000) );
  AOI221_X1 U2091 ( .B1(n1001), .B2(n931), .C1(n1002), .C2(n1003), .A(n1004), 
        .ZN(n997) );
  NAND3_X1 U2092 ( .A1(n6041), .A2(n6042), .A3(n6043), .ZN(n1003) );
  NAND2_X1 U2093 ( .A1(n6051), .A2(n857), .ZN(n1001) );
  AOI21_X1 U2094 ( .B1(n1005), .B2(n6030), .A(net54933), .ZN(n984) );
  OR3_X1 U2095 ( .A1(n998), .A2(n931), .A3(n1004), .ZN(n1005) );
  INV_X1 U2096 ( .A(\UUT/Mcontrol/x_rd[4] ), .ZN(n993) );
  NAND3_X1 U2097 ( .A1(n6044), .A2(n1006), .A3(n1007), .ZN(n982) );
  NOR3_X1 U2098 ( .A1(n1008), .A2(n6079), .A3(n6067), .ZN(n1007) );
  INV_X1 U2099 ( .A(n995), .ZN(n1006) );
  NAND3_X1 U2100 ( .A1(n921), .A2(net54869), .A3(n1002), .ZN(n995) );
  NOR3_X1 U2101 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2019 ), .A2(n6048), 
        .A3(n1004), .ZN(n1002) );
  INV_X1 U2102 ( .A(n998), .ZN(n921) );
  NAND3_X1 U2103 ( .A1(n929), .A2(n6030), .A3(n6075), .ZN(n998) );
  OAI22_X1 U2104 ( .A1(net54911), .A2(n1009), .B1(net54861), .B2(
        \UUT/Mpath/the_mult/N231 ), .ZN(n4202) );
  OAI22_X1 U2105 ( .A1(net54911), .A2(n1010), .B1(net54861), .B2(n1009), .ZN(
        n4203) );
  INV_X1 U2106 ( .A(\UUT/Mpath/the_mult/x_mul_command[0] ), .ZN(n1009) );
  OAI22_X1 U2107 ( .A1(n546), .A2(n1011), .B1(n5428), .B2(n295), .ZN(n4204) );
  INV_X1 U2108 ( .A(I_DATA_INBUS[0]), .ZN(n1011) );
  OAI22_X1 U2109 ( .A1(net54911), .A2(n1012), .B1(net54861), .B2(
        \UUT/Mpath/the_mult/N230 ), .ZN(n4205) );
  OAI22_X1 U2110 ( .A1(net54911), .A2(n1013), .B1(net54861), .B2(n1012), .ZN(
        n4206) );
  INV_X1 U2111 ( .A(\UUT/Mpath/the_mult/x_mul_command[1] ), .ZN(n1012) );
  OAI22_X1 U2112 ( .A1(net54911), .A2(n1013), .B1(net54861), .B2(
        \UUT/Mcontrol/st_logic/N27 ), .ZN(n4207) );
  INV_X1 U2113 ( .A(\UUT/d_mul_command [1]), .ZN(n1013) );
  OAI22_X1 U2114 ( .A1(n546), .A2(n1014), .B1(n5427), .B2(n295), .ZN(n4208) );
  INV_X1 U2115 ( .A(I_DATA_INBUS[1]), .ZN(n1014) );
  OAI22_X1 U2116 ( .A1(net54911), .A2(n1015), .B1(net54861), .B2(
        \UUT/Mpath/the_mult/N244 ), .ZN(n4209) );
  OAI22_X1 U2117 ( .A1(net54911), .A2(n1016), .B1(net54861), .B2(n1015), .ZN(
        n4210) );
  INV_X1 U2118 ( .A(\UUT/Mpath/the_mult/x_mul_command[2] ), .ZN(n1015) );
  OAI22_X1 U2119 ( .A1(net54911), .A2(n1016), .B1(net54861), .B2(
        \UUT/Mcontrol/st_logic/N26 ), .ZN(n4211) );
  INV_X1 U2120 ( .A(\UUT/d_mul_command [2]), .ZN(n1016) );
  OAI22_X1 U2121 ( .A1(n546), .A2(n1017), .B1(n5426), .B2(n295), .ZN(n4212) );
  INV_X1 U2122 ( .A(I_DATA_INBUS[2]), .ZN(n1017) );
  OAI22_X1 U2123 ( .A1(net54913), .A2(n1018), .B1(net54861), .B2(
        \UUT/Mpath/the_mult/N229 ), .ZN(n4213) );
  OAI22_X1 U2124 ( .A1(net54913), .A2(n1019), .B1(net54861), .B2(n1018), .ZN(
        n4214) );
  INV_X1 U2125 ( .A(\UUT/Mpath/the_mult/x_mul_command[3] ), .ZN(n1018) );
  OAI22_X1 U2126 ( .A1(net54913), .A2(n1019), .B1(net54859), .B2(n2748), .ZN(
        n4215) );
  INV_X1 U2127 ( .A(\UUT/d_mul_command [3]), .ZN(n1019) );
  OAI22_X1 U2128 ( .A1(n546), .A2(n1020), .B1(n5425), .B2(n295), .ZN(n4216) );
  INV_X1 U2129 ( .A(I_DATA_INBUS[3]), .ZN(n1020) );
  OAI22_X1 U2130 ( .A1(net54913), .A2(n1021), .B1(net54863), .B2(n2750), .ZN(
        n4217) );
  OAI22_X1 U2131 ( .A1(net54913), .A2(n1022), .B1(net54859), .B2(n1021), .ZN(
        n4218) );
  INV_X1 U2132 ( .A(\UUT/Mpath/the_mult/x_mul_command[4] ), .ZN(n1021) );
  OAI22_X1 U2133 ( .A1(net54913), .A2(n1022), .B1(net54859), .B2(n2752), .ZN(
        n4219) );
  OAI22_X1 U2134 ( .A1(n546), .A2(n1023), .B1(n5424), .B2(n295), .ZN(n4220) );
  INV_X1 U2135 ( .A(I_DATA_INBUS[4]), .ZN(n1023) );
  OAI22_X1 U2136 ( .A1(net54913), .A2(n1024), .B1(net54859), .B2(n2754), .ZN(
        n4221) );
  OAI22_X1 U2137 ( .A1(net54913), .A2(n1025), .B1(net54861), .B2(n1024), .ZN(
        n4222) );
  INV_X1 U2138 ( .A(\UUT/Mpath/the_mult/x_mul_command[5] ), .ZN(n1024) );
  OAI22_X1 U2139 ( .A1(net54913), .A2(n1025), .B1(net54859), .B2(n2756), .ZN(
        n4223) );
  OAI22_X1 U2140 ( .A1(n546), .A2(n1026), .B1(n5423), .B2(n295), .ZN(n4224) );
  INV_X1 U2141 ( .A(I_DATA_INBUS[5]), .ZN(n1026) );
  OAI22_X1 U2142 ( .A1(n546), .A2(n1027), .B1(n6143), .B2(n295), .ZN(n4225) );
  INV_X1 U2143 ( .A(I_DATA_INBUS[6]), .ZN(n1027) );
  OAI22_X1 U2144 ( .A1(n546), .A2(n1028), .B1(n6094), .B2(n295), .ZN(n4226) );
  INV_X1 U2145 ( .A(I_DATA_INBUS[7]), .ZN(n1028) );
  OAI22_X1 U2146 ( .A1(n546), .A2(n1029), .B1(n5897), .B2(n295), .ZN(n4227) );
  INV_X1 U2147 ( .A(I_DATA_INBUS[8]), .ZN(n1029) );
  OAI22_X1 U2148 ( .A1(n546), .A2(n1030), .B1(n5889), .B2(n295), .ZN(n4228) );
  INV_X1 U2149 ( .A(I_DATA_INBUS[9]), .ZN(n1030) );
  OAI22_X1 U2150 ( .A1(n546), .A2(n1031), .B1(n5881), .B2(n295), .ZN(n4229) );
  INV_X1 U2151 ( .A(I_DATA_INBUS[10]), .ZN(n1031) );
  OAI22_X1 U2152 ( .A1(n546), .A2(n1032), .B1(n6036), .B2(n295), .ZN(n4230) );
  INV_X1 U2153 ( .A(I_DATA_INBUS[11]), .ZN(n1032) );
  OAI22_X1 U2154 ( .A1(n546), .A2(n1033), .B1(n6035), .B2(n295), .ZN(n4231) );
  INV_X1 U2155 ( .A(I_DATA_INBUS[12]), .ZN(n1033) );
  OAI22_X1 U2156 ( .A1(n546), .A2(n1034), .B1(n6033), .B2(n295), .ZN(n4232) );
  INV_X1 U2157 ( .A(I_DATA_INBUS[13]), .ZN(n1034) );
  OAI22_X1 U2158 ( .A1(n546), .A2(n1035), .B1(n6032), .B2(n295), .ZN(n4233) );
  INV_X1 U2159 ( .A(I_DATA_INBUS[14]), .ZN(n1035) );
  OAI22_X1 U2160 ( .A1(n546), .A2(n1036), .B1(n5831), .B2(n295), .ZN(n4234) );
  INV_X1 U2161 ( .A(I_DATA_INBUS[15]), .ZN(n1036) );
  OAI22_X1 U2162 ( .A1(n546), .A2(n1037), .B1(n6027), .B2(n295), .ZN(n4235) );
  INV_X1 U2163 ( .A(I_DATA_INBUS[16]), .ZN(n1037) );
  OAI22_X1 U2164 ( .A1(n546), .A2(n1038), .B1(n6034), .B2(n295), .ZN(n4236) );
  INV_X1 U2165 ( .A(I_DATA_INBUS[17]), .ZN(n1038) );
  OAI22_X1 U2166 ( .A1(n546), .A2(n1039), .B1(n6026), .B2(n295), .ZN(n4237) );
  INV_X1 U2167 ( .A(I_DATA_INBUS[18]), .ZN(n1039) );
  OAI22_X1 U2168 ( .A1(n546), .A2(n1040), .B1(n6031), .B2(n295), .ZN(n4238) );
  INV_X1 U2169 ( .A(I_DATA_INBUS[19]), .ZN(n1040) );
  OAI22_X1 U2170 ( .A1(n546), .A2(n1041), .B1(n6029), .B2(n295), .ZN(n4239) );
  INV_X1 U2171 ( .A(I_DATA_INBUS[20]), .ZN(n1041) );
  OAI22_X1 U2172 ( .A1(n546), .A2(n1042), .B1(n6037), .B2(n295), .ZN(n4240) );
  INV_X1 U2173 ( .A(I_DATA_INBUS[21]), .ZN(n1042) );
  OAI22_X1 U2174 ( .A1(n546), .A2(n1043), .B1(n5896), .B2(n295), .ZN(n4241) );
  INV_X1 U2175 ( .A(I_DATA_INBUS[22]), .ZN(n1043) );
  OAI22_X1 U2176 ( .A1(n546), .A2(n1044), .B1(n5888), .B2(n295), .ZN(n4242) );
  INV_X1 U2177 ( .A(I_DATA_INBUS[23]), .ZN(n1044) );
  OAI22_X1 U2178 ( .A1(n546), .A2(n1045), .B1(n5879), .B2(n295), .ZN(n4243) );
  INV_X1 U2179 ( .A(I_DATA_INBUS[24]), .ZN(n1045) );
  OAI22_X1 U2180 ( .A1(n546), .A2(n1046), .B1(n5871), .B2(n295), .ZN(n4244) );
  INV_X1 U2181 ( .A(I_DATA_INBUS[25]), .ZN(n1046) );
  OAI21_X1 U2182 ( .B1(net54847), .B2(n1047), .A(n1048), .ZN(n4245) );
  OAI21_X1 U2183 ( .B1(n1049), .B2(n1050), .A(net54859), .ZN(n1048) );
  INV_X1 U2184 ( .A(n1051), .ZN(n1050) );
  NOR3_X1 U2185 ( .A1(n1052), .A2(\UUT/Mcontrol/Operation_decoding32/N2007 ), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N1995 ), .ZN(n1049) );
  OAI221_X1 U2186 ( .B1(net54931), .B2(n1053), .C1(net54891), .C2(n1054), .A(
        n1055), .ZN(n4246) );
  AOI21_X1 U2187 ( .B1(n1056), .B2(n6042), .A(
        \UUT/Mcontrol/Operation_decoding32/N2019 ), .ZN(n1053) );
  OAI21_X1 U2188 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2001 ), .B2(n1057), 
        .A(n1058), .ZN(n1056) );
  NOR3_X1 U2189 ( .A1(n1052), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N1995 ), .ZN(n1057) );
  INV_X1 U2190 ( .A(\UUT/Mcontrol/Operation_decoding32/N1987 ), .ZN(n1052) );
  OAI211_X1 U2191 ( .C1(net54877), .C2(n1059), .A(n1060), .B(n1055), .ZN(n4247) );
  NAND4_X1 U2192 ( .A1(n1061), .A2(net54869), .A3(n6042), .A4(
        \UUT/Mcontrol/Operation_decoding32/N1994 ), .ZN(n1060) );
  OAI22_X1 U2193 ( .A1(net54847), .A2(n2781), .B1(net54919), .B2(n116), .ZN(
        n4248) );
  AND4_X1 U2194 ( .A1(n1051), .A2(n1062), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1994 ), .A4(n1058), .ZN(n116) );
  INV_X1 U2195 ( .A(\UUT/Mcontrol/Operation_decoding32/N2007 ), .ZN(n1058) );
  NAND3_X1 U2196 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1987 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1981 ), .ZN(n1062) );
  NOR4_X1 U2197 ( .A1(n1063), .A2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
        .A3(n1064), .A4(\UUT/Mcontrol/Operation_decoding32/N2001 ), .ZN(n1051)
         );
  OAI221_X1 U2198 ( .B1(n1065), .B2(n1066), .C1(net54889), .C2(n1067), .A(
        n1055), .ZN(n4249) );
  NAND2_X1 U2199 ( .A1(net54877), .A2(n1063), .ZN(n1055) );
  INV_X1 U2200 ( .A(n6050), .ZN(n1063) );
  INV_X1 U2201 ( .A(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), .ZN(n1067)
         );
  NAND2_X1 U2202 ( .A1(net54875), .A2(n6042), .ZN(n1066) );
  AOI21_X1 U2203 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2017 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N2005 ), .A(
        \UUT/Mcontrol/d_instr [26]), .ZN(n1065) );
  OAI21_X1 U2204 ( .B1(n295), .B2(n2783), .A(n1068), .ZN(n4250) );
  NAND2_X1 U2205 ( .A1(I_DATA_INBUS[26]), .A2(n295), .ZN(n1068) );
  OAI21_X1 U2206 ( .B1(n295), .B2(n2784), .A(n1069), .ZN(n4251) );
  NAND2_X1 U2207 ( .A1(I_DATA_INBUS[27]), .A2(n295), .ZN(n1069) );
  OAI21_X1 U2208 ( .B1(n295), .B2(n2785), .A(n1070), .ZN(n4252) );
  NAND2_X1 U2209 ( .A1(I_DATA_INBUS[28]), .A2(n295), .ZN(n1070) );
  OAI22_X1 U2210 ( .A1(n546), .A2(n1071), .B1(n6071), .B2(n295), .ZN(n4253) );
  INV_X1 U2211 ( .A(I_DATA_INBUS[29]), .ZN(n1071) );
  OAI22_X1 U2212 ( .A1(n546), .A2(n1072), .B1(n6070), .B2(n295), .ZN(n4254) );
  INV_X1 U2213 ( .A(I_DATA_INBUS[30]), .ZN(n1072) );
  OAI22_X1 U2214 ( .A1(net54917), .A2(n1010), .B1(net54863), .B2(
        \UUT/Mcontrol/st_logic/N34 ), .ZN(n4255) );
  INV_X1 U2215 ( .A(\UUT/d_mul_command [0]), .ZN(n1010) );
  OAI221_X1 U2216 ( .B1(n1073), .B2(n316), .C1(\UUT/Mpath/the_alu/N83 ), .C2(
        net54889), .A(n1074), .ZN(n4256) );
  AOI22_X1 U2217 ( .A1(n318), .A2(n1075), .B1(n319), .B2(n1076), .ZN(n1074) );
  NAND2_X1 U2220 ( .A1(net54875), .A2(n1077), .ZN(n316) );
  OAI22_X1 U2221 ( .A1(net54917), .A2(n1078), .B1(net54863), .B2(n968), .ZN(
        n4257) );
  INV_X1 U2222 ( .A(n6869), .ZN(n968) );
  INV_X1 U2223 ( .A(\UUT/Mpath/the_mult/x_mult_out[0] ), .ZN(n1078) );
  OAI22_X1 U2224 ( .A1(net54915), .A2(n1079), .B1(net54863), .B2(n794), .ZN(
        n4258) );
  INV_X1 U2225 ( .A(n6517), .ZN(n794) );
  INV_X1 U2226 ( .A(\UUT/Mpath/the_mult/x_mult_out[1] ), .ZN(n1079) );
  OAI22_X1 U2227 ( .A1(net54915), .A2(n1080), .B1(net54863), .B2(n772), .ZN(
        n4259) );
  INV_X1 U2228 ( .A(n6518), .ZN(n772) );
  INV_X1 U2229 ( .A(\UUT/Mpath/the_mult/x_mult_out[2] ), .ZN(n1080) );
  OAI22_X1 U2230 ( .A1(net54917), .A2(n1081), .B1(net54867), .B2(n749), .ZN(
        n4260) );
  INV_X1 U2231 ( .A(\UUT/Mpath/the_mult/Mult_out[3] ), .ZN(n749) );
  INV_X1 U2232 ( .A(\UUT/Mpath/the_mult/x_mult_out[3] ), .ZN(n1081) );
  OAI22_X1 U2233 ( .A1(net54917), .A2(n1082), .B1(net54863), .B2(n726), .ZN(
        n4261) );
  INV_X1 U2234 ( .A(\UUT/Mpath/the_mult/Mult_out[4] ), .ZN(n726) );
  INV_X1 U2235 ( .A(\UUT/Mpath/the_mult/x_mult_out[4] ), .ZN(n1082) );
  OAI22_X1 U2236 ( .A1(net54917), .A2(n1083), .B1(net54865), .B2(n703), .ZN(
        n4262) );
  INV_X1 U2237 ( .A(\UUT/Mpath/the_mult/Mult_out[5] ), .ZN(n703) );
  INV_X1 U2238 ( .A(\UUT/Mpath/the_mult/x_mult_out[5] ), .ZN(n1083) );
  OAI22_X1 U2239 ( .A1(net54919), .A2(n1084), .B1(net54863), .B2(n675), .ZN(
        n4263) );
  INV_X1 U2240 ( .A(\UUT/Mpath/the_mult/Mult_out[6] ), .ZN(n675) );
  INV_X1 U2241 ( .A(\UUT/Mpath/the_mult/x_mult_out[6] ), .ZN(n1084) );
  OAI22_X1 U2242 ( .A1(net54917), .A2(n1085), .B1(net54865), .B2(n652), .ZN(
        n4264) );
  INV_X1 U2243 ( .A(\UUT/Mpath/the_mult/Mult_out[7] ), .ZN(n652) );
  INV_X1 U2244 ( .A(\UUT/Mpath/the_mult/x_mult_out[7] ), .ZN(n1085) );
  OAI22_X1 U2245 ( .A1(net54917), .A2(n1086), .B1(net54865), .B2(n635), .ZN(
        n4265) );
  INV_X1 U2246 ( .A(\UUT/Mpath/the_mult/Mult_out[8] ), .ZN(n635) );
  INV_X1 U2247 ( .A(\UUT/Mpath/the_mult/x_mult_out[8] ), .ZN(n1086) );
  OAI22_X1 U2248 ( .A1(net54913), .A2(n1087), .B1(net54865), .B2(n615), .ZN(
        n4266) );
  INV_X1 U2249 ( .A(\UUT/Mpath/the_mult/Mult_out[9] ), .ZN(n615) );
  INV_X1 U2250 ( .A(\UUT/Mpath/the_mult/x_mult_out[9] ), .ZN(n1087) );
  OAI22_X1 U2251 ( .A1(net54919), .A2(n1088), .B1(net54865), .B2(n599), .ZN(
        n4267) );
  INV_X1 U2252 ( .A(\UUT/Mpath/the_mult/Mult_out[10] ), .ZN(n599) );
  INV_X1 U2253 ( .A(\UUT/Mpath/the_mult/x_mult_out[10] ), .ZN(n1088) );
  OAI22_X1 U2254 ( .A1(net54919), .A2(n1089), .B1(net54865), .B2(n580), .ZN(
        n4268) );
  INV_X1 U2255 ( .A(\UUT/Mpath/the_mult/Mult_out[11] ), .ZN(n580) );
  INV_X1 U2256 ( .A(\UUT/Mpath/the_mult/x_mult_out[11] ), .ZN(n1089) );
  OAI22_X1 U2257 ( .A1(net54919), .A2(n1090), .B1(net54865), .B2(n555), .ZN(
        n4269) );
  INV_X1 U2258 ( .A(\UUT/Mpath/the_mult/Mult_out[12] ), .ZN(n555) );
  INV_X1 U2259 ( .A(\UUT/Mpath/the_mult/x_mult_out[12] ), .ZN(n1090) );
  OAI22_X1 U2260 ( .A1(net54919), .A2(n1091), .B1(net54865), .B2(n529), .ZN(
        n4270) );
  INV_X1 U2261 ( .A(\UUT/Mpath/the_mult/Mult_out[13] ), .ZN(n529) );
  INV_X1 U2262 ( .A(\UUT/Mpath/the_mult/x_mult_out[13] ), .ZN(n1091) );
  OAI22_X1 U2263 ( .A1(net54919), .A2(n1092), .B1(net54865), .B2(n504), .ZN(
        n4271) );
  INV_X1 U2264 ( .A(\UUT/Mpath/the_mult/Mult_out[14] ), .ZN(n504) );
  INV_X1 U2265 ( .A(\UUT/Mpath/the_mult/x_mult_out[14] ), .ZN(n1092) );
  OAI22_X1 U2266 ( .A1(net54917), .A2(n1093), .B1(net54865), .B2(n475), .ZN(
        n4272) );
  INV_X1 U2267 ( .A(\UUT/Mpath/the_mult/Mult_out[15] ), .ZN(n475) );
  INV_X1 U2268 ( .A(\UUT/Mpath/the_mult/x_mult_out[15] ), .ZN(n1093) );
  OAI22_X1 U2269 ( .A1(net54917), .A2(n1094), .B1(net54867), .B2(n454), .ZN(
        n4273) );
  INV_X1 U2270 ( .A(\UUT/Mpath/the_mult/Mult_out[16] ), .ZN(n454) );
  INV_X1 U2271 ( .A(\UUT/Mpath/the_mult/x_mult_out[16] ), .ZN(n1094) );
  OAI22_X1 U2272 ( .A1(net54919), .A2(n1095), .B1(net54867), .B2(n427), .ZN(
        n4274) );
  INV_X1 U2273 ( .A(\UUT/Mpath/the_mult/Mult_out[17] ), .ZN(n427) );
  INV_X1 U2274 ( .A(\UUT/Mpath/the_mult/x_mult_out[17] ), .ZN(n1095) );
  OAI22_X1 U2275 ( .A1(net54915), .A2(n1096), .B1(net54867), .B2(n405), .ZN(
        n4275) );
  INV_X1 U2276 ( .A(\UUT/Mpath/the_mult/Mult_out[18] ), .ZN(n405) );
  INV_X1 U2277 ( .A(\UUT/Mpath/the_mult/x_mult_out[18] ), .ZN(n1096) );
  OAI22_X1 U2278 ( .A1(net54917), .A2(n1097), .B1(net54867), .B2(n383), .ZN(
        n4276) );
  INV_X1 U2279 ( .A(\UUT/Mpath/the_mult/Mult_out[19] ), .ZN(n383) );
  INV_X1 U2280 ( .A(\UUT/Mpath/the_mult/x_mult_out[19] ), .ZN(n1097) );
  OAI22_X1 U2281 ( .A1(net54917), .A2(n1098), .B1(net54867), .B2(n357), .ZN(
        n4277) );
  INV_X1 U2282 ( .A(\UUT/Mpath/the_mult/Mult_out[20] ), .ZN(n357) );
  INV_X1 U2283 ( .A(\UUT/Mpath/the_mult/x_mult_out[20] ), .ZN(n1098) );
  OAI22_X1 U2284 ( .A1(net54915), .A2(n1099), .B1(net54867), .B2(n336), .ZN(
        n4278) );
  INV_X1 U2285 ( .A(\UUT/Mpath/the_mult/Mult_out[21] ), .ZN(n336) );
  INV_X1 U2286 ( .A(\UUT/Mpath/the_mult/x_mult_out[21] ), .ZN(n1099) );
  OAI22_X1 U2287 ( .A1(net54917), .A2(n1100), .B1(net54867), .B2(n307), .ZN(
        n4279) );
  INV_X1 U2288 ( .A(\UUT/Mpath/the_mult/Mult_out[22] ), .ZN(n307) );
  INV_X1 U2289 ( .A(\UUT/Mpath/the_mult/x_mult_out[22] ), .ZN(n1100) );
  OAI22_X1 U2290 ( .A1(net54915), .A2(n1101), .B1(net54867), .B2(n806), .ZN(
        n4280) );
  INV_X1 U2291 ( .A(\UUT/Mpath/the_mult/Mult_out[23] ), .ZN(n806) );
  INV_X1 U2292 ( .A(\UUT/Mpath/the_mult/x_mult_out[23] ), .ZN(n1101) );
  OAI22_X1 U2293 ( .A1(net54915), .A2(n1102), .B1(net54867), .B2(n213), .ZN(
        n4281) );
  INV_X1 U2294 ( .A(\UUT/Mpath/the_mult/Mult_out[24] ), .ZN(n213) );
  INV_X1 U2295 ( .A(\UUT/Mpath/the_mult/x_mult_out[24] ), .ZN(n1102) );
  OAI22_X1 U2296 ( .A1(net54915), .A2(n1103), .B1(net54867), .B2(n198), .ZN(
        n4282) );
  INV_X1 U2297 ( .A(\UUT/Mpath/the_mult/Mult_out[25] ), .ZN(n198) );
  INV_X1 U2298 ( .A(\UUT/Mpath/the_mult/x_mult_out[25] ), .ZN(n1103) );
  OAI22_X1 U2299 ( .A1(net54915), .A2(n1104), .B1(net54869), .B2(n185), .ZN(
        n4283) );
  INV_X1 U2300 ( .A(\UUT/Mpath/the_mult/Mult_out[26] ), .ZN(n185) );
  INV_X1 U2301 ( .A(\UUT/Mpath/the_mult/x_mult_out[26] ), .ZN(n1104) );
  OAI22_X1 U2302 ( .A1(net54915), .A2(n1105), .B1(net54869), .B2(n169), .ZN(
        n4284) );
  INV_X1 U2303 ( .A(\UUT/Mpath/the_mult/Mult_out[27] ), .ZN(n169) );
  INV_X1 U2304 ( .A(\UUT/Mpath/the_mult/x_mult_out[27] ), .ZN(n1105) );
  OAI22_X1 U2305 ( .A1(net54915), .A2(n1106), .B1(net54869), .B2(n157), .ZN(
        n4285) );
  INV_X1 U2306 ( .A(\UUT/Mpath/the_mult/Mult_out[28] ), .ZN(n157) );
  INV_X1 U2307 ( .A(\UUT/Mpath/the_mult/x_mult_out[28] ), .ZN(n1106) );
  OAI22_X1 U2308 ( .A1(net54913), .A2(n1107), .B1(net54869), .B2(n141), .ZN(
        n4286) );
  INV_X1 U2309 ( .A(\UUT/Mpath/the_mult/Mult_out[29] ), .ZN(n141) );
  INV_X1 U2310 ( .A(\UUT/Mpath/the_mult/x_mult_out[29] ), .ZN(n1107) );
  OAI22_X1 U2311 ( .A1(net54915), .A2(n1108), .B1(net54869), .B2(n864), .ZN(
        n4287) );
  INV_X1 U2312 ( .A(\UUT/Mpath/the_mult/Mult_out[30] ), .ZN(n864) );
  INV_X1 U2313 ( .A(\UUT/Mpath/the_mult/x_mult_out[30] ), .ZN(n1108) );
  OAI22_X1 U2314 ( .A1(net54915), .A2(n1109), .B1(net54869), .B2(n946), .ZN(
        n4288) );
  INV_X1 U2315 ( .A(\UUT/Mpath/the_mult/Mult_out[31] ), .ZN(n946) );
  INV_X1 U2316 ( .A(\UUT/Mpath/the_mult/x_mult_out[31] ), .ZN(n1109) );
  OAI21_X1 U2317 ( .B1(net54847), .B2(n1110), .A(n1111), .ZN(n4289) );
  NAND2_X1 U2318 ( .A1(\UUT/Mpath/the_mult/x_mult_out[32] ), .A2(net54855), 
        .ZN(n1111) );
  OAI21_X1 U2319 ( .B1(net54847), .B2(n791), .A(n1112), .ZN(n4290) );
  NAND2_X1 U2320 ( .A1(\UUT/Mpath/the_mult/x_mult_out[33] ), .A2(net54855), 
        .ZN(n1112) );
  INV_X1 U2321 ( .A(\UUT/Mpath/the_mult/Mult_out[33] ), .ZN(n791) );
  OAI21_X1 U2322 ( .B1(net54847), .B2(n769), .A(n1113), .ZN(n4291) );
  NAND2_X1 U2323 ( .A1(\UUT/Mpath/the_mult/x_mult_out[34] ), .A2(net54855), 
        .ZN(n1113) );
  INV_X1 U2324 ( .A(\UUT/Mpath/the_mult/Mult_out[34] ), .ZN(n769) );
  OAI21_X1 U2325 ( .B1(net54847), .B2(n746), .A(n1114), .ZN(n4292) );
  NAND2_X1 U2326 ( .A1(\UUT/Mpath/the_mult/x_mult_out[35] ), .A2(net54855), 
        .ZN(n1114) );
  INV_X1 U2327 ( .A(\UUT/Mpath/the_mult/Mult_out[35] ), .ZN(n746) );
  OAI21_X1 U2328 ( .B1(net54847), .B2(n723), .A(n1115), .ZN(n4293) );
  NAND2_X1 U2329 ( .A1(\UUT/Mpath/the_mult/x_mult_out[36] ), .A2(net54855), 
        .ZN(n1115) );
  INV_X1 U2330 ( .A(\UUT/Mpath/the_mult/Mult_out[36] ), .ZN(n723) );
  OAI21_X1 U2331 ( .B1(net54849), .B2(n700), .A(n1116), .ZN(n4294) );
  NAND2_X1 U2332 ( .A1(\UUT/Mpath/the_mult/x_mult_out[37] ), .A2(net54853), 
        .ZN(n1116) );
  INV_X1 U2333 ( .A(\UUT/Mpath/the_mult/Mult_out[37] ), .ZN(n700) );
  OAI21_X1 U2334 ( .B1(net54849), .B2(n672), .A(n1117), .ZN(n4295) );
  NAND2_X1 U2335 ( .A1(\UUT/Mpath/the_mult/x_mult_out[38] ), .A2(net54855), 
        .ZN(n1117) );
  INV_X1 U2336 ( .A(\UUT/Mpath/the_mult/Mult_out[38] ), .ZN(n672) );
  OAI21_X1 U2337 ( .B1(net54849), .B2(n649), .A(n1118), .ZN(n4296) );
  NAND2_X1 U2338 ( .A1(\UUT/Mpath/the_mult/x_mult_out[39] ), .A2(net54853), 
        .ZN(n1118) );
  INV_X1 U2339 ( .A(\UUT/Mpath/the_mult/Mult_out[39] ), .ZN(n649) );
  OAI21_X1 U2340 ( .B1(net54849), .B2(n632), .A(n1119), .ZN(n4297) );
  NAND2_X1 U2341 ( .A1(\UUT/Mpath/the_mult/x_mult_out[40] ), .A2(net54853), 
        .ZN(n1119) );
  INV_X1 U2342 ( .A(\UUT/Mpath/the_mult/Mult_out[40] ), .ZN(n632) );
  OAI21_X1 U2343 ( .B1(net54849), .B2(n612), .A(n1120), .ZN(n4298) );
  NAND2_X1 U2344 ( .A1(\UUT/Mpath/the_mult/x_mult_out[41] ), .A2(net54855), 
        .ZN(n1120) );
  INV_X1 U2345 ( .A(\UUT/Mpath/the_mult/Mult_out[41] ), .ZN(n612) );
  OAI21_X1 U2346 ( .B1(net54849), .B2(n596), .A(n1121), .ZN(n4299) );
  NAND2_X1 U2347 ( .A1(\UUT/Mpath/the_mult/x_mult_out[42] ), .A2(net54853), 
        .ZN(n1121) );
  INV_X1 U2348 ( .A(\UUT/Mpath/the_mult/Mult_out[42] ), .ZN(n596) );
  OAI21_X1 U2349 ( .B1(net54849), .B2(n577), .A(n1122), .ZN(n4300) );
  NAND2_X1 U2350 ( .A1(\UUT/Mpath/the_mult/x_mult_out[43] ), .A2(net54853), 
        .ZN(n1122) );
  INV_X1 U2351 ( .A(\UUT/Mpath/the_mult/Mult_out[43] ), .ZN(n577) );
  OAI21_X1 U2352 ( .B1(net54849), .B2(n552), .A(n1123), .ZN(n4301) );
  NAND2_X1 U2353 ( .A1(\UUT/Mpath/the_mult/x_mult_out[44] ), .A2(net54853), 
        .ZN(n1123) );
  INV_X1 U2354 ( .A(\UUT/Mpath/the_mult/Mult_out[44] ), .ZN(n552) );
  OAI21_X1 U2355 ( .B1(net54849), .B2(n526), .A(n1124), .ZN(n4302) );
  NAND2_X1 U2356 ( .A1(\UUT/Mpath/the_mult/x_mult_out[45] ), .A2(net54853), 
        .ZN(n1124) );
  INV_X1 U2357 ( .A(\UUT/Mpath/the_mult/Mult_out[45] ), .ZN(n526) );
  OAI21_X1 U2358 ( .B1(net54851), .B2(n501), .A(n1125), .ZN(n4303) );
  NAND2_X1 U2359 ( .A1(\UUT/Mpath/the_mult/x_mult_out[46] ), .A2(net54855), 
        .ZN(n1125) );
  INV_X1 U2360 ( .A(\UUT/Mpath/the_mult/Mult_out[46] ), .ZN(n501) );
  OAI21_X1 U2361 ( .B1(net54851), .B2(n472), .A(n1126), .ZN(n4304) );
  NAND2_X1 U2362 ( .A1(\UUT/Mpath/the_mult/x_mult_out[47] ), .A2(net54853), 
        .ZN(n1126) );
  INV_X1 U2363 ( .A(\UUT/Mpath/the_mult/Mult_out[47] ), .ZN(n472) );
  OAI21_X1 U2364 ( .B1(net54851), .B2(n451), .A(n1127), .ZN(n4305) );
  NAND2_X1 U2365 ( .A1(\UUT/Mpath/the_mult/x_mult_out[48] ), .A2(net54853), 
        .ZN(n1127) );
  INV_X1 U2366 ( .A(\UUT/Mpath/the_mult/Mult_out[48] ), .ZN(n451) );
  OAI21_X1 U2367 ( .B1(net54849), .B2(n424), .A(n1128), .ZN(n4306) );
  NAND2_X1 U2368 ( .A1(\UUT/Mpath/the_mult/x_mult_out[49] ), .A2(net54855), 
        .ZN(n1128) );
  INV_X1 U2369 ( .A(\UUT/Mpath/the_mult/Mult_out[49] ), .ZN(n424) );
  OAI21_X1 U2370 ( .B1(net54851), .B2(n402), .A(n1129), .ZN(n4307) );
  NAND2_X1 U2371 ( .A1(\UUT/Mpath/the_mult/x_mult_out[50] ), .A2(net54855), 
        .ZN(n1129) );
  INV_X1 U2372 ( .A(\UUT/Mpath/the_mult/Mult_out[50] ), .ZN(n402) );
  OAI21_X1 U2373 ( .B1(net54851), .B2(n380), .A(n1130), .ZN(n4308) );
  NAND2_X1 U2374 ( .A1(\UUT/Mpath/the_mult/x_mult_out[51] ), .A2(net54855), 
        .ZN(n1130) );
  INV_X1 U2375 ( .A(\UUT/Mpath/the_mult/Mult_out[51] ), .ZN(n380) );
  OAI21_X1 U2376 ( .B1(net54851), .B2(n354), .A(n1131), .ZN(n4309) );
  NAND2_X1 U2377 ( .A1(\UUT/Mpath/the_mult/x_mult_out[52] ), .A2(net54857), 
        .ZN(n1131) );
  INV_X1 U2378 ( .A(\UUT/Mpath/the_mult/Mult_out[52] ), .ZN(n354) );
  OAI21_X1 U2379 ( .B1(net54851), .B2(n333), .A(n1132), .ZN(n4310) );
  NAND2_X1 U2380 ( .A1(\UUT/Mpath/the_mult/x_mult_out[53] ), .A2(net54855), 
        .ZN(n1132) );
  INV_X1 U2381 ( .A(\UUT/Mpath/the_mult/Mult_out[53] ), .ZN(n333) );
  OAI21_X1 U2382 ( .B1(net54849), .B2(n304), .A(n1133), .ZN(n4311) );
  NAND2_X1 U2383 ( .A1(\UUT/Mpath/the_mult/x_mult_out[54] ), .A2(net54857), 
        .ZN(n1133) );
  INV_X1 U2384 ( .A(\UUT/Mpath/the_mult/Mult_out[54] ), .ZN(n304) );
  OAI21_X1 U2385 ( .B1(net54851), .B2(n803), .A(n1134), .ZN(n4312) );
  NAND2_X1 U2386 ( .A1(\UUT/Mpath/the_mult/x_mult_out[55] ), .A2(net54857), 
        .ZN(n1134) );
  INV_X1 U2387 ( .A(\UUT/Mpath/the_mult/Mult_out[55] ), .ZN(n803) );
  OAI21_X1 U2388 ( .B1(net54851), .B2(n210), .A(n1135), .ZN(n4313) );
  NAND2_X1 U2389 ( .A1(\UUT/Mpath/the_mult/x_mult_out[56] ), .A2(net54857), 
        .ZN(n1135) );
  INV_X1 U2390 ( .A(\UUT/Mpath/the_mult/Mult_out[56] ), .ZN(n210) );
  OAI21_X1 U2391 ( .B1(net54851), .B2(n195), .A(n1136), .ZN(n4314) );
  NAND2_X1 U2392 ( .A1(\UUT/Mpath/the_mult/x_mult_out[57] ), .A2(net54857), 
        .ZN(n1136) );
  INV_X1 U2393 ( .A(\UUT/Mpath/the_mult/Mult_out[57] ), .ZN(n195) );
  OAI21_X1 U2394 ( .B1(net54851), .B2(n182), .A(n1137), .ZN(n4315) );
  NAND2_X1 U2395 ( .A1(\UUT/Mpath/the_mult/x_mult_out[58] ), .A2(net54857), 
        .ZN(n1137) );
  INV_X1 U2396 ( .A(\UUT/Mpath/the_mult/Mult_out[58] ), .ZN(n182) );
  OAI21_X1 U2397 ( .B1(net54853), .B2(n166), .A(n1138), .ZN(n4316) );
  NAND2_X1 U2398 ( .A1(\UUT/Mpath/the_mult/x_mult_out[59] ), .A2(net54857), 
        .ZN(n1138) );
  INV_X1 U2399 ( .A(\UUT/Mpath/the_mult/Mult_out[59] ), .ZN(n166) );
  OAI21_X1 U2400 ( .B1(net54849), .B2(n154), .A(n1139), .ZN(n4317) );
  NAND2_X1 U2401 ( .A1(\UUT/Mpath/the_mult/x_mult_out[60] ), .A2(net54857), 
        .ZN(n1139) );
  INV_X1 U2402 ( .A(\UUT/Mpath/the_mult/Mult_out[60] ), .ZN(n154) );
  OAI21_X1 U2403 ( .B1(net54853), .B2(n134), .A(n1140), .ZN(n4318) );
  NAND2_X1 U2404 ( .A1(\UUT/Mpath/the_mult/x_mult_out[61] ), .A2(net54857), 
        .ZN(n1140) );
  INV_X1 U2405 ( .A(\UUT/Mpath/the_mult/Mult_out[61] ), .ZN(n134) );
  OAI21_X1 U2406 ( .B1(net54853), .B2(n861), .A(n1141), .ZN(n4319) );
  NAND2_X1 U2407 ( .A1(\UUT/Mpath/the_mult/x_mult_out[62] ), .A2(net54857), 
        .ZN(n1141) );
  INV_X1 U2408 ( .A(\UUT/Mpath/the_mult/Mult_out[62] ), .ZN(n861) );
  OAI21_X1 U2409 ( .B1(net54851), .B2(n1142), .A(n1143), .ZN(n4320) );
  NAND2_X1 U2410 ( .A1(\UUT/Mpath/the_mult/x_mult_out[63] ), .A2(net54857), 
        .ZN(n1143) );
  OAI22_X1 U2411 ( .A1(n5527), .A2(net54879), .B1(n1073), .B2(net54933), .ZN(
        n4321) );
  OAI22_X1 U2412 ( .A1(n1144), .A2(net54937), .B1(
        \UUT/Mpath/the_memhandle/N240 ), .B2(net54875), .ZN(n4322) );
  INV_X1 U2413 ( .A(\UUT/daddr_out [0]), .ZN(n1144) );
  OAI222_X1 U2414 ( .A1(n80), .A2(n123), .B1(n79), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N68 ), .C2(net54893), .ZN(n4324) );
  INV_X1 U2415 ( .A(\UUT/break_code[8] ), .ZN(n79) );
  INV_X1 U2416 ( .A(n1145), .ZN(n80) );
  OAI222_X1 U2417 ( .A1(n638), .A2(n129), .B1(n958), .B2(n131), .C1(n5436), 
        .C2(n132), .ZN(n1145) );
  OAI211_X1 U2419 ( .C1(n1146), .C2(n482), .A(n484), .B(n1147), .ZN(n641) );
  AOI22_X1 U2420 ( .A1(n486), .A2(n1148), .B1(n1149), .B2(n489), .ZN(n1147) );
  INV_X1 U2421 ( .A(n5437), .ZN(n1149) );
  INV_X1 U2422 ( .A(n5747), .ZN(n1146) );
  INV_X1 U2423 ( .A(n1150), .ZN(n638) );
  OAI211_X1 U2424 ( .C1(n5616), .C2(n321), .A(n1151), .B(n1152), .ZN(n1150) );
  AOI222_X1 U2425 ( .A1(n285), .A2(n1153), .B1(\UUT/Mpath/out_jar[8] ), .B2(
        n325), .C1(n284), .C2(n1154), .ZN(n1152) );
  INV_X1 U2426 ( .A(n5679), .ZN(n1154) );
  AOI22_X1 U2427 ( .A1(n6379), .A2(n6190), .B1(
        \UUT/Mpath/the_mult/x_mult_out[8] ), .B2(n291), .ZN(n1151) );
  OAI222_X1 U2428 ( .A1(n77), .A2(n123), .B1(n76), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N64 ), .C2(net54895), .ZN(n4325) );
  INV_X1 U2429 ( .A(\UUT/break_code[10] ), .ZN(n76) );
  INV_X1 U2430 ( .A(n1155), .ZN(n77) );
  OAI222_X1 U2431 ( .A1(n602), .A2(n129), .B1(n959), .B2(n131), .C1(n5523), 
        .C2(n132), .ZN(n1155) );
  OAI211_X1 U2433 ( .C1(n482), .C2(n1156), .A(n484), .B(n1157), .ZN(n605) );
  AOI22_X1 U2434 ( .A1(n486), .A2(n781), .B1(n1158), .B2(n489), .ZN(n1157) );
  INV_X1 U2435 ( .A(n5524), .ZN(n1158) );
  INV_X1 U2436 ( .A(n5845), .ZN(n781) );
  AND2_X1 U2437 ( .A1(n5713), .A2(n5710), .ZN(n486) );
  INV_X1 U2438 ( .A(n5838), .ZN(n1156) );
  NAND2_X1 U2439 ( .A1(n5711), .A2(n5710), .ZN(n482) );
  INV_X1 U2440 ( .A(n1159), .ZN(n602) );
  OAI211_X1 U2441 ( .C1(n5674), .C2(n321), .A(n1160), .B(n1161), .ZN(n1159) );
  AOI222_X1 U2442 ( .A1(n285), .A2(n1162), .B1(\UUT/Mpath/out_jar[10] ), .B2(
        n325), .C1(n284), .C2(n1163), .ZN(n1161) );
  INV_X1 U2443 ( .A(n5708), .ZN(n1163) );
  AOI22_X1 U2444 ( .A1(n6379), .A2(n6205), .B1(
        \UUT/Mpath/the_mult/x_mult_out[10] ), .B2(n291), .ZN(n1160) );
  OAI22_X1 U2445 ( .A1(\UUT/Mpath/the_alu/N22 ), .A2(net54877), .B1(net54921), 
        .B2(n74), .ZN(n4327) );
  INV_X1 U2446 ( .A(n1164), .ZN(n74) );
  OAI211_X1 U2447 ( .C1(n789), .C2(n115), .A(n856), .B(n1165), .ZN(n1164) );
  NOR2_X1 U2448 ( .A1(n854), .A2(n1166), .ZN(n1165) );
  NOR3_X1 U2449 ( .A1(n450), .A2(n5831), .A3(n1167), .ZN(n1166) );
  AND2_X1 U2450 ( .A1(n5869), .A2(n207), .ZN(n854) );
  AOI21_X1 U2451 ( .B1(n5870), .B2(n207), .A(n448), .ZN(n856) );
  NOR2_X1 U2452 ( .A1(n450), .A2(n1168), .ZN(n207) );
  OR2_X1 U2453 ( .A1(n1169), .A2(n175), .ZN(n450) );
  INV_X1 U2454 ( .A(n1170), .ZN(n115) );
  OAI222_X1 U2455 ( .A1(n953), .A2(n129), .B1(n952), .B2(n131), .C1(n5454), 
        .C2(n132), .ZN(n1170) );
  AND2_X1 U2458 ( .A1(n484), .A2(n1172), .ZN(n282) );
  NAND2_X1 U2459 ( .A1(n5945), .A2(n5710), .ZN(n1172) );
  NAND2_X1 U2460 ( .A1(n5715), .A2(n5710), .ZN(n484) );
  NAND3_X1 U2461 ( .A1(n5950), .A2(n5710), .A3(n5951), .ZN(n281) );
  INV_X1 U2462 ( .A(n175), .ZN(n789) );
  OAI22_X1 U2463 ( .A1(n5455), .A2(net54877), .B1(net54919), .B2(n953), .ZN(
        n4328) );
  AOI221_X1 U2464 ( .B1(n1173), .B2(n284), .C1(n6197), .C2(n285), .A(n1174), 
        .ZN(n953) );
  INV_X1 U2465 ( .A(n1175), .ZN(n1174) );
  AOI222_X1 U2466 ( .A1(n288), .A2(n1176), .B1(n6379), .B2(n6644), .C1(
        \UUT/Mpath/the_mult/x_mult_out[31] ), .C2(n291), .ZN(n1175) );
  INV_X1 U2467 ( .A(n5628), .ZN(n1176) );
  INV_X1 U2468 ( .A(n321), .ZN(n288) );
  INV_X1 U2469 ( .A(n5685), .ZN(n1173) );
  INV_X1 U2472 ( .A(n5629), .ZN(n948) );
  INV_X1 U2473 ( .A(\UUT/Mpath/the_mult/Mult_out[63] ), .ZN(n1142) );
  OAI221_X1 U2474 ( .B1(n133), .B2(n1110), .C1(n5709), .C2(n135), .A(n1178), 
        .ZN(n4330) );
  AOI22_X1 U2475 ( .A1(n137), .A2(n970), .B1(\UUT/Mpath/the_mult/Mad_out [32]), 
        .B2(n139), .ZN(n1178) );
  INV_X1 U2478 ( .A(n5677), .ZN(n970) );
  INV_X1 U2485 ( .A(\UUT/Mpath/the_mult/Mult_out[32] ), .ZN(n1110) );
  AND2_X1 U2487 ( .A1(n5413), .A2(net54895), .ZN(n975) );
  OAI22_X1 U2488 ( .A1(net54913), .A2(n1184), .B1(n5677), .B2(net54875), .ZN(
        n4331) );
  OAI221_X1 U2489 ( .B1(n1073), .B2(n310), .C1(n147), .C2(n1184), .A(n1185), 
        .ZN(n4332) );
  AOI22_X1 U2490 ( .A1(n312), .A2(n1075), .B1(n314), .B2(n1076), .ZN(n1185) );
  INV_X1 U2493 ( .A(\UUT/Mpath/the_mult/x_operand1[0] ), .ZN(n1184) );
  NAND2_X1 U2494 ( .A1(n147), .A2(n1077), .ZN(n310) );
  INV_X1 U2495 ( .A(n5528), .ZN(n1077) );
  OAI21_X1 U2497 ( .B1(\UUT/Mpath/the_mult/N227 ), .B2(
        \UUT/Mpath/the_mult/N223 ), .A(net54859), .ZN(n73) );
  OAI22_X1 U2498 ( .A1(net54847), .A2(\UUT/Mpath/N111 ), .B1(n6069), .B2(n945), 
        .ZN(n4333) );
  NAND2_X1 U2499 ( .A1(n1186), .A2(net54857), .ZN(n945) );
  NAND4_X1 U2500 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2025 ), .A2(n935), 
        .A3(n931), .A4(n937), .ZN(n1186) );
  OAI22_X1 U2501 ( .A1(n546), .A2(n1187), .B1(n6069), .B2(n295), .ZN(n4334) );
  INV_X1 U2503 ( .A(I_DATA_INBUS[31]), .ZN(n1187) );
  INV_X1 U2505 ( .A(\UUT/Mcontrol/st_logic/N10 ), .ZN(n978) );
  OAI222_X1 U2506 ( .A1(n70), .A2(n123), .B1(n68), .B2(n300), .C1(
        \UUT/Mpath/the_alu/N84 ), .C2(net54895), .ZN(n4335) );
  INV_X1 U2507 ( .A(n449), .ZN(n300) );
  NOR2_X1 U2508 ( .A1(n175), .A2(net54933), .ZN(n449) );
  INV_X1 U2510 ( .A(n6588), .ZN(n68) );
  NAND2_X1 U2511 ( .A1(n175), .A2(net54859), .ZN(n123) );
  OAI21_X1 U2512 ( .B1(n6206), .B2(n6170), .A(n6030), .ZN(n175) );
  INV_X1 U2513 ( .A(n1188), .ZN(n70) );
  OAI222_X1 U2514 ( .A1(n5526), .A2(n132), .B1(n960), .B2(n131), .C1(n1073), 
        .C2(n129), .ZN(n1188) );
  INV_X1 U2516 ( .A(n1189), .ZN(n1073) );
  OAI211_X1 U2517 ( .C1(n5676), .C2(n321), .A(n1190), .B(n1191), .ZN(n1189) );
  AOI222_X1 U2518 ( .A1(n285), .A2(n5613), .B1(\UUT/Mpath/out_jar[0] ), .B2(
        n325), .C1(n284), .C2(n1192), .ZN(n1191) );
  INV_X1 U2519 ( .A(n5709), .ZN(n1192) );
  INV_X1 U2521 ( .A(n1194), .ZN(n1193) );
  AOI22_X1 U2523 ( .A1(n6379), .A2(\UUT/daddr_out [0]), .B1(
        \UUT/Mpath/the_mult/x_mult_out[0] ), .B2(n291), .ZN(n1190) );
  NOR3_X1 U2525 ( .A1(n1195), .A2(n285), .A3(n1196), .ZN(n290) );
  INV_X1 U2526 ( .A(\UUT/Mpath/N128 ), .ZN(n1196) );
  INV_X1 U2527 ( .A(\UUT/Mpath/N125 ), .ZN(n1195) );
  NAND3_X1 U2528 ( .A1(n1194), .A2(n1197), .A3(\UUT/Mpath/the_mult/N216 ), 
        .ZN(n321) );
  INV_X1 U2529 ( .A(\UUT/Mpath/the_mult/N198 ), .ZN(n1197) );
  NOR2_X1 U2530 ( .A1(n285), .A2(\UUT/Mpath/N125 ), .ZN(n1194) );
  OAI211_X1 U2534 ( .C1(n5710), .C2(n5527), .A(n1198), .B(n1199), .ZN(n1076)
         );
  AOI222_X1 U2535 ( .A1(n5747), .A2(n684), .B1(n685), .B2(n1148), .C1(n6000), 
        .C2(n686), .ZN(n1199) );
  AND2_X1 U2536 ( .A1(n687), .A2(\UUT/Mpath/the_memhandle/N37 ), .ZN(n686) );
  INV_X1 U2537 ( .A(n5999), .ZN(n1148) );
  AND2_X1 U2538 ( .A1(n5757), .A2(n688), .ZN(n685) );
  AND2_X1 U2539 ( .A1(n5710), .A2(n1200), .ZN(n684) );
  OAI22_X1 U2540 ( .A1(n5985), .A2(n1201), .B1(\UUT/Mpath/the_memhandle/N34 ), 
        .B2(n1202), .ZN(n1200) );
  INV_X1 U2541 ( .A(n5755), .ZN(n1202) );
  AOI22_X1 U2542 ( .A1(n6001), .A2(n687), .B1(n5994), .B2(n688), .ZN(n1198) );
  INV_X1 U2543 ( .A(n660), .ZN(n688) );
  NAND2_X1 U2544 ( .A1(n5710), .A2(n1201), .ZN(n660) );
  NOR2_X1 U2545 ( .A1(n1201), .A2(n489), .ZN(n687) );
  INV_X1 U2546 ( .A(n5710), .ZN(n489) );
  INV_X1 U2547 ( .A(\UUT/Mpath/the_memhandle/N34 ), .ZN(n1201) );
  NAND2_X1 U2549 ( .A1(n1203), .A2(n1204), .ZN(n6197) );
  AOI222_X1 U2550 ( .A1(\UUT/Mpath/the_shift/sh_ror [31]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [31]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [31]), .C2(n6199), .ZN(n1204) );
  AOI22_X1 U2551 ( .A1(\UUT/Mpath/the_shift/sh_sll [31]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [31]), .B2(n6198), .ZN(n1203) );
  INV_X1 U2554 ( .A(\UUT/Mpath/the_alu/N21 ), .ZN(n1209) );
  AOI22_X1 U2555 ( .A1(\UUT/Mpath/the_alu/N126 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N94 ), .B2(n1213), .ZN(n1206) );
  AOI22_X1 U2556 ( .A1(\UUT/Mpath/the_alu/N158 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N190 ), .B2(n1215), .ZN(n1205) );
  INV_X1 U2557 ( .A(n1216), .ZN(n6116) );
  NOR4_X1 U2558 ( .A1(n1217), .A2(n1008), .A3(n6067), .A4(n6079), .ZN(n6076)
         );
  INV_X1 U2559 ( .A(\UUT/Mcontrol/Operation_decoding32/N1945 ), .ZN(n1008) );
  INV_X1 U2560 ( .A(n6285), .ZN(n1217) );
  NAND3_X1 U2561 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1975 ), .A2(n445), 
        .A3(n857), .ZN(n6074) );
  INV_X1 U2562 ( .A(n937), .ZN(n6073) );
  NOR2_X1 U2563 ( .A1(n1218), .A2(n1219), .ZN(n937) );
  INV_X1 U2564 ( .A(n932), .ZN(n1218) );
  INV_X1 U2565 ( .A(\UUT/Mcontrol/d_sampled_finstr [29]), .ZN(n6071) );
  INV_X1 U2566 ( .A(\UUT/Mcontrol/d_sampled_finstr [30]), .ZN(n6070) );
  INV_X1 U2567 ( .A(\UUT/Mcontrol/d_sampled_finstr [31]), .ZN(n6069) );
  INV_X1 U2568 ( .A(\UUT/Mcontrol/Operation_decoding32/N2019 ), .ZN(n6051) );
  INV_X1 U2570 ( .A(n6078), .ZN(n6048) );
  INV_X1 U2571 ( .A(\UUT/Mcontrol/d_sampled_finstr [21]), .ZN(n6037) );
  INV_X1 U2572 ( .A(\UUT/Mcontrol/d_sampled_finstr [17]), .ZN(n6034) );
  INV_X1 U2573 ( .A(\UUT/Mcontrol/d_sampled_finstr [19]), .ZN(n6031) );
  INV_X1 U2574 ( .A(\UUT/Mcontrol/d_sampled_finstr [20]), .ZN(n6029) );
  INV_X1 U2575 ( .A(\UUT/Mcontrol/Operation_decoding32/N2043 ), .ZN(n6028) );
  INV_X1 U2576 ( .A(\UUT/Mcontrol/d_sampled_finstr [16]), .ZN(n6027) );
  INV_X1 U2577 ( .A(\UUT/Mcontrol/d_sampled_finstr [18]), .ZN(n6026) );
  AOI22_X1 U2578 ( .A1(dram_data_inbus[16]), .A2(n5779), .B1(
        BUS_DATA_INBUS[16]), .B2(n6377), .ZN(n5944) );
  AOI22_X1 U2579 ( .A1(dram_data_inbus[17]), .A2(n5779), .B1(
        BUS_DATA_INBUS[17]), .B2(n6377), .ZN(n5919) );
  INV_X1 U2580 ( .A(\UUT/Mcontrol/d_sampled_finstr [22]), .ZN(n5896) );
  AOI22_X1 U2581 ( .A1(dram_data_inbus[24]), .A2(n5779), .B1(
        BUS_DATA_INBUS[24]), .B2(n6377), .ZN(n5890) );
  INV_X1 U2582 ( .A(\UUT/Mcontrol/d_sampled_finstr [23]), .ZN(n5888) );
  AOI22_X1 U2583 ( .A1(dram_data_inbus[25]), .A2(n5779), .B1(
        BUS_DATA_INBUS[25]), .B2(n6377), .ZN(n5882) );
  INV_X1 U2584 ( .A(n5870), .ZN(n5880) );
  INV_X1 U2585 ( .A(\UUT/Mcontrol/d_sampled_finstr [24]), .ZN(n5879) );
  AOI22_X1 U2586 ( .A1(dram_data_inbus[26]), .A2(n5779), .B1(
        BUS_DATA_INBUS[26]), .B2(n6377), .ZN(n5873) );
  NAND2_X1 U2587 ( .A1(n1220), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .ZN(n5872) );
  INV_X1 U2588 ( .A(n6118), .ZN(n1220) );
  INV_X1 U2589 ( .A(\UUT/Mcontrol/d_sampled_finstr [25]), .ZN(n5871) );
  AOI22_X1 U2590 ( .A1(dram_data_inbus[27]), .A2(n5779), .B1(
        BUS_DATA_INBUS[27]), .B2(n6377), .ZN(n5863) );
  AOI22_X1 U2591 ( .A1(dram_data_inbus[28]), .A2(n5779), .B1(
        BUS_DATA_INBUS[28]), .B2(n6377), .ZN(n5857) );
  AOI22_X1 U2592 ( .A1(dram_data_inbus[29]), .A2(n5779), .B1(
        BUS_DATA_INBUS[29]), .B2(n6377), .ZN(n5851) );
  AOI22_X1 U2593 ( .A1(dram_data_inbus[18]), .A2(n5779), .B1(
        BUS_DATA_INBUS[18]), .B2(n6377), .ZN(n5841) );
  AOI22_X1 U2594 ( .A1(dram_data_inbus[30]), .A2(n5779), .B1(
        BUS_DATA_INBUS[30]), .B2(n6377), .ZN(n5832) );
  AOI22_X1 U2595 ( .A1(n5779), .A2(dram_data_inbus[31]), .B1(n6377), .B2(
        BUS_DATA_INBUS[31]), .ZN(n5825) );
  AOI22_X1 U2596 ( .A1(dram_data_inbus[19]), .A2(n5779), .B1(
        BUS_DATA_INBUS[19]), .B2(n6377), .ZN(n5815) );
  AOI22_X1 U2597 ( .A1(dram_data_inbus[20]), .A2(n5779), .B1(
        BUS_DATA_INBUS[20]), .B2(n6377), .ZN(n5802) );
  AOI22_X1 U2598 ( .A1(dram_data_inbus[21]), .A2(n5779), .B1(
        BUS_DATA_INBUS[21]), .B2(n6377), .ZN(n5789) );
  AOI22_X1 U2599 ( .A1(dram_data_inbus[22]), .A2(n5779), .B1(
        BUS_DATA_INBUS[22]), .B2(n6377), .ZN(n5772) );
  AOI22_X1 U2600 ( .A1(dram_data_inbus[23]), .A2(n5779), .B1(
        BUS_DATA_INBUS[23]), .B2(n6377), .ZN(n5760) );
  OAI21_X1 U2601 ( .B1(n5984), .B2(n5983), .A(\UUT/Mpath/the_memhandle/N34 ), 
        .ZN(n5754) );
  NAND2_X1 U2602 ( .A1(n1221), .A2(n1222), .ZN(n5613) );
  AOI222_X1 U2603 ( .A1(n6378), .A2(\UUT/Mpath/the_shift/sh_ror [0]), .B1(
        \UUT/Mpath/the_shift/sh_srl [0]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(n6199), .C2(\UUT/Mpath/the_shift/sh_rol [0]), .ZN(n1222) );
  AOI22_X1 U2604 ( .A1(n6200), .A2(\UUT/Mpath/the_shift/sh_sll [0]), .B1(n6198), .B2(\UUT/Mpath/the_shift/sh_sra [0]), .ZN(n1221) );
  NAND3_X1 U2605 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n5606) );
  AOI222_X1 U2606 ( .A1(n1208), .A2(n1226), .B1(\UUT/Mpath/the_alu/diff[24] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[24] ), .C2(n1211), .ZN(n1225)
         );
  INV_X1 U2607 ( .A(\UUT/Mpath/the_alu/N35 ), .ZN(n1226) );
  AOI22_X1 U2608 ( .A1(\UUT/Mpath/the_alu/N133 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N101 ), .B2(n1213), .ZN(n1224) );
  AOI22_X1 U2609 ( .A1(\UUT/Mpath/the_alu/N165 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N197 ), .B2(n1215), .ZN(n1223) );
  NAND2_X1 U2610 ( .A1(n1227), .A2(n1228), .ZN(n5605) );
  AOI222_X1 U2611 ( .A1(\UUT/Mpath/the_shift/sh_ror [24]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [24]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [24]), .C2(n6199), .ZN(n1228) );
  AOI22_X1 U2612 ( .A1(\UUT/Mpath/the_shift/sh_sll [24]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [24]), .B2(n6198), .ZN(n1227) );
  NAND3_X1 U2613 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n5599) );
  AOI222_X1 U2614 ( .A1(n1208), .A2(n1232), .B1(\UUT/Mpath/the_alu/diff[25] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[25] ), .C2(n1211), .ZN(n1231)
         );
  INV_X1 U2615 ( .A(\UUT/Mpath/the_alu/N33 ), .ZN(n1232) );
  AOI22_X1 U2616 ( .A1(\UUT/Mpath/the_alu/N132 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N100 ), .B2(n1213), .ZN(n1230) );
  AOI22_X1 U2617 ( .A1(\UUT/Mpath/the_alu/N164 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N196 ), .B2(n1215), .ZN(n1229) );
  NAND2_X1 U2618 ( .A1(n1233), .A2(n1234), .ZN(n5598) );
  AOI222_X1 U2619 ( .A1(\UUT/Mpath/the_shift/sh_ror [25]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [25]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [25]), .C2(n6199), .ZN(n1234) );
  AOI22_X1 U2620 ( .A1(\UUT/Mpath/the_shift/sh_sll [25]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [25]), .B2(n6198), .ZN(n1233) );
  INV_X1 U2623 ( .A(\UUT/Mpath/the_alu/N31 ), .ZN(n1238) );
  AOI22_X1 U2624 ( .A1(\UUT/Mpath/the_alu/N131 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N99 ), .B2(n1213), .ZN(n1236) );
  AOI22_X1 U2625 ( .A1(\UUT/Mpath/the_alu/N163 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N195 ), .B2(n1215), .ZN(n1235) );
  NAND2_X1 U2626 ( .A1(n1239), .A2(n1240), .ZN(n5591) );
  AOI222_X1 U2627 ( .A1(\UUT/Mpath/the_shift/sh_ror [26]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [26]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [26]), .C2(n6199), .ZN(n1240) );
  AOI22_X1 U2628 ( .A1(\UUT/Mpath/the_shift/sh_sll [26]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [26]), .B2(n6198), .ZN(n1239) );
  INV_X1 U2631 ( .A(\UUT/Mpath/the_alu/N29 ), .ZN(n1244) );
  AOI22_X1 U2632 ( .A1(\UUT/Mpath/the_alu/N130 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N98 ), .B2(n1213), .ZN(n1242) );
  AOI22_X1 U2633 ( .A1(\UUT/Mpath/the_alu/N162 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N194 ), .B2(n1215), .ZN(n1241) );
  NAND2_X1 U2634 ( .A1(n1245), .A2(n1246), .ZN(n5584) );
  AOI222_X1 U2635 ( .A1(\UUT/Mpath/the_shift/sh_ror [27]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [27]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [27]), .C2(n6199), .ZN(n1246) );
  AOI22_X1 U2636 ( .A1(\UUT/Mpath/the_shift/sh_sll [27]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [27]), .B2(n6198), .ZN(n1245) );
  INV_X1 U2639 ( .A(\UUT/Mpath/the_alu/N27 ), .ZN(n1250) );
  AOI22_X1 U2640 ( .A1(\UUT/Mpath/the_alu/N129 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N97 ), .B2(n1213), .ZN(n1248) );
  AOI22_X1 U2641 ( .A1(\UUT/Mpath/the_alu/N161 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N193 ), .B2(n1215), .ZN(n1247) );
  NAND2_X1 U2642 ( .A1(n1251), .A2(n1252), .ZN(n5577) );
  AOI222_X1 U2643 ( .A1(\UUT/Mpath/the_shift/sh_ror [28]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [28]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [28]), .C2(n6199), .ZN(n1252) );
  AOI22_X1 U2644 ( .A1(\UUT/Mpath/the_shift/sh_sll [28]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [28]), .B2(n6198), .ZN(n1251) );
  INV_X1 U2647 ( .A(\UUT/Mpath/the_alu/N25 ), .ZN(n1256) );
  AOI22_X1 U2648 ( .A1(\UUT/Mpath/the_alu/N128 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N96 ), .B2(n1213), .ZN(n1254) );
  AOI22_X1 U2649 ( .A1(\UUT/Mpath/the_alu/N160 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N192 ), .B2(n1215), .ZN(n1253) );
  NAND2_X1 U2650 ( .A1(n1257), .A2(n1258), .ZN(n5570) );
  AOI222_X1 U2651 ( .A1(\UUT/Mpath/the_shift/sh_ror [29]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [29]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [29]), .C2(n6199), .ZN(n1258) );
  AOI22_X1 U2652 ( .A1(\UUT/Mpath/the_shift/sh_sll [29]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [29]), .B2(n6198), .ZN(n1257) );
  INV_X1 U2655 ( .A(\UUT/Mpath/the_alu/N23 ), .ZN(n1262) );
  AOI22_X1 U2656 ( .A1(\UUT/Mpath/the_alu/N127 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N95 ), .B2(n1213), .ZN(n1260) );
  AOI22_X1 U2657 ( .A1(\UUT/Mpath/the_alu/N159 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N191 ), .B2(n1215), .ZN(n1259) );
  NAND2_X1 U2658 ( .A1(n1263), .A2(n1264), .ZN(n5562) );
  AOI222_X1 U2659 ( .A1(\UUT/Mpath/the_shift/sh_ror [30]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [30]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [30]), .C2(n6199), .ZN(n1264) );
  AOI22_X1 U2660 ( .A1(\UUT/Mpath/the_shift/sh_sll [30]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [30]), .B2(n6198), .ZN(n1263) );
  AND4_X1 U2661 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n5526)
         );
  NOR4_X1 U2662 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1268)
         );
  NAND3_X1 U2663 ( .A1(n6019), .A2(n6015), .A3(n6024), .ZN(n1272) );
  OAI211_X1 U2664 ( .C1(n5745), .C2(n5412), .A(n6004), .B(n6011), .ZN(n1271)
         );
  OAI222_X1 U2665 ( .A1(n5743), .A2(n5284), .B1(n5744), .B2(n5252), .C1(n5746), 
        .C2(n5380), .ZN(n1270) );
  OAI221_X1 U2666 ( .B1(n5716), .B2(n5188), .C1(n5717), .C2(n5220), .A(n1273), 
        .ZN(n1269) );
  AOI22_X1 U2667 ( .A1(n1274), .A2(n1275), .B1(n1276), .B2(n1277), .ZN(n1273)
         );
  AOI211_X1 U2668 ( .C1(n1278), .C2(n1279), .A(n1280), .B(n1281), .ZN(n1267)
         );
  OAI22_X1 U2669 ( .A1(n5726), .A2(n4836), .B1(n5736), .B2(n4740), .ZN(n1281)
         );
  OAI222_X1 U2670 ( .A1(n5731), .A2(n4676), .B1(n5737), .B2(n4644), .C1(n5732), 
        .C2(n4708), .ZN(n1280) );
  AOI221_X1 U2671 ( .B1(n1282), .B2(n1283), .C1(n1284), .C2(n1285), .A(n1286), 
        .ZN(n1266) );
  OAI22_X1 U2672 ( .A1(n4484), .A2(n1287), .B1(n5316), .B2(n1288), .ZN(n1286)
         );
  INV_X1 U2673 ( .A(n5092), .ZN(n1283) );
  AOI222_X1 U2674 ( .A1(n1289), .A2(n1290), .B1(n1291), .B2(n1292), .C1(n1293), 
        .C2(n1294), .ZN(n1265) );
  AND4_X1 U2675 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n5523)
         );
  NOR4_X1 U2676 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1298)
         );
  NAND3_X1 U2677 ( .A1(n5992), .A2(n5991), .A3(n5993), .ZN(n1302) );
  OAI211_X1 U2678 ( .C1(n5745), .C2(n5411), .A(n5989), .B(n5990), .ZN(n1301)
         );
  OAI222_X1 U2679 ( .A1(n5743), .A2(n5283), .B1(n5744), .B2(n5251), .C1(n5746), 
        .C2(n5379), .ZN(n1300) );
  OAI221_X1 U2680 ( .B1(n5716), .B2(n5187), .C1(n5717), .C2(n5219), .A(n1303), 
        .ZN(n1299) );
  AOI22_X1 U2681 ( .A1(n1304), .A2(n1275), .B1(n1305), .B2(n1277), .ZN(n1303)
         );
  AOI211_X1 U2682 ( .C1(n1306), .C2(n1279), .A(n1307), .B(n1308), .ZN(n1297)
         );
  OAI22_X1 U2683 ( .A1(n5726), .A2(n4835), .B1(n5736), .B2(n4739), .ZN(n1308)
         );
  OAI222_X1 U2684 ( .A1(n5731), .A2(n4675), .B1(n5737), .B2(n4643), .C1(n5732), 
        .C2(n4707), .ZN(n1307) );
  AOI221_X1 U2685 ( .B1(n1282), .B2(n1309), .C1(n1284), .C2(n1310), .A(n1311), 
        .ZN(n1296) );
  OAI22_X1 U2686 ( .A1(n4483), .A2(n1287), .B1(n5315), .B2(n1288), .ZN(n1311)
         );
  INV_X1 U2687 ( .A(n5091), .ZN(n1309) );
  AOI222_X1 U2688 ( .A1(n1312), .A2(n1290), .B1(n1291), .B2(n1313), .C1(n1314), 
        .C2(n1294), .ZN(n1295) );
  AND4_X1 U2689 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n5520)
         );
  NOR4_X1 U2690 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1318)
         );
  NAND3_X1 U2691 ( .A1(n5981), .A2(n5980), .A3(n5982), .ZN(n1322) );
  OAI211_X1 U2692 ( .C1(n5745), .C2(n5410), .A(n5978), .B(n5979), .ZN(n1321)
         );
  OAI222_X1 U2693 ( .A1(n5743), .A2(n5282), .B1(n5744), .B2(n5250), .C1(n5746), 
        .C2(n5378), .ZN(n1320) );
  OAI221_X1 U2694 ( .B1(n5716), .B2(n5186), .C1(n5717), .C2(n5218), .A(n1323), 
        .ZN(n1319) );
  AOI22_X1 U2695 ( .A1(n1324), .A2(n1275), .B1(n1325), .B2(n1277), .ZN(n1323)
         );
  AOI211_X1 U2696 ( .C1(n1326), .C2(n1279), .A(n1327), .B(n1328), .ZN(n1317)
         );
  OAI22_X1 U2697 ( .A1(n5726), .A2(n4834), .B1(n5736), .B2(n4738), .ZN(n1328)
         );
  OAI222_X1 U2698 ( .A1(n5731), .A2(n4674), .B1(n5737), .B2(n4642), .C1(n5732), 
        .C2(n4706), .ZN(n1327) );
  AOI221_X1 U2699 ( .B1(n1282), .B2(n1329), .C1(n1284), .C2(n1330), .A(n1331), 
        .ZN(n1316) );
  OAI22_X1 U2700 ( .A1(n4482), .A2(n1287), .B1(n5314), .B2(n1288), .ZN(n1331)
         );
  INV_X1 U2701 ( .A(n5090), .ZN(n1329) );
  AOI222_X1 U2702 ( .A1(n1332), .A2(n1290), .B1(n1291), .B2(n1333), .C1(n1334), 
        .C2(n1294), .ZN(n1315) );
  AND4_X1 U2703 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n5517)
         );
  NOR4_X1 U2704 ( .A1(n1339), .A2(n1340), .A3(n1341), .A4(n1342), .ZN(n1338)
         );
  NAND3_X1 U2705 ( .A1(n5976), .A2(n5975), .A3(n5977), .ZN(n1342) );
  OAI211_X1 U2706 ( .C1(n5745), .C2(n5409), .A(n5973), .B(n5974), .ZN(n1341)
         );
  OAI222_X1 U2707 ( .A1(n5743), .A2(n5281), .B1(n5744), .B2(n5249), .C1(n5746), 
        .C2(n5377), .ZN(n1340) );
  OAI221_X1 U2708 ( .B1(n5716), .B2(n5185), .C1(n5717), .C2(n5217), .A(n1343), 
        .ZN(n1339) );
  AOI22_X1 U2709 ( .A1(n1344), .A2(n1275), .B1(n1345), .B2(n1277), .ZN(n1343)
         );
  AOI211_X1 U2710 ( .C1(n1346), .C2(n1279), .A(n1347), .B(n1348), .ZN(n1337)
         );
  OAI22_X1 U2711 ( .A1(n5726), .A2(n4833), .B1(n5736), .B2(n4737), .ZN(n1348)
         );
  OAI222_X1 U2712 ( .A1(n5731), .A2(n4673), .B1(n5737), .B2(n4641), .C1(n5732), 
        .C2(n4705), .ZN(n1347) );
  AOI221_X1 U2713 ( .B1(n1282), .B2(n1349), .C1(n1284), .C2(n1350), .A(n1351), 
        .ZN(n1336) );
  OAI22_X1 U2714 ( .A1(n4481), .A2(n1287), .B1(n5313), .B2(n1288), .ZN(n1351)
         );
  INV_X1 U2715 ( .A(n5089), .ZN(n1349) );
  AOI222_X1 U2716 ( .A1(n1352), .A2(n1290), .B1(n1291), .B2(n1353), .C1(n1354), 
        .C2(n1294), .ZN(n1335) );
  AND4_X1 U2717 ( .A1(n1355), .A2(n1356), .A3(n1357), .A4(n1358), .ZN(n5514)
         );
  NOR4_X1 U2718 ( .A1(n1359), .A2(n1360), .A3(n1361), .A4(n1362), .ZN(n1358)
         );
  NAND3_X1 U2719 ( .A1(n5971), .A2(n5970), .A3(n5972), .ZN(n1362) );
  OAI211_X1 U2720 ( .C1(n5745), .C2(n5408), .A(n5968), .B(n5969), .ZN(n1361)
         );
  OAI222_X1 U2721 ( .A1(n5743), .A2(n5280), .B1(n5744), .B2(n5248), .C1(n5746), 
        .C2(n5376), .ZN(n1360) );
  OAI221_X1 U2722 ( .B1(n5716), .B2(n5184), .C1(n5717), .C2(n5216), .A(n1363), 
        .ZN(n1359) );
  AOI22_X1 U2723 ( .A1(n1364), .A2(n1275), .B1(n1365), .B2(n1277), .ZN(n1363)
         );
  AOI211_X1 U2724 ( .C1(n1366), .C2(n1279), .A(n1367), .B(n1368), .ZN(n1357)
         );
  OAI22_X1 U2725 ( .A1(n5726), .A2(n4832), .B1(n5736), .B2(n4736), .ZN(n1368)
         );
  OAI222_X1 U2726 ( .A1(n5731), .A2(n4672), .B1(n5737), .B2(n4640), .C1(n5732), 
        .C2(n4704), .ZN(n1367) );
  AOI221_X1 U2727 ( .B1(n1282), .B2(n1369), .C1(n1284), .C2(n1370), .A(n1371), 
        .ZN(n1356) );
  OAI22_X1 U2728 ( .A1(n4480), .A2(n1287), .B1(n5312), .B2(n1288), .ZN(n1371)
         );
  INV_X1 U2729 ( .A(n5088), .ZN(n1369) );
  AOI222_X1 U2730 ( .A1(n1372), .A2(n1290), .B1(n1291), .B2(n1373), .C1(n1374), 
        .C2(n1294), .ZN(n1355) );
  AND4_X1 U2731 ( .A1(n1375), .A2(n1376), .A3(n1377), .A4(n1378), .ZN(n5511)
         );
  NOR4_X1 U2732 ( .A1(n1379), .A2(n1380), .A3(n1381), .A4(n1382), .ZN(n1378)
         );
  NAND3_X1 U2733 ( .A1(n5966), .A2(n5965), .A3(n5967), .ZN(n1382) );
  OAI211_X1 U2734 ( .C1(n5745), .C2(n5407), .A(n5963), .B(n5964), .ZN(n1381)
         );
  OAI222_X1 U2735 ( .A1(n5743), .A2(n5279), .B1(n5744), .B2(n5247), .C1(n5746), 
        .C2(n5375), .ZN(n1380) );
  OAI221_X1 U2736 ( .B1(n5716), .B2(n5183), .C1(n5717), .C2(n5215), .A(n1383), 
        .ZN(n1379) );
  AOI22_X1 U2737 ( .A1(n1384), .A2(n1275), .B1(n1385), .B2(n1277), .ZN(n1383)
         );
  AOI211_X1 U2738 ( .C1(n1386), .C2(n1279), .A(n1387), .B(n1388), .ZN(n1377)
         );
  OAI22_X1 U2739 ( .A1(n5726), .A2(n4831), .B1(n5736), .B2(n4735), .ZN(n1388)
         );
  OAI222_X1 U2740 ( .A1(n5731), .A2(n4671), .B1(n5737), .B2(n4639), .C1(n5732), 
        .C2(n4703), .ZN(n1387) );
  AOI221_X1 U2741 ( .B1(n1282), .B2(n1389), .C1(n1284), .C2(n1390), .A(n1391), 
        .ZN(n1376) );
  OAI22_X1 U2742 ( .A1(n4479), .A2(n1287), .B1(n5311), .B2(n1288), .ZN(n1391)
         );
  INV_X1 U2743 ( .A(n5087), .ZN(n1389) );
  AOI222_X1 U2744 ( .A1(n1392), .A2(n1290), .B1(n1291), .B2(n1393), .C1(n1394), 
        .C2(n1294), .ZN(n1375) );
  AND4_X1 U2745 ( .A1(n1395), .A2(n1396), .A3(n1397), .A4(n1398), .ZN(n5508)
         );
  NOR4_X1 U2746 ( .A1(n1399), .A2(n1400), .A3(n1401), .A4(n1402), .ZN(n1398)
         );
  NAND3_X1 U2747 ( .A1(n5961), .A2(n5960), .A3(n5962), .ZN(n1402) );
  OAI211_X1 U2748 ( .C1(n5745), .C2(n5406), .A(n5958), .B(n5959), .ZN(n1401)
         );
  OAI222_X1 U2749 ( .A1(n5743), .A2(n5278), .B1(n5744), .B2(n5246), .C1(n5746), 
        .C2(n5374), .ZN(n1400) );
  OAI221_X1 U2750 ( .B1(n5716), .B2(n5182), .C1(n5717), .C2(n5214), .A(n1403), 
        .ZN(n1399) );
  AOI22_X1 U2751 ( .A1(n1404), .A2(n1275), .B1(n1405), .B2(n1277), .ZN(n1403)
         );
  AOI211_X1 U2752 ( .C1(n1406), .C2(n1279), .A(n1407), .B(n1408), .ZN(n1397)
         );
  OAI22_X1 U2753 ( .A1(n5726), .A2(n4830), .B1(n5736), .B2(n4734), .ZN(n1408)
         );
  OAI222_X1 U2754 ( .A1(n5731), .A2(n4670), .B1(n5737), .B2(n4638), .C1(n5732), 
        .C2(n4702), .ZN(n1407) );
  AOI221_X1 U2755 ( .B1(n1282), .B2(n1409), .C1(n1284), .C2(n1410), .A(n1411), 
        .ZN(n1396) );
  OAI22_X1 U2756 ( .A1(n4478), .A2(n1287), .B1(n5310), .B2(n1288), .ZN(n1411)
         );
  INV_X1 U2757 ( .A(n5086), .ZN(n1409) );
  AOI222_X1 U2758 ( .A1(n1412), .A2(n1290), .B1(n1291), .B2(n1413), .C1(n1414), 
        .C2(n1294), .ZN(n1395) );
  AND4_X1 U2759 ( .A1(n1415), .A2(n1416), .A3(n1417), .A4(n1418), .ZN(n5505)
         );
  NOR4_X1 U2760 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1418)
         );
  NAND3_X1 U2761 ( .A1(n5955), .A2(n5954), .A3(n5956), .ZN(n1422) );
  OAI211_X1 U2762 ( .C1(n5745), .C2(n5405), .A(n5952), .B(n5953), .ZN(n1421)
         );
  OAI222_X1 U2763 ( .A1(n5743), .A2(n5277), .B1(n5744), .B2(n5245), .C1(n5746), 
        .C2(n5373), .ZN(n1420) );
  OAI221_X1 U2764 ( .B1(n5716), .B2(n5181), .C1(n5717), .C2(n5213), .A(n1423), 
        .ZN(n1419) );
  AOI22_X1 U2765 ( .A1(n1424), .A2(n1275), .B1(n1425), .B2(n1277), .ZN(n1423)
         );
  AOI211_X1 U2766 ( .C1(n1426), .C2(n1279), .A(n1427), .B(n1428), .ZN(n1417)
         );
  OAI22_X1 U2767 ( .A1(n5726), .A2(n4829), .B1(n5736), .B2(n4733), .ZN(n1428)
         );
  OAI222_X1 U2768 ( .A1(n5731), .A2(n4669), .B1(n5737), .B2(n4637), .C1(n5732), 
        .C2(n4701), .ZN(n1427) );
  AOI221_X1 U2769 ( .B1(n1282), .B2(n1429), .C1(n1284), .C2(n1430), .A(n1431), 
        .ZN(n1416) );
  OAI22_X1 U2770 ( .A1(n4477), .A2(n1287), .B1(n5309), .B2(n1288), .ZN(n1431)
         );
  INV_X1 U2771 ( .A(n5085), .ZN(n1429) );
  AOI222_X1 U2772 ( .A1(n1432), .A2(n1290), .B1(n1291), .B2(n1433), .C1(n1434), 
        .C2(n1294), .ZN(n1415) );
  AND4_X1 U2773 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .ZN(n5502)
         );
  NOR4_X1 U2774 ( .A1(n1439), .A2(n1440), .A3(n1441), .A4(n1442), .ZN(n1438)
         );
  NAND3_X1 U2775 ( .A1(n5942), .A2(n5941), .A3(n5943), .ZN(n1442) );
  OAI211_X1 U2776 ( .C1(n5745), .C2(n5404), .A(n5939), .B(n5940), .ZN(n1441)
         );
  OAI222_X1 U2777 ( .A1(n5743), .A2(n5276), .B1(n5744), .B2(n5244), .C1(n5746), 
        .C2(n5372), .ZN(n1440) );
  OAI221_X1 U2778 ( .B1(n5716), .B2(n5180), .C1(n5717), .C2(n5212), .A(n1443), 
        .ZN(n1439) );
  AOI22_X1 U2779 ( .A1(n1444), .A2(n1275), .B1(n1445), .B2(n1277), .ZN(n1443)
         );
  AOI211_X1 U2780 ( .C1(n1446), .C2(n1279), .A(n1447), .B(n1448), .ZN(n1437)
         );
  OAI22_X1 U2781 ( .A1(n5726), .A2(n4828), .B1(n5736), .B2(n4732), .ZN(n1448)
         );
  OAI222_X1 U2782 ( .A1(n5731), .A2(n4668), .B1(n5737), .B2(n4636), .C1(n5732), 
        .C2(n4700), .ZN(n1447) );
  AOI221_X1 U2783 ( .B1(n1282), .B2(n1449), .C1(n1284), .C2(n1450), .A(n1451), 
        .ZN(n1436) );
  OAI22_X1 U2784 ( .A1(n4476), .A2(n1287), .B1(n5308), .B2(n1288), .ZN(n1451)
         );
  INV_X1 U2785 ( .A(n5084), .ZN(n1449) );
  AOI222_X1 U2786 ( .A1(n1452), .A2(n1290), .B1(n1291), .B2(n1453), .C1(n1454), 
        .C2(n1294), .ZN(n1435) );
  AND4_X1 U2787 ( .A1(n1455), .A2(n1456), .A3(n1457), .A4(n1458), .ZN(n5499)
         );
  NOR4_X1 U2788 ( .A1(n1459), .A2(n1460), .A3(n1461), .A4(n1462), .ZN(n1458)
         );
  NAND3_X1 U2789 ( .A1(n5937), .A2(n5936), .A3(n5938), .ZN(n1462) );
  OAI211_X1 U2790 ( .C1(n5745), .C2(n5403), .A(n5934), .B(n5935), .ZN(n1461)
         );
  OAI222_X1 U2791 ( .A1(n5743), .A2(n5275), .B1(n5744), .B2(n5243), .C1(n5746), 
        .C2(n5371), .ZN(n1460) );
  OAI221_X1 U2792 ( .B1(n5716), .B2(n5179), .C1(n5717), .C2(n5211), .A(n1463), 
        .ZN(n1459) );
  AOI22_X1 U2793 ( .A1(n1464), .A2(n1275), .B1(n1465), .B2(n1277), .ZN(n1463)
         );
  AOI211_X1 U2794 ( .C1(n1466), .C2(n1279), .A(n1467), .B(n1468), .ZN(n1457)
         );
  OAI22_X1 U2795 ( .A1(n5726), .A2(n4827), .B1(n5736), .B2(n4731), .ZN(n1468)
         );
  OAI222_X1 U2796 ( .A1(n5731), .A2(n4667), .B1(n5737), .B2(n4635), .C1(n5732), 
        .C2(n4699), .ZN(n1467) );
  AOI221_X1 U2797 ( .B1(n1282), .B2(n1469), .C1(n1284), .C2(n1470), .A(n1471), 
        .ZN(n1456) );
  OAI22_X1 U2798 ( .A1(n4475), .A2(n1287), .B1(n5307), .B2(n1288), .ZN(n1471)
         );
  INV_X1 U2799 ( .A(n5083), .ZN(n1469) );
  AOI222_X1 U2800 ( .A1(n1472), .A2(n1290), .B1(n1291), .B2(n1473), .C1(n1474), 
        .C2(n1294), .ZN(n1455) );
  AND4_X1 U2801 ( .A1(n1475), .A2(n1476), .A3(n1477), .A4(n1478), .ZN(n5496)
         );
  NOR4_X1 U2802 ( .A1(n1479), .A2(n1480), .A3(n1481), .A4(n1482), .ZN(n1478)
         );
  NAND3_X1 U2803 ( .A1(n5932), .A2(n5931), .A3(n5933), .ZN(n1482) );
  OAI211_X1 U2804 ( .C1(n5745), .C2(n5402), .A(n5929), .B(n5930), .ZN(n1481)
         );
  OAI222_X1 U2805 ( .A1(n5743), .A2(n5274), .B1(n5744), .B2(n5242), .C1(n5746), 
        .C2(n5370), .ZN(n1480) );
  OAI221_X1 U2806 ( .B1(n5716), .B2(n5178), .C1(n5717), .C2(n5210), .A(n1483), 
        .ZN(n1479) );
  AOI22_X1 U2807 ( .A1(n1484), .A2(n1275), .B1(n1485), .B2(n1277), .ZN(n1483)
         );
  AOI211_X1 U2808 ( .C1(n1486), .C2(n1279), .A(n1487), .B(n1488), .ZN(n1477)
         );
  OAI22_X1 U2809 ( .A1(n5726), .A2(n4826), .B1(n5736), .B2(n4730), .ZN(n1488)
         );
  OAI222_X1 U2810 ( .A1(n5731), .A2(n4666), .B1(n5737), .B2(n4634), .C1(n5732), 
        .C2(n4698), .ZN(n1487) );
  AOI221_X1 U2811 ( .B1(n1282), .B2(n1489), .C1(n1284), .C2(n1490), .A(n1491), 
        .ZN(n1476) );
  OAI22_X1 U2812 ( .A1(n4474), .A2(n1287), .B1(n5306), .B2(n1288), .ZN(n1491)
         );
  INV_X1 U2813 ( .A(n5082), .ZN(n1489) );
  AOI222_X1 U2814 ( .A1(n1492), .A2(n1290), .B1(n1291), .B2(n1493), .C1(n1494), 
        .C2(n1294), .ZN(n1475) );
  AND4_X1 U2815 ( .A1(n1495), .A2(n1496), .A3(n1497), .A4(n1498), .ZN(n5493)
         );
  NOR4_X1 U2816 ( .A1(n1499), .A2(n1500), .A3(n1501), .A4(n1502), .ZN(n1498)
         );
  NAND3_X1 U2817 ( .A1(n5927), .A2(n5926), .A3(n5928), .ZN(n1502) );
  OAI211_X1 U2818 ( .C1(n5745), .C2(n5401), .A(n5924), .B(n5925), .ZN(n1501)
         );
  OAI222_X1 U2819 ( .A1(n5743), .A2(n5273), .B1(n5744), .B2(n5241), .C1(n5746), 
        .C2(n5369), .ZN(n1500) );
  OAI221_X1 U2820 ( .B1(n5716), .B2(n5177), .C1(n5717), .C2(n5209), .A(n1503), 
        .ZN(n1499) );
  AOI22_X1 U2821 ( .A1(n1504), .A2(n1275), .B1(n1505), .B2(n1277), .ZN(n1503)
         );
  AOI211_X1 U2822 ( .C1(n1506), .C2(n1279), .A(n1507), .B(n1508), .ZN(n1497)
         );
  OAI22_X1 U2823 ( .A1(n5726), .A2(n4825), .B1(n5736), .B2(n4729), .ZN(n1508)
         );
  OAI222_X1 U2824 ( .A1(n5731), .A2(n4665), .B1(n5737), .B2(n4633), .C1(n5732), 
        .C2(n4697), .ZN(n1507) );
  AOI221_X1 U2825 ( .B1(n1282), .B2(n1509), .C1(n1284), .C2(n1510), .A(n1511), 
        .ZN(n1496) );
  OAI22_X1 U2826 ( .A1(n4473), .A2(n1287), .B1(n5305), .B2(n1288), .ZN(n1511)
         );
  INV_X1 U2827 ( .A(n5081), .ZN(n1509) );
  AOI222_X1 U2828 ( .A1(n1512), .A2(n1290), .B1(n1291), .B2(n1513), .C1(n1514), 
        .C2(n1294), .ZN(n1495) );
  AND4_X1 U2829 ( .A1(n1515), .A2(n1516), .A3(n1517), .A4(n1518), .ZN(n5490)
         );
  NOR4_X1 U2830 ( .A1(n1519), .A2(n1520), .A3(n1521), .A4(n1522), .ZN(n1518)
         );
  NAND3_X1 U2831 ( .A1(n5916), .A2(n5915), .A3(n5917), .ZN(n1522) );
  OAI211_X1 U2832 ( .C1(n5745), .C2(n5400), .A(n5913), .B(n5914), .ZN(n1521)
         );
  OAI222_X1 U2833 ( .A1(n5743), .A2(n5272), .B1(n5744), .B2(n5240), .C1(n5746), 
        .C2(n5368), .ZN(n1520) );
  OAI221_X1 U2834 ( .B1(n5716), .B2(n5176), .C1(n5717), .C2(n5208), .A(n1523), 
        .ZN(n1519) );
  AOI22_X1 U2835 ( .A1(n1524), .A2(n1275), .B1(n1525), .B2(n1277), .ZN(n1523)
         );
  AOI211_X1 U2836 ( .C1(n1526), .C2(n1279), .A(n1527), .B(n1528), .ZN(n1517)
         );
  OAI22_X1 U2837 ( .A1(n5726), .A2(n4824), .B1(n5736), .B2(n4728), .ZN(n1528)
         );
  OAI222_X1 U2838 ( .A1(n5731), .A2(n4664), .B1(n5737), .B2(n4632), .C1(n5732), 
        .C2(n4696), .ZN(n1527) );
  AOI221_X1 U2839 ( .B1(n1282), .B2(n1529), .C1(n1284), .C2(n1530), .A(n1531), 
        .ZN(n1516) );
  OAI22_X1 U2840 ( .A1(n4472), .A2(n1287), .B1(n5304), .B2(n1288), .ZN(n1531)
         );
  INV_X1 U2841 ( .A(n5080), .ZN(n1529) );
  AOI222_X1 U2842 ( .A1(n1532), .A2(n1290), .B1(n1291), .B2(n1533), .C1(n1534), 
        .C2(n1294), .ZN(n1515) );
  AND4_X1 U2843 ( .A1(n1535), .A2(n1536), .A3(n1537), .A4(n1538), .ZN(n5487)
         );
  NOR4_X1 U2844 ( .A1(n1539), .A2(n1540), .A3(n1541), .A4(n1542), .ZN(n1538)
         );
  NAND3_X1 U2845 ( .A1(n5911), .A2(n5910), .A3(n5912), .ZN(n1542) );
  OAI211_X1 U2846 ( .C1(n5745), .C2(n5399), .A(n5908), .B(n5909), .ZN(n1541)
         );
  OAI222_X1 U2847 ( .A1(n5743), .A2(n5271), .B1(n5744), .B2(n5239), .C1(n5746), 
        .C2(n5367), .ZN(n1540) );
  OAI221_X1 U2848 ( .B1(n5716), .B2(n5175), .C1(n5717), .C2(n5207), .A(n1543), 
        .ZN(n1539) );
  AOI22_X1 U2849 ( .A1(n1544), .A2(n1275), .B1(n1545), .B2(n1277), .ZN(n1543)
         );
  AOI211_X1 U2850 ( .C1(n1546), .C2(n1279), .A(n1547), .B(n1548), .ZN(n1537)
         );
  OAI22_X1 U2851 ( .A1(n5726), .A2(n4823), .B1(n5736), .B2(n4727), .ZN(n1548)
         );
  OAI222_X1 U2852 ( .A1(n5731), .A2(n4663), .B1(n5737), .B2(n4631), .C1(n5732), 
        .C2(n4695), .ZN(n1547) );
  AOI221_X1 U2853 ( .B1(n1282), .B2(n1549), .C1(n1284), .C2(n1550), .A(n1551), 
        .ZN(n1536) );
  OAI22_X1 U2854 ( .A1(n4471), .A2(n1287), .B1(n5303), .B2(n1288), .ZN(n1551)
         );
  INV_X1 U2855 ( .A(n5079), .ZN(n1549) );
  AOI222_X1 U2856 ( .A1(n1552), .A2(n1290), .B1(n1291), .B2(n1553), .C1(n1554), 
        .C2(n1294), .ZN(n1535) );
  AND4_X1 U2857 ( .A1(n1555), .A2(n1556), .A3(n1557), .A4(n1558), .ZN(n5484)
         );
  NOR4_X1 U2858 ( .A1(n1559), .A2(n1560), .A3(n1561), .A4(n1562), .ZN(n1558)
         );
  NAND3_X1 U2859 ( .A1(n5906), .A2(n5905), .A3(n5907), .ZN(n1562) );
  OAI211_X1 U2860 ( .C1(n5745), .C2(n5398), .A(n5903), .B(n5904), .ZN(n1561)
         );
  OAI222_X1 U2861 ( .A1(n5743), .A2(n5270), .B1(n5744), .B2(n5238), .C1(n5746), 
        .C2(n5366), .ZN(n1560) );
  OAI221_X1 U2862 ( .B1(n5716), .B2(n5174), .C1(n5717), .C2(n5206), .A(n1563), 
        .ZN(n1559) );
  AOI22_X1 U2863 ( .A1(n1564), .A2(n1275), .B1(n1565), .B2(n1277), .ZN(n1563)
         );
  AOI211_X1 U2864 ( .C1(n1566), .C2(n1279), .A(n1567), .B(n1568), .ZN(n1557)
         );
  OAI22_X1 U2865 ( .A1(n5726), .A2(n4822), .B1(n5736), .B2(n4726), .ZN(n1568)
         );
  OAI222_X1 U2866 ( .A1(n5731), .A2(n4662), .B1(n5737), .B2(n4630), .C1(n5732), 
        .C2(n4694), .ZN(n1567) );
  AOI221_X1 U2867 ( .B1(n1282), .B2(n1569), .C1(n1284), .C2(n1570), .A(n1571), 
        .ZN(n1556) );
  OAI22_X1 U2868 ( .A1(n4470), .A2(n1287), .B1(n5302), .B2(n1288), .ZN(n1571)
         );
  INV_X1 U2869 ( .A(n5078), .ZN(n1569) );
  AOI222_X1 U2870 ( .A1(n1572), .A2(n1290), .B1(n1291), .B2(n1573), .C1(n1574), 
        .C2(n1294), .ZN(n1555) );
  AND4_X1 U2871 ( .A1(n1575), .A2(n1576), .A3(n1577), .A4(n1578), .ZN(n5481)
         );
  NOR4_X1 U2872 ( .A1(n1579), .A2(n1580), .A3(n1581), .A4(n1582), .ZN(n1578)
         );
  NAND3_X1 U2873 ( .A1(n5901), .A2(n5900), .A3(n5902), .ZN(n1582) );
  OAI211_X1 U2874 ( .C1(n5745), .C2(n5397), .A(n5898), .B(n5899), .ZN(n1581)
         );
  OAI222_X1 U2875 ( .A1(n5743), .A2(n5269), .B1(n5744), .B2(n5237), .C1(n5746), 
        .C2(n5365), .ZN(n1580) );
  OAI221_X1 U2876 ( .B1(n5716), .B2(n5173), .C1(n5717), .C2(n5205), .A(n1583), 
        .ZN(n1579) );
  AOI22_X1 U2877 ( .A1(n1584), .A2(n1275), .B1(n1585), .B2(n1277), .ZN(n1583)
         );
  AOI211_X1 U2878 ( .C1(n1586), .C2(n1279), .A(n1587), .B(n1588), .ZN(n1577)
         );
  OAI22_X1 U2879 ( .A1(n5726), .A2(n4821), .B1(n5736), .B2(n4725), .ZN(n1588)
         );
  OAI222_X1 U2880 ( .A1(n5731), .A2(n4661), .B1(n5737), .B2(n4629), .C1(n5732), 
        .C2(n4693), .ZN(n1587) );
  AOI221_X1 U2881 ( .B1(n1282), .B2(n1589), .C1(n1284), .C2(n1590), .A(n1591), 
        .ZN(n1576) );
  OAI22_X1 U2882 ( .A1(n4469), .A2(n1287), .B1(n5301), .B2(n1288), .ZN(n1591)
         );
  INV_X1 U2883 ( .A(n5077), .ZN(n1589) );
  AOI222_X1 U2884 ( .A1(n1592), .A2(n1290), .B1(n1291), .B2(n1593), .C1(n1594), 
        .C2(n1294), .ZN(n1575) );
  AND4_X1 U2885 ( .A1(n1595), .A2(n1596), .A3(n1597), .A4(n1598), .ZN(n5478)
         );
  NOR4_X1 U2886 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .ZN(n1598)
         );
  NAND3_X1 U2887 ( .A1(n5894), .A2(n5893), .A3(n5895), .ZN(n1602) );
  OAI211_X1 U2888 ( .C1(n5745), .C2(n5396), .A(n5891), .B(n5892), .ZN(n1601)
         );
  OAI222_X1 U2889 ( .A1(n5743), .A2(n5268), .B1(n5744), .B2(n5236), .C1(n5746), 
        .C2(n5364), .ZN(n1600) );
  OAI221_X1 U2890 ( .B1(n5716), .B2(n5172), .C1(n5717), .C2(n5204), .A(n1603), 
        .ZN(n1599) );
  AOI22_X1 U2891 ( .A1(n1604), .A2(n1275), .B1(n1605), .B2(n1277), .ZN(n1603)
         );
  AOI211_X1 U2892 ( .C1(n1606), .C2(n1279), .A(n1607), .B(n1608), .ZN(n1597)
         );
  OAI22_X1 U2893 ( .A1(n5726), .A2(n4820), .B1(n5736), .B2(n4724), .ZN(n1608)
         );
  OAI222_X1 U2894 ( .A1(n5731), .A2(n4660), .B1(n5737), .B2(n4628), .C1(n5732), 
        .C2(n4692), .ZN(n1607) );
  AOI221_X1 U2895 ( .B1(n1282), .B2(n1609), .C1(n1284), .C2(n1610), .A(n1611), 
        .ZN(n1596) );
  OAI22_X1 U2896 ( .A1(n4468), .A2(n1287), .B1(n5300), .B2(n1288), .ZN(n1611)
         );
  INV_X1 U2897 ( .A(n5076), .ZN(n1609) );
  AOI222_X1 U2898 ( .A1(n1612), .A2(n1290), .B1(n1291), .B2(n1613), .C1(n1614), 
        .C2(n1294), .ZN(n1595) );
  AND4_X1 U2899 ( .A1(n1615), .A2(n1616), .A3(n1617), .A4(n1618), .ZN(n5475)
         );
  NOR4_X1 U2900 ( .A1(n1619), .A2(n1620), .A3(n1621), .A4(n1622), .ZN(n1618)
         );
  NAND3_X1 U2901 ( .A1(n5886), .A2(n5885), .A3(n5887), .ZN(n1622) );
  OAI211_X1 U2902 ( .C1(n5745), .C2(n5395), .A(n5883), .B(n5884), .ZN(n1621)
         );
  OAI222_X1 U2903 ( .A1(n5743), .A2(n5267), .B1(n5744), .B2(n5235), .C1(n5746), 
        .C2(n5363), .ZN(n1620) );
  OAI221_X1 U2904 ( .B1(n5716), .B2(n5171), .C1(n5717), .C2(n5203), .A(n1623), 
        .ZN(n1619) );
  AOI22_X1 U2905 ( .A1(n1624), .A2(n1275), .B1(n1625), .B2(n1277), .ZN(n1623)
         );
  AOI211_X1 U2906 ( .C1(n1626), .C2(n1279), .A(n1627), .B(n1628), .ZN(n1617)
         );
  OAI22_X1 U2907 ( .A1(n5726), .A2(n4819), .B1(n5736), .B2(n4723), .ZN(n1628)
         );
  OAI222_X1 U2908 ( .A1(n5731), .A2(n4659), .B1(n5737), .B2(n4627), .C1(n5732), 
        .C2(n4691), .ZN(n1627) );
  AOI221_X1 U2909 ( .B1(n1282), .B2(n1629), .C1(n1284), .C2(n1630), .A(n1631), 
        .ZN(n1616) );
  OAI22_X1 U2910 ( .A1(n4467), .A2(n1287), .B1(n5299), .B2(n1288), .ZN(n1631)
         );
  INV_X1 U2911 ( .A(n5075), .ZN(n1629) );
  AOI222_X1 U2912 ( .A1(n1632), .A2(n1290), .B1(n1291), .B2(n1633), .C1(n1634), 
        .C2(n1294), .ZN(n1615) );
  AND4_X1 U2913 ( .A1(n1635), .A2(n1636), .A3(n1637), .A4(n1638), .ZN(n5472)
         );
  NOR4_X1 U2914 ( .A1(n1639), .A2(n1640), .A3(n1641), .A4(n1642), .ZN(n1638)
         );
  NAND3_X1 U2915 ( .A1(n5877), .A2(n5876), .A3(n5878), .ZN(n1642) );
  OAI211_X1 U2916 ( .C1(n5745), .C2(n5394), .A(n5874), .B(n5875), .ZN(n1641)
         );
  OAI222_X1 U2917 ( .A1(n5743), .A2(n5266), .B1(n5744), .B2(n5234), .C1(n5746), 
        .C2(n5362), .ZN(n1640) );
  OAI221_X1 U2918 ( .B1(n5716), .B2(n5170), .C1(n5717), .C2(n5202), .A(n1643), 
        .ZN(n1639) );
  AOI22_X1 U2919 ( .A1(n1644), .A2(n1275), .B1(n1645), .B2(n1277), .ZN(n1643)
         );
  AOI211_X1 U2920 ( .C1(n1646), .C2(n1279), .A(n1647), .B(n1648), .ZN(n1637)
         );
  OAI22_X1 U2921 ( .A1(n5726), .A2(n4818), .B1(n5736), .B2(n4722), .ZN(n1648)
         );
  OAI222_X1 U2922 ( .A1(n5731), .A2(n4658), .B1(n5737), .B2(n4626), .C1(n5732), 
        .C2(n4690), .ZN(n1647) );
  AOI221_X1 U2923 ( .B1(n1282), .B2(n1649), .C1(n1284), .C2(n1650), .A(n1651), 
        .ZN(n1636) );
  OAI22_X1 U2924 ( .A1(n4466), .A2(n1287), .B1(n5298), .B2(n1288), .ZN(n1651)
         );
  INV_X1 U2925 ( .A(n5074), .ZN(n1649) );
  AOI222_X1 U2926 ( .A1(n1652), .A2(n1290), .B1(n1291), .B2(n1653), .C1(n1654), 
        .C2(n1294), .ZN(n1635) );
  AND4_X1 U2927 ( .A1(n1655), .A2(n1656), .A3(n1657), .A4(n1658), .ZN(n5469)
         );
  NOR4_X1 U2928 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1658)
         );
  NAND3_X1 U2929 ( .A1(n5867), .A2(n5866), .A3(n5868), .ZN(n1662) );
  OAI211_X1 U2930 ( .C1(n5745), .C2(n5393), .A(n5864), .B(n5865), .ZN(n1661)
         );
  OAI222_X1 U2931 ( .A1(n5743), .A2(n5265), .B1(n5744), .B2(n5233), .C1(n5746), 
        .C2(n5361), .ZN(n1660) );
  OAI221_X1 U2932 ( .B1(n5716), .B2(n5169), .C1(n5717), .C2(n5201), .A(n1663), 
        .ZN(n1659) );
  AOI22_X1 U2933 ( .A1(n1664), .A2(n1275), .B1(n1665), .B2(n1277), .ZN(n1663)
         );
  AOI211_X1 U2934 ( .C1(n1666), .C2(n1279), .A(n1667), .B(n1668), .ZN(n1657)
         );
  OAI22_X1 U2935 ( .A1(n5726), .A2(n4817), .B1(n5736), .B2(n4721), .ZN(n1668)
         );
  OAI222_X1 U2936 ( .A1(n5731), .A2(n4657), .B1(n5737), .B2(n4625), .C1(n5732), 
        .C2(n4689), .ZN(n1667) );
  AOI221_X1 U2937 ( .B1(n1282), .B2(n1669), .C1(n1284), .C2(n1670), .A(n1671), 
        .ZN(n1656) );
  OAI22_X1 U2938 ( .A1(n4465), .A2(n1287), .B1(n5297), .B2(n1288), .ZN(n1671)
         );
  INV_X1 U2939 ( .A(n5073), .ZN(n1669) );
  AOI222_X1 U2940 ( .A1(n1672), .A2(n1290), .B1(n1291), .B2(n1673), .C1(n1674), 
        .C2(n1294), .ZN(n1655) );
  AND4_X1 U2941 ( .A1(n1675), .A2(n1676), .A3(n1677), .A4(n1678), .ZN(n5466)
         );
  NOR4_X1 U2942 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .ZN(n1678)
         );
  NAND3_X1 U2943 ( .A1(n5861), .A2(n5860), .A3(n5862), .ZN(n1682) );
  OAI211_X1 U2944 ( .C1(n5745), .C2(n5392), .A(n5858), .B(n5859), .ZN(n1681)
         );
  OAI222_X1 U2945 ( .A1(n5743), .A2(n5264), .B1(n5744), .B2(n5232), .C1(n5746), 
        .C2(n5360), .ZN(n1680) );
  OAI221_X1 U2946 ( .B1(n5716), .B2(n5168), .C1(n5717), .C2(n5200), .A(n1683), 
        .ZN(n1679) );
  AOI22_X1 U2947 ( .A1(n1684), .A2(n1275), .B1(n1685), .B2(n1277), .ZN(n1683)
         );
  AOI211_X1 U2948 ( .C1(n1686), .C2(n1279), .A(n1687), .B(n1688), .ZN(n1677)
         );
  OAI22_X1 U2949 ( .A1(n5726), .A2(n4816), .B1(n5736), .B2(n4720), .ZN(n1688)
         );
  OAI222_X1 U2950 ( .A1(n5731), .A2(n4656), .B1(n5737), .B2(n4624), .C1(n5732), 
        .C2(n4688), .ZN(n1687) );
  AOI221_X1 U2951 ( .B1(n1282), .B2(n1689), .C1(n1284), .C2(n1690), .A(n1691), 
        .ZN(n1676) );
  OAI22_X1 U2952 ( .A1(n4464), .A2(n1287), .B1(n5296), .B2(n1288), .ZN(n1691)
         );
  INV_X1 U2953 ( .A(n5072), .ZN(n1689) );
  AOI222_X1 U2954 ( .A1(n1692), .A2(n1290), .B1(n1291), .B2(n1693), .C1(n1694), 
        .C2(n1294), .ZN(n1675) );
  AND4_X1 U2955 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n5463)
         );
  NOR4_X1 U2956 ( .A1(n1699), .A2(n1700), .A3(n1701), .A4(n1702), .ZN(n1698)
         );
  NAND3_X1 U2957 ( .A1(n5855), .A2(n5854), .A3(n5856), .ZN(n1702) );
  OAI211_X1 U2958 ( .C1(n5745), .C2(n5391), .A(n5852), .B(n5853), .ZN(n1701)
         );
  OAI222_X1 U2959 ( .A1(n5743), .A2(n5263), .B1(n5744), .B2(n5231), .C1(n5746), 
        .C2(n5359), .ZN(n1700) );
  OAI221_X1 U2960 ( .B1(n5716), .B2(n5167), .C1(n5717), .C2(n5199), .A(n1703), 
        .ZN(n1699) );
  AOI22_X1 U2961 ( .A1(n1704), .A2(n1275), .B1(n1705), .B2(n1277), .ZN(n1703)
         );
  AOI211_X1 U2962 ( .C1(n1706), .C2(n1279), .A(n1707), .B(n1708), .ZN(n1697)
         );
  OAI22_X1 U2963 ( .A1(n5726), .A2(n4815), .B1(n5736), .B2(n4719), .ZN(n1708)
         );
  OAI222_X1 U2964 ( .A1(n5731), .A2(n4655), .B1(n5737), .B2(n4623), .C1(n5732), 
        .C2(n4687), .ZN(n1707) );
  AOI221_X1 U2965 ( .B1(n1282), .B2(n1709), .C1(n1284), .C2(n1710), .A(n1711), 
        .ZN(n1696) );
  OAI22_X1 U2966 ( .A1(n4463), .A2(n1287), .B1(n5295), .B2(n1288), .ZN(n1711)
         );
  INV_X1 U2967 ( .A(n5071), .ZN(n1709) );
  AOI222_X1 U2968 ( .A1(n1712), .A2(n1290), .B1(n1291), .B2(n1713), .C1(n1714), 
        .C2(n1294), .ZN(n1695) );
  AND4_X1 U2969 ( .A1(n1715), .A2(n1716), .A3(n1717), .A4(n1718), .ZN(n5460)
         );
  NOR4_X1 U2970 ( .A1(n1719), .A2(n1720), .A3(n1721), .A4(n1722), .ZN(n1718)
         );
  NAND3_X1 U2971 ( .A1(n5849), .A2(n5848), .A3(n5850), .ZN(n1722) );
  OAI211_X1 U2972 ( .C1(n5745), .C2(n5390), .A(n5846), .B(n5847), .ZN(n1721)
         );
  OAI222_X1 U2973 ( .A1(n5743), .A2(n5262), .B1(n5744), .B2(n5230), .C1(n5746), 
        .C2(n5358), .ZN(n1720) );
  OAI221_X1 U2974 ( .B1(n5716), .B2(n5166), .C1(n5717), .C2(n5198), .A(n1723), 
        .ZN(n1719) );
  AOI22_X1 U2975 ( .A1(n1724), .A2(n1275), .B1(n1725), .B2(n1277), .ZN(n1723)
         );
  AOI211_X1 U2976 ( .C1(n1726), .C2(n1279), .A(n1727), .B(n1728), .ZN(n1717)
         );
  OAI22_X1 U2977 ( .A1(n5726), .A2(n4814), .B1(n5736), .B2(n4718), .ZN(n1728)
         );
  OAI222_X1 U2978 ( .A1(n5731), .A2(n4654), .B1(n5737), .B2(n4622), .C1(n5732), 
        .C2(n4686), .ZN(n1727) );
  AOI221_X1 U2979 ( .B1(n1282), .B2(n1729), .C1(n1284), .C2(n1730), .A(n1731), 
        .ZN(n1716) );
  OAI22_X1 U2980 ( .A1(n4462), .A2(n1287), .B1(n5294), .B2(n1288), .ZN(n1731)
         );
  INV_X1 U2981 ( .A(n5070), .ZN(n1729) );
  AOI222_X1 U2982 ( .A1(n1732), .A2(n1290), .B1(n1291), .B2(n1733), .C1(n1734), 
        .C2(n1294), .ZN(n1715) );
  AND4_X1 U2983 ( .A1(n1735), .A2(n1736), .A3(n1737), .A4(n1738), .ZN(n5457)
         );
  NOR4_X1 U2984 ( .A1(n1739), .A2(n1740), .A3(n1741), .A4(n1742), .ZN(n1738)
         );
  NAND3_X1 U2985 ( .A1(n5836), .A2(n5835), .A3(n5837), .ZN(n1742) );
  OAI211_X1 U2986 ( .C1(n5745), .C2(n5389), .A(n5833), .B(n5834), .ZN(n1741)
         );
  OAI222_X1 U2987 ( .A1(n5743), .A2(n5261), .B1(n5744), .B2(n5229), .C1(n5746), 
        .C2(n5357), .ZN(n1740) );
  OAI221_X1 U2988 ( .B1(n5716), .B2(n5165), .C1(n5717), .C2(n5197), .A(n1743), 
        .ZN(n1739) );
  AOI22_X1 U2989 ( .A1(n1744), .A2(n1275), .B1(n1745), .B2(n1277), .ZN(n1743)
         );
  AOI211_X1 U2990 ( .C1(n1746), .C2(n1279), .A(n1747), .B(n1748), .ZN(n1737)
         );
  OAI22_X1 U2991 ( .A1(n5726), .A2(n4813), .B1(n5736), .B2(n4717), .ZN(n1748)
         );
  OAI222_X1 U2992 ( .A1(n5731), .A2(n4653), .B1(n5737), .B2(n4621), .C1(n5732), 
        .C2(n4685), .ZN(n1747) );
  AOI221_X1 U2993 ( .B1(n1282), .B2(n1749), .C1(n1284), .C2(n1750), .A(n1751), 
        .ZN(n1736) );
  OAI22_X1 U2994 ( .A1(n4461), .A2(n1287), .B1(n5293), .B2(n1288), .ZN(n1751)
         );
  INV_X1 U2995 ( .A(n5069), .ZN(n1749) );
  AOI222_X1 U2996 ( .A1(n1752), .A2(n1290), .B1(n1291), .B2(n1753), .C1(n1754), 
        .C2(n1294), .ZN(n1735) );
  AND4_X1 U2997 ( .A1(n1755), .A2(n1756), .A3(n1757), .A4(n1758), .ZN(n5454)
         );
  NOR4_X1 U2998 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(n1758)
         );
  NAND3_X1 U2999 ( .A1(n5829), .A2(n5828), .A3(n5830), .ZN(n1762) );
  OAI211_X1 U3000 ( .C1(n5745), .C2(n5388), .A(n5826), .B(n5827), .ZN(n1761)
         );
  OAI222_X1 U3001 ( .A1(n5743), .A2(n5260), .B1(n5744), .B2(n5228), .C1(n5746), 
        .C2(n5356), .ZN(n1760) );
  OAI221_X1 U3002 ( .B1(n5716), .B2(n5164), .C1(n5717), .C2(n5196), .A(n1763), 
        .ZN(n1759) );
  AOI22_X1 U3003 ( .A1(n1764), .A2(n1275), .B1(n1765), .B2(n1277), .ZN(n1763)
         );
  AOI211_X1 U3004 ( .C1(n1766), .C2(n1279), .A(n1767), .B(n1768), .ZN(n1757)
         );
  OAI22_X1 U3005 ( .A1(n5726), .A2(n4812), .B1(n5736), .B2(n4716), .ZN(n1768)
         );
  OAI222_X1 U3006 ( .A1(n5731), .A2(n4652), .B1(n5737), .B2(n4620), .C1(n5732), 
        .C2(n4684), .ZN(n1767) );
  AOI221_X1 U3007 ( .B1(n1282), .B2(n1769), .C1(n1284), .C2(n1770), .A(n1771), 
        .ZN(n1756) );
  OAI22_X1 U3008 ( .A1(n4460), .A2(n1287), .B1(n5292), .B2(n1288), .ZN(n1771)
         );
  INV_X1 U3009 ( .A(n5068), .ZN(n1769) );
  AOI222_X1 U3010 ( .A1(n1772), .A2(n1290), .B1(n1291), .B2(n1773), .C1(n1774), 
        .C2(n1294), .ZN(n1755) );
  AND4_X1 U3011 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .ZN(n5451)
         );
  NOR4_X1 U3012 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .ZN(n1778)
         );
  NAND3_X1 U3013 ( .A1(n5823), .A2(n5822), .A3(n5824), .ZN(n1782) );
  OAI211_X1 U3014 ( .C1(n5745), .C2(n5387), .A(n5820), .B(n5821), .ZN(n1781)
         );
  OAI222_X1 U3015 ( .A1(n5743), .A2(n5259), .B1(n5744), .B2(n5227), .C1(n5746), 
        .C2(n5355), .ZN(n1780) );
  OAI221_X1 U3016 ( .B1(n5716), .B2(n5163), .C1(n5717), .C2(n5195), .A(n1783), 
        .ZN(n1779) );
  AOI22_X1 U3017 ( .A1(n1784), .A2(n1275), .B1(n1785), .B2(n1277), .ZN(n1783)
         );
  AOI211_X1 U3018 ( .C1(n1786), .C2(n1279), .A(n1787), .B(n1788), .ZN(n1777)
         );
  OAI22_X1 U3019 ( .A1(n5726), .A2(n4811), .B1(n5736), .B2(n4715), .ZN(n1788)
         );
  OAI222_X1 U3020 ( .A1(n5731), .A2(n4651), .B1(n5737), .B2(n4619), .C1(n5732), 
        .C2(n4683), .ZN(n1787) );
  AOI221_X1 U3021 ( .B1(n1282), .B2(n1789), .C1(n1284), .C2(n1790), .A(n1791), 
        .ZN(n1776) );
  OAI22_X1 U3022 ( .A1(n4459), .A2(n1287), .B1(n5291), .B2(n1288), .ZN(n1791)
         );
  INV_X1 U3023 ( .A(n5067), .ZN(n1789) );
  AOI222_X1 U3024 ( .A1(n1792), .A2(n1290), .B1(n1291), .B2(n1793), .C1(n1794), 
        .C2(n1294), .ZN(n1775) );
  AND4_X1 U3025 ( .A1(n1795), .A2(n1796), .A3(n1797), .A4(n1798), .ZN(n5448)
         );
  NOR4_X1 U3026 ( .A1(n1799), .A2(n1800), .A3(n1801), .A4(n1802), .ZN(n1798)
         );
  NAND3_X1 U3027 ( .A1(n5810), .A2(n5809), .A3(n5811), .ZN(n1802) );
  OAI211_X1 U3028 ( .C1(n5745), .C2(n5386), .A(n5807), .B(n5808), .ZN(n1801)
         );
  OAI222_X1 U3029 ( .A1(n5743), .A2(n5258), .B1(n5744), .B2(n5226), .C1(n5746), 
        .C2(n5354), .ZN(n1800) );
  OAI221_X1 U3030 ( .B1(n5716), .B2(n5162), .C1(n5717), .C2(n5194), .A(n1803), 
        .ZN(n1799) );
  AOI22_X1 U3031 ( .A1(n1804), .A2(n1275), .B1(n1805), .B2(n1277), .ZN(n1803)
         );
  AOI211_X1 U3032 ( .C1(n1806), .C2(n1279), .A(n1807), .B(n1808), .ZN(n1797)
         );
  OAI22_X1 U3033 ( .A1(n5726), .A2(n4810), .B1(n5736), .B2(n4714), .ZN(n1808)
         );
  OAI222_X1 U3034 ( .A1(n5731), .A2(n4650), .B1(n5737), .B2(n4618), .C1(n5732), 
        .C2(n4682), .ZN(n1807) );
  AOI221_X1 U3035 ( .B1(n1282), .B2(n1809), .C1(n1284), .C2(n1810), .A(n1811), 
        .ZN(n1796) );
  OAI22_X1 U3036 ( .A1(n4458), .A2(n1287), .B1(n5290), .B2(n1288), .ZN(n1811)
         );
  INV_X1 U3037 ( .A(n5066), .ZN(n1809) );
  AOI222_X1 U3038 ( .A1(n1812), .A2(n1290), .B1(n1291), .B2(n1813), .C1(n1814), 
        .C2(n1294), .ZN(n1795) );
  AND4_X1 U3039 ( .A1(n1815), .A2(n1816), .A3(n1817), .A4(n1818), .ZN(n5445)
         );
  NOR4_X1 U3040 ( .A1(n1819), .A2(n1820), .A3(n1821), .A4(n1822), .ZN(n1818)
         );
  NAND3_X1 U3041 ( .A1(n5797), .A2(n5796), .A3(n5798), .ZN(n1822) );
  OAI211_X1 U3042 ( .C1(n5745), .C2(n5385), .A(n5794), .B(n5795), .ZN(n1821)
         );
  OAI222_X1 U3043 ( .A1(n5743), .A2(n5257), .B1(n5744), .B2(n5225), .C1(n5746), 
        .C2(n5353), .ZN(n1820) );
  OAI221_X1 U3044 ( .B1(n5716), .B2(n5161), .C1(n5717), .C2(n5193), .A(n1823), 
        .ZN(n1819) );
  AOI22_X1 U3045 ( .A1(n1824), .A2(n1275), .B1(n1825), .B2(n1277), .ZN(n1823)
         );
  AOI211_X1 U3046 ( .C1(n1826), .C2(n1279), .A(n1827), .B(n1828), .ZN(n1817)
         );
  OAI22_X1 U3047 ( .A1(n5726), .A2(n4809), .B1(n5736), .B2(n4713), .ZN(n1828)
         );
  OAI222_X1 U3048 ( .A1(n5731), .A2(n4649), .B1(n5737), .B2(n4617), .C1(n5732), 
        .C2(n4681), .ZN(n1827) );
  AOI221_X1 U3049 ( .B1(n1282), .B2(n1829), .C1(n1284), .C2(n1830), .A(n1831), 
        .ZN(n1816) );
  OAI22_X1 U3050 ( .A1(n4457), .A2(n1287), .B1(n5289), .B2(n1288), .ZN(n1831)
         );
  INV_X1 U3051 ( .A(n5065), .ZN(n1829) );
  AOI222_X1 U3052 ( .A1(n1832), .A2(n1290), .B1(n1291), .B2(n1833), .C1(n1834), 
        .C2(n1294), .ZN(n1815) );
  AND4_X1 U3053 ( .A1(n1835), .A2(n1836), .A3(n1837), .A4(n1838), .ZN(n5442)
         );
  NOR4_X1 U3054 ( .A1(n1839), .A2(n1840), .A3(n1841), .A4(n1842), .ZN(n1838)
         );
  NAND3_X1 U3055 ( .A1(n5784), .A2(n5783), .A3(n5785), .ZN(n1842) );
  OAI211_X1 U3056 ( .C1(n5745), .C2(n5384), .A(n5781), .B(n5782), .ZN(n1841)
         );
  OAI222_X1 U3057 ( .A1(n5743), .A2(n5256), .B1(n5744), .B2(n5224), .C1(n5746), 
        .C2(n5352), .ZN(n1840) );
  OAI221_X1 U3058 ( .B1(n5716), .B2(n5160), .C1(n5717), .C2(n5192), .A(n1843), 
        .ZN(n1839) );
  AOI22_X1 U3059 ( .A1(n1844), .A2(n1275), .B1(n1845), .B2(n1277), .ZN(n1843)
         );
  AOI211_X1 U3060 ( .C1(n1846), .C2(n1279), .A(n1847), .B(n1848), .ZN(n1837)
         );
  OAI22_X1 U3061 ( .A1(n5726), .A2(n4808), .B1(n5736), .B2(n4712), .ZN(n1848)
         );
  OAI222_X1 U3062 ( .A1(n5731), .A2(n4648), .B1(n5737), .B2(n4616), .C1(n5732), 
        .C2(n4680), .ZN(n1847) );
  AOI221_X1 U3063 ( .B1(n1282), .B2(n1849), .C1(n1284), .C2(n1850), .A(n1851), 
        .ZN(n1836) );
  OAI22_X1 U3064 ( .A1(n4456), .A2(n1287), .B1(n5288), .B2(n1288), .ZN(n1851)
         );
  INV_X1 U3065 ( .A(n5064), .ZN(n1849) );
  AOI222_X1 U3066 ( .A1(n1852), .A2(n1290), .B1(n1291), .B2(n1853), .C1(n1854), 
        .C2(n1294), .ZN(n1835) );
  AND4_X1 U3067 ( .A1(n1855), .A2(n1856), .A3(n1857), .A4(n1858), .ZN(n5439)
         );
  NOR4_X1 U3068 ( .A1(n1859), .A2(n1860), .A3(n1861), .A4(n1862), .ZN(n1858)
         );
  NAND3_X1 U3069 ( .A1(n5767), .A2(n5766), .A3(n5768), .ZN(n1862) );
  OAI211_X1 U3070 ( .C1(n5745), .C2(n5383), .A(n5764), .B(n5765), .ZN(n1861)
         );
  OAI222_X1 U3071 ( .A1(n5743), .A2(n5255), .B1(n5744), .B2(n5223), .C1(n5746), 
        .C2(n5351), .ZN(n1860) );
  OAI221_X1 U3072 ( .B1(n5716), .B2(n5159), .C1(n5717), .C2(n5191), .A(n1863), 
        .ZN(n1859) );
  AOI22_X1 U3073 ( .A1(n1864), .A2(n1275), .B1(n1865), .B2(n1277), .ZN(n1863)
         );
  AOI211_X1 U3074 ( .C1(n1866), .C2(n1279), .A(n1867), .B(n1868), .ZN(n1857)
         );
  OAI22_X1 U3075 ( .A1(n5726), .A2(n4807), .B1(n5736), .B2(n4711), .ZN(n1868)
         );
  OAI222_X1 U3076 ( .A1(n5731), .A2(n4647), .B1(n5737), .B2(n4615), .C1(n5732), 
        .C2(n4679), .ZN(n1867) );
  AOI221_X1 U3077 ( .B1(n1282), .B2(n1869), .C1(n1284), .C2(n1870), .A(n1871), 
        .ZN(n1856) );
  OAI22_X1 U3078 ( .A1(n4455), .A2(n1287), .B1(n5287), .B2(n1288), .ZN(n1871)
         );
  INV_X1 U3079 ( .A(n5063), .ZN(n1869) );
  AOI222_X1 U3080 ( .A1(n1872), .A2(n1290), .B1(n1291), .B2(n1873), .C1(n1874), 
        .C2(n1294), .ZN(n1855) );
  AND4_X1 U3081 ( .A1(n1875), .A2(n1876), .A3(n1877), .A4(n1878), .ZN(n5436)
         );
  NOR4_X1 U3082 ( .A1(n1879), .A2(n1880), .A3(n1881), .A4(n1882), .ZN(n1878)
         );
  NAND3_X1 U3083 ( .A1(n5752), .A2(n5751), .A3(n5753), .ZN(n1882) );
  OAI211_X1 U3084 ( .C1(n5745), .C2(n5382), .A(n5749), .B(n5750), .ZN(n1881)
         );
  OAI222_X1 U3085 ( .A1(n5743), .A2(n5254), .B1(n5744), .B2(n5222), .C1(n5746), 
        .C2(n5350), .ZN(n1880) );
  OAI221_X1 U3086 ( .B1(n5716), .B2(n5158), .C1(n5717), .C2(n5190), .A(n1883), 
        .ZN(n1879) );
  AOI22_X1 U3087 ( .A1(n1884), .A2(n1275), .B1(n1885), .B2(n1277), .ZN(n1883)
         );
  AOI211_X1 U3088 ( .C1(n1886), .C2(n1279), .A(n1887), .B(n1888), .ZN(n1877)
         );
  OAI22_X1 U3089 ( .A1(n5726), .A2(n4806), .B1(n5736), .B2(n4710), .ZN(n1888)
         );
  OAI222_X1 U3090 ( .A1(n5731), .A2(n4646), .B1(n5737), .B2(n4614), .C1(n5732), 
        .C2(n4678), .ZN(n1887) );
  AOI221_X1 U3091 ( .B1(n1282), .B2(n1889), .C1(n1284), .C2(n1890), .A(n1891), 
        .ZN(n1876) );
  OAI22_X1 U3092 ( .A1(n4454), .A2(n1287), .B1(n5286), .B2(n1288), .ZN(n1891)
         );
  INV_X1 U3093 ( .A(n5062), .ZN(n1889) );
  AOI222_X1 U3094 ( .A1(n1892), .A2(n1290), .B1(n1291), .B2(n1893), .C1(n1894), 
        .C2(n1294), .ZN(n1875) );
  AND4_X1 U3095 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(n5431)
         );
  NOR4_X1 U3096 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898)
         );
  NAND3_X1 U3097 ( .A1(n5733), .A2(n5728), .A3(n5740), .ZN(n1902) );
  OAI211_X1 U3098 ( .C1(n5745), .C2(n5381), .A(n5718), .B(n5723), .ZN(n1901)
         );
  OAI222_X1 U3099 ( .A1(n5743), .A2(n5253), .B1(n5744), .B2(n5221), .C1(n5746), 
        .C2(n5349), .ZN(n1900) );
  OAI221_X1 U3100 ( .B1(n5716), .B2(n5157), .C1(n5717), .C2(n5189), .A(n1903), 
        .ZN(n1899) );
  AOI22_X1 U3101 ( .A1(n1904), .A2(n1275), .B1(n1905), .B2(n1277), .ZN(n1903)
         );
  AOI211_X1 U3104 ( .C1(n1906), .C2(n1279), .A(n1907), .B(n1908), .ZN(n1897)
         );
  OAI22_X1 U3105 ( .A1(n5726), .A2(n4805), .B1(n5736), .B2(n4709), .ZN(n1908)
         );
  OAI222_X1 U3106 ( .A1(n5731), .A2(n4645), .B1(n5737), .B2(n4613), .C1(n5732), 
        .C2(n4677), .ZN(n1907) );
  AOI221_X1 U3108 ( .B1(n1282), .B2(n1909), .C1(n1284), .C2(n1910), .A(n1911), 
        .ZN(n1896) );
  OAI22_X1 U3109 ( .A1(n4453), .A2(n1287), .B1(n5285), .B2(n1288), .ZN(n1911)
         );
  INV_X1 U3113 ( .A(n6022), .ZN(n1912) );
  INV_X1 U3114 ( .A(n5061), .ZN(n1909) );
  AOI222_X1 U3116 ( .A1(n1913), .A2(n1290), .B1(n1291), .B2(n1914), .C1(n1915), 
        .C2(n1294), .ZN(n1895) );
  INV_X1 U3120 ( .A(\UUT/Mcontrol/d_sampled_finstr [4]), .ZN(n5424) );
  INV_X1 U3121 ( .A(n1075), .ZN(n5422) );
  NAND4_X1 U3122 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1075)
         );
  NOR4_X1 U3123 ( .A1(n1920), .A2(n1921), .A3(n1922), .A4(n1923), .ZN(n1919)
         );
  NAND3_X1 U3124 ( .A1(n5610), .A2(n5609), .A3(n5611), .ZN(n1923) );
  OAI211_X1 U3125 ( .C1(n5560), .C2(n5412), .A(n5607), .B(n5608), .ZN(n1922)
         );
  OAI222_X1 U3126 ( .A1(n5558), .A2(n5284), .B1(n5559), .B2(n5252), .C1(n5561), 
        .C2(n5380), .ZN(n1921) );
  OAI221_X1 U3127 ( .B1(n5531), .B2(n5188), .C1(n5532), .C2(n5220), .A(n1924), 
        .ZN(n1920) );
  AOI22_X1 U3128 ( .A1(n1274), .A2(n1925), .B1(n1276), .B2(n1926), .ZN(n1924)
         );
  INV_X1 U3129 ( .A(n4996), .ZN(n1276) );
  INV_X1 U3130 ( .A(n4964), .ZN(n1274) );
  AOI211_X1 U3131 ( .C1(n1278), .C2(n1927), .A(n1928), .B(n1929), .ZN(n1918)
         );
  OAI22_X1 U3132 ( .A1(n5541), .A2(n4836), .B1(n5551), .B2(n4740), .ZN(n1929)
         );
  OAI222_X1 U3133 ( .A1(n5546), .A2(n4676), .B1(n5552), .B2(n4644), .C1(n5547), 
        .C2(n4708), .ZN(n1928) );
  INV_X1 U3134 ( .A(n4868), .ZN(n1278) );
  AOI221_X1 U3135 ( .B1(n1930), .B2(n1285), .C1(n1931), .C2(n1932), .A(n1933), 
        .ZN(n1917) );
  OAI22_X1 U3136 ( .A1(n4484), .A2(n1934), .B1(n5092), .B2(n1935), .ZN(n1933)
         );
  INV_X1 U3137 ( .A(n5316), .ZN(n1932) );
  INV_X1 U3138 ( .A(n5348), .ZN(n1285) );
  AOI222_X1 U3139 ( .A1(n1289), .A2(n1936), .B1(n1937), .B2(n1292), .C1(n1293), 
        .C2(n1938), .ZN(n1916) );
  INV_X1 U3140 ( .A(n4516), .ZN(n1293) );
  INV_X1 U3141 ( .A(n4452), .ZN(n1292) );
  INV_X1 U3142 ( .A(n4548), .ZN(n1289) );
  AND4_X1 U3143 ( .A1(n1939), .A2(n1940), .A3(n1941), .A4(n1942), .ZN(n5421)
         );
  NOR4_X1 U3144 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(n1942)
         );
  NAND3_X1 U3145 ( .A1(n5603), .A2(n5602), .A3(n5604), .ZN(n1946) );
  OAI211_X1 U3146 ( .C1(n5560), .C2(n5396), .A(n5600), .B(n5601), .ZN(n1945)
         );
  OAI222_X1 U3147 ( .A1(n5558), .A2(n5268), .B1(n5559), .B2(n5236), .C1(n5561), 
        .C2(n5364), .ZN(n1944) );
  OAI221_X1 U3148 ( .B1(n5531), .B2(n5172), .C1(n5532), .C2(n5204), .A(n1947), 
        .ZN(n1943) );
  AOI22_X1 U3149 ( .A1(n1604), .A2(n1925), .B1(n1605), .B2(n1926), .ZN(n1947)
         );
  INV_X1 U3150 ( .A(n4980), .ZN(n1605) );
  INV_X1 U3151 ( .A(n4948), .ZN(n1604) );
  AOI211_X1 U3152 ( .C1(n1606), .C2(n1927), .A(n1948), .B(n1949), .ZN(n1941)
         );
  OAI22_X1 U3153 ( .A1(n5541), .A2(n4820), .B1(n5551), .B2(n4724), .ZN(n1949)
         );
  OAI222_X1 U3154 ( .A1(n5546), .A2(n4660), .B1(n5552), .B2(n4628), .C1(n5547), 
        .C2(n4692), .ZN(n1948) );
  INV_X1 U3155 ( .A(n4852), .ZN(n1606) );
  AOI221_X1 U3156 ( .B1(n1930), .B2(n1610), .C1(n1931), .C2(n1950), .A(n1951), 
        .ZN(n1940) );
  OAI22_X1 U3157 ( .A1(n4468), .A2(n1934), .B1(n5076), .B2(n6373), .ZN(n1951)
         );
  INV_X1 U3158 ( .A(n5300), .ZN(n1950) );
  INV_X1 U3159 ( .A(n5332), .ZN(n1610) );
  AOI222_X1 U3160 ( .A1(n1612), .A2(n1936), .B1(n1937), .B2(n1613), .C1(n1614), 
        .C2(n1938), .ZN(n1939) );
  INV_X1 U3161 ( .A(n4500), .ZN(n1614) );
  INV_X1 U3162 ( .A(n4436), .ZN(n1613) );
  INV_X1 U3163 ( .A(n4532), .ZN(n1612) );
  AND4_X1 U3164 ( .A1(n1952), .A2(n1953), .A3(n1954), .A4(n1955), .ZN(n5420)
         );
  NOR4_X1 U3165 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .ZN(n1955)
         );
  NAND3_X1 U3166 ( .A1(n5596), .A2(n5595), .A3(n5597), .ZN(n1959) );
  OAI211_X1 U3167 ( .C1(n5560), .C2(n5395), .A(n5593), .B(n5594), .ZN(n1958)
         );
  OAI222_X1 U3168 ( .A1(n5558), .A2(n5267), .B1(n5559), .B2(n5235), .C1(n5561), 
        .C2(n5363), .ZN(n1957) );
  OAI221_X1 U3169 ( .B1(n5531), .B2(n5171), .C1(n5532), .C2(n5203), .A(n1960), 
        .ZN(n1956) );
  AOI22_X1 U3170 ( .A1(n1624), .A2(n1925), .B1(n1625), .B2(n1926), .ZN(n1960)
         );
  INV_X1 U3171 ( .A(n4979), .ZN(n1625) );
  INV_X1 U3172 ( .A(n4947), .ZN(n1624) );
  AOI211_X1 U3173 ( .C1(n1626), .C2(n1927), .A(n1961), .B(n1962), .ZN(n1954)
         );
  OAI22_X1 U3174 ( .A1(n5541), .A2(n4819), .B1(n5551), .B2(n4723), .ZN(n1962)
         );
  OAI222_X1 U3175 ( .A1(n5546), .A2(n4659), .B1(n5552), .B2(n4627), .C1(n5547), 
        .C2(n4691), .ZN(n1961) );
  INV_X1 U3176 ( .A(n4851), .ZN(n1626) );
  AOI221_X1 U3177 ( .B1(n1930), .B2(n1630), .C1(n1931), .C2(n1963), .A(n1964), 
        .ZN(n1953) );
  OAI22_X1 U3178 ( .A1(n4467), .A2(n1934), .B1(n5075), .B2(n6373), .ZN(n1964)
         );
  INV_X1 U3179 ( .A(n5299), .ZN(n1963) );
  INV_X1 U3180 ( .A(n5331), .ZN(n1630) );
  AOI222_X1 U3181 ( .A1(n1632), .A2(n1936), .B1(n1937), .B2(n1633), .C1(n1634), 
        .C2(n1938), .ZN(n1952) );
  INV_X1 U3182 ( .A(n4499), .ZN(n1634) );
  INV_X1 U3183 ( .A(n4435), .ZN(n1633) );
  INV_X1 U3184 ( .A(n4531), .ZN(n1632) );
  AND4_X1 U3185 ( .A1(n1965), .A2(n1966), .A3(n1967), .A4(n1968), .ZN(n5419)
         );
  NOR4_X1 U3186 ( .A1(n1969), .A2(n1970), .A3(n1971), .A4(n1972), .ZN(n1968)
         );
  NAND3_X1 U3187 ( .A1(n5589), .A2(n5588), .A3(n5590), .ZN(n1972) );
  OAI211_X1 U3188 ( .C1(n5560), .C2(n5394), .A(n5586), .B(n5587), .ZN(n1971)
         );
  OAI222_X1 U3189 ( .A1(n5558), .A2(n5266), .B1(n5559), .B2(n5234), .C1(n5561), 
        .C2(n5362), .ZN(n1970) );
  OAI221_X1 U3190 ( .B1(n5531), .B2(n5170), .C1(n5532), .C2(n5202), .A(n1973), 
        .ZN(n1969) );
  AOI22_X1 U3191 ( .A1(n1644), .A2(n1925), .B1(n1645), .B2(n1926), .ZN(n1973)
         );
  INV_X1 U3192 ( .A(n4978), .ZN(n1645) );
  INV_X1 U3193 ( .A(n4946), .ZN(n1644) );
  AOI211_X1 U3194 ( .C1(n1646), .C2(n1927), .A(n1974), .B(n1975), .ZN(n1967)
         );
  OAI22_X1 U3195 ( .A1(n5541), .A2(n4818), .B1(n5551), .B2(n4722), .ZN(n1975)
         );
  OAI222_X1 U3196 ( .A1(n5546), .A2(n4658), .B1(n5552), .B2(n4626), .C1(n5547), 
        .C2(n4690), .ZN(n1974) );
  INV_X1 U3197 ( .A(n4850), .ZN(n1646) );
  AOI221_X1 U3198 ( .B1(n1930), .B2(n1650), .C1(n1931), .C2(n1976), .A(n1977), 
        .ZN(n1966) );
  OAI22_X1 U3199 ( .A1(n4466), .A2(n1934), .B1(n5074), .B2(n6373), .ZN(n1977)
         );
  INV_X1 U3200 ( .A(n5298), .ZN(n1976) );
  INV_X1 U3201 ( .A(n5330), .ZN(n1650) );
  AOI222_X1 U3202 ( .A1(n1652), .A2(n1936), .B1(n1937), .B2(n1653), .C1(n1654), 
        .C2(n1938), .ZN(n1965) );
  INV_X1 U3203 ( .A(n4498), .ZN(n1654) );
  INV_X1 U3204 ( .A(n4434), .ZN(n1653) );
  INV_X1 U3205 ( .A(n4530), .ZN(n1652) );
  AND4_X1 U3206 ( .A1(n1978), .A2(n1979), .A3(n1980), .A4(n1981), .ZN(n5418)
         );
  NOR4_X1 U3207 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(n1981)
         );
  NAND3_X1 U3208 ( .A1(n5582), .A2(n5581), .A3(n5583), .ZN(n1985) );
  OAI211_X1 U3209 ( .C1(n5560), .C2(n5393), .A(n5579), .B(n5580), .ZN(n1984)
         );
  OAI222_X1 U3210 ( .A1(n5558), .A2(n5265), .B1(n5559), .B2(n5233), .C1(n5561), 
        .C2(n5361), .ZN(n1983) );
  OAI221_X1 U3211 ( .B1(n5531), .B2(n5169), .C1(n5532), .C2(n5201), .A(n1986), 
        .ZN(n1982) );
  AOI22_X1 U3212 ( .A1(n1664), .A2(n1925), .B1(n1665), .B2(n1926), .ZN(n1986)
         );
  INV_X1 U3213 ( .A(n4977), .ZN(n1665) );
  INV_X1 U3214 ( .A(n4945), .ZN(n1664) );
  AOI211_X1 U3215 ( .C1(n1666), .C2(n1927), .A(n1987), .B(n1988), .ZN(n1980)
         );
  OAI22_X1 U3216 ( .A1(n5541), .A2(n4817), .B1(n5551), .B2(n4721), .ZN(n1988)
         );
  OAI222_X1 U3217 ( .A1(n5546), .A2(n4657), .B1(n5552), .B2(n4625), .C1(n5547), 
        .C2(n4689), .ZN(n1987) );
  INV_X1 U3218 ( .A(n4849), .ZN(n1666) );
  AOI221_X1 U3219 ( .B1(n1930), .B2(n1670), .C1(n1931), .C2(n1989), .A(n1990), 
        .ZN(n1979) );
  OAI22_X1 U3220 ( .A1(n4465), .A2(n1934), .B1(n5073), .B2(n6373), .ZN(n1990)
         );
  INV_X1 U3221 ( .A(n5297), .ZN(n1989) );
  INV_X1 U3222 ( .A(n5329), .ZN(n1670) );
  AOI222_X1 U3223 ( .A1(n1672), .A2(n1936), .B1(n1937), .B2(n1673), .C1(n1674), 
        .C2(n1938), .ZN(n1978) );
  INV_X1 U3224 ( .A(n4497), .ZN(n1674) );
  INV_X1 U3225 ( .A(n4433), .ZN(n1673) );
  INV_X1 U3226 ( .A(n4529), .ZN(n1672) );
  AND4_X1 U3227 ( .A1(n1991), .A2(n1992), .A3(n1993), .A4(n1994), .ZN(n5417)
         );
  NOR4_X1 U3228 ( .A1(n1995), .A2(n1996), .A3(n1997), .A4(n1998), .ZN(n1994)
         );
  NAND3_X1 U3229 ( .A1(n5575), .A2(n5574), .A3(n5576), .ZN(n1998) );
  OAI211_X1 U3230 ( .C1(n5560), .C2(n5392), .A(n5572), .B(n5573), .ZN(n1997)
         );
  OAI222_X1 U3231 ( .A1(n5558), .A2(n5264), .B1(n5559), .B2(n5232), .C1(n5561), 
        .C2(n5360), .ZN(n1996) );
  OAI221_X1 U3232 ( .B1(n5531), .B2(n5168), .C1(n5532), .C2(n5200), .A(n1999), 
        .ZN(n1995) );
  AOI22_X1 U3233 ( .A1(n1684), .A2(n1925), .B1(n1685), .B2(n1926), .ZN(n1999)
         );
  INV_X1 U3234 ( .A(n4976), .ZN(n1685) );
  INV_X1 U3235 ( .A(n4944), .ZN(n1684) );
  AOI211_X1 U3236 ( .C1(n1686), .C2(n1927), .A(n2000), .B(n2001), .ZN(n1993)
         );
  OAI22_X1 U3237 ( .A1(n5541), .A2(n4816), .B1(n5551), .B2(n4720), .ZN(n2001)
         );
  OAI222_X1 U3238 ( .A1(n5546), .A2(n4656), .B1(n5552), .B2(n4624), .C1(n5547), 
        .C2(n4688), .ZN(n2000) );
  INV_X1 U3239 ( .A(n4848), .ZN(n1686) );
  AOI221_X1 U3240 ( .B1(n1930), .B2(n1690), .C1(n1931), .C2(n2002), .A(n2003), 
        .ZN(n1992) );
  OAI22_X1 U3241 ( .A1(n4464), .A2(n1934), .B1(n5072), .B2(n6373), .ZN(n2003)
         );
  INV_X1 U3242 ( .A(n5296), .ZN(n2002) );
  INV_X1 U3243 ( .A(n5328), .ZN(n1690) );
  AOI222_X1 U3244 ( .A1(n1692), .A2(n1936), .B1(n1937), .B2(n1693), .C1(n1694), 
        .C2(n1938), .ZN(n1991) );
  INV_X1 U3245 ( .A(n4496), .ZN(n1694) );
  INV_X1 U3246 ( .A(n4432), .ZN(n1693) );
  INV_X1 U3247 ( .A(n4528), .ZN(n1692) );
  AND4_X1 U3248 ( .A1(n2004), .A2(n2005), .A3(n2006), .A4(n2007), .ZN(n5416)
         );
  NOR4_X1 U3249 ( .A1(n2008), .A2(n2009), .A3(n2010), .A4(n2011), .ZN(n2007)
         );
  NAND3_X1 U3250 ( .A1(n5568), .A2(n5567), .A3(n5569), .ZN(n2011) );
  OAI211_X1 U3251 ( .C1(n5560), .C2(n5391), .A(n5565), .B(n5566), .ZN(n2010)
         );
  OAI222_X1 U3252 ( .A1(n5558), .A2(n5263), .B1(n5559), .B2(n5231), .C1(n5561), 
        .C2(n5359), .ZN(n2009) );
  OAI221_X1 U3253 ( .B1(n5531), .B2(n5167), .C1(n5532), .C2(n5199), .A(n2012), 
        .ZN(n2008) );
  AOI22_X1 U3254 ( .A1(n1704), .A2(n1925), .B1(n1705), .B2(n1926), .ZN(n2012)
         );
  INV_X1 U3255 ( .A(n4975), .ZN(n1705) );
  INV_X1 U3256 ( .A(n4943), .ZN(n1704) );
  AOI211_X1 U3257 ( .C1(n1706), .C2(n1927), .A(n2013), .B(n2014), .ZN(n2006)
         );
  OAI22_X1 U3258 ( .A1(n5541), .A2(n4815), .B1(n5551), .B2(n4719), .ZN(n2014)
         );
  OAI222_X1 U3259 ( .A1(n5546), .A2(n4655), .B1(n5552), .B2(n4623), .C1(n5547), 
        .C2(n4687), .ZN(n2013) );
  INV_X1 U3260 ( .A(n4847), .ZN(n1706) );
  AOI221_X1 U3261 ( .B1(n1930), .B2(n1710), .C1(n1931), .C2(n2015), .A(n2016), 
        .ZN(n2005) );
  OAI22_X1 U3262 ( .A1(n4463), .A2(n1934), .B1(n5071), .B2(n6373), .ZN(n2016)
         );
  INV_X1 U3263 ( .A(n5295), .ZN(n2015) );
  INV_X1 U3264 ( .A(n5327), .ZN(n1710) );
  AOI222_X1 U3265 ( .A1(n1712), .A2(n1936), .B1(n1937), .B2(n1713), .C1(n1714), 
        .C2(n1938), .ZN(n2004) );
  INV_X1 U3266 ( .A(n4495), .ZN(n1714) );
  INV_X1 U3267 ( .A(n4431), .ZN(n1713) );
  INV_X1 U3268 ( .A(n4527), .ZN(n1712) );
  AND4_X1 U3269 ( .A1(n2017), .A2(n2018), .A3(n2019), .A4(n2020), .ZN(n5415)
         );
  NOR4_X1 U3270 ( .A1(n2021), .A2(n2022), .A3(n2023), .A4(n2024), .ZN(n2020)
         );
  NAND3_X1 U3271 ( .A1(n5548), .A2(n5543), .A3(n5555), .ZN(n2024) );
  OAI211_X1 U3272 ( .C1(n5560), .C2(n5389), .A(n5533), .B(n5538), .ZN(n2023)
         );
  OAI222_X1 U3273 ( .A1(n5558), .A2(n5261), .B1(n5559), .B2(n5229), .C1(n5561), 
        .C2(n5357), .ZN(n2022) );
  OAI221_X1 U3274 ( .B1(n5531), .B2(n5165), .C1(n5532), .C2(n5197), .A(n2025), 
        .ZN(n2021) );
  AOI22_X1 U3275 ( .A1(n1744), .A2(n1925), .B1(n1745), .B2(n1926), .ZN(n2025)
         );
  INV_X1 U3276 ( .A(n4973), .ZN(n1745) );
  INV_X1 U3277 ( .A(n4941), .ZN(n1744) );
  AOI211_X1 U3278 ( .C1(n1746), .C2(n1927), .A(n2026), .B(n2027), .ZN(n2019)
         );
  OAI22_X1 U3279 ( .A1(n5541), .A2(n4813), .B1(n5551), .B2(n4717), .ZN(n2027)
         );
  OAI222_X1 U3280 ( .A1(n5546), .A2(n4653), .B1(n5552), .B2(n4621), .C1(n5547), 
        .C2(n4685), .ZN(n2026) );
  INV_X1 U3281 ( .A(n4845), .ZN(n1746) );
  AOI221_X1 U3282 ( .B1(n1930), .B2(n1750), .C1(n1931), .C2(n2028), .A(n2029), 
        .ZN(n2018) );
  OAI22_X1 U3283 ( .A1(n4461), .A2(n1934), .B1(n5069), .B2(n6373), .ZN(n2029)
         );
  INV_X1 U3284 ( .A(n5293), .ZN(n2028) );
  INV_X1 U3285 ( .A(n5325), .ZN(n1750) );
  AOI222_X1 U3286 ( .A1(n1752), .A2(n1936), .B1(n1937), .B2(n1753), .C1(n1754), 
        .C2(n1938), .ZN(n2017) );
  INV_X1 U3287 ( .A(n4493), .ZN(n1754) );
  INV_X1 U3288 ( .A(n4429), .ZN(n1753) );
  INV_X1 U3289 ( .A(n4525), .ZN(n1752) );
  AND4_X1 U3290 ( .A1(n2030), .A2(n2031), .A3(n2032), .A4(n2033), .ZN(n5414)
         );
  NOR4_X1 U3291 ( .A1(n2034), .A2(n2035), .A3(n2036), .A4(n2037), .ZN(n2033)
         );
  NAND3_X1 U3292 ( .A1(n6315), .A2(n6311), .A3(n6320), .ZN(n2037) );
  OAI211_X1 U3293 ( .C1(n5560), .C2(n5388), .A(n6300), .B(n6307), .ZN(n2036)
         );
  OAI222_X1 U3294 ( .A1(n5558), .A2(n5260), .B1(n5559), .B2(n5228), .C1(n5561), 
        .C2(n5356), .ZN(n2035) );
  OAI221_X1 U3295 ( .B1(n5531), .B2(n5164), .C1(n5532), .C2(n5196), .A(n2038), 
        .ZN(n2034) );
  AOI22_X1 U3296 ( .A1(n1764), .A2(n1925), .B1(n1765), .B2(n1926), .ZN(n2038)
         );
  INV_X1 U3297 ( .A(n4972), .ZN(n1765) );
  INV_X1 U3298 ( .A(n4940), .ZN(n1764) );
  AOI211_X1 U3299 ( .C1(n1766), .C2(n1927), .A(n2039), .B(n2040), .ZN(n2032)
         );
  OAI22_X1 U3300 ( .A1(n5541), .A2(n4812), .B1(n5551), .B2(n4716), .ZN(n2040)
         );
  OAI222_X1 U3301 ( .A1(n5546), .A2(n4652), .B1(n5552), .B2(n4620), .C1(n5547), 
        .C2(n4684), .ZN(n2039) );
  INV_X1 U3302 ( .A(n4844), .ZN(n1766) );
  AOI221_X1 U3303 ( .B1(n1930), .B2(n1770), .C1(n1931), .C2(n2041), .A(n2042), 
        .ZN(n2031) );
  OAI22_X1 U3304 ( .A1(n4460), .A2(n1934), .B1(n5068), .B2(n6373), .ZN(n2042)
         );
  INV_X1 U3305 ( .A(n5292), .ZN(n2041) );
  INV_X1 U3306 ( .A(n5324), .ZN(n1770) );
  AOI222_X1 U3307 ( .A1(n1772), .A2(n1936), .B1(n1937), .B2(n1773), .C1(n1774), 
        .C2(n1938), .ZN(n2030) );
  INV_X1 U3308 ( .A(n4492), .ZN(n1774) );
  INV_X1 U3309 ( .A(n4428), .ZN(n1773) );
  INV_X1 U3310 ( .A(n4524), .ZN(n1772) );
  NAND2_X1 U3311 ( .A1(n977), .A2(n1059), .ZN(dmem_read) );
  INV_X1 U3312 ( .A(\UUT/Mcontrol/x_sampled_dmem_command[MR] ), .ZN(n1059) );
  NAND2_X1 U3313 ( .A1(n977), .A2(n1054), .ZN(dmem_ishalf) );
  INV_X1 U3314 ( .A(\UUT/Mcontrol/x_sampled_dmem_command[MH] ), .ZN(n1054) );
  NAND2_X1 U3315 ( .A1(n977), .A2(n1047), .ZN(dmem_isbyte) );
  INV_X1 U3316 ( .A(\UUT/Mcontrol/x_sampled_dmem_command[MB] ), .ZN(n1047) );
  INV_X1 U3317 ( .A(\UUT/x_we ), .ZN(n977) );
  NOR2_X1 U3318 ( .A1(\UUT/regfile/N267 ), .A2(n2043), .ZN(\UUT/regfile/N269 )
         );
  INV_X1 U3319 ( .A(n6007), .ZN(n2043) );
  NAND2_X1 U3320 ( .A1(n2044), .A2(n2045), .ZN(\UUT/daddr_out [0]) );
  AOI21_X1 U3321 ( .B1(\UUT/Mpath/the_alu/diff[0] ), .B2(n1210), .A(n2046), 
        .ZN(n2045) );
  NOR3_X1 U3322 ( .A1(n2047), .A2(n2048), .A3(n1211), .ZN(n2046) );
  AOI22_X1 U3323 ( .A1(n2049), .A2(\UUT/Mpath/the_alu/N93 ), .B1(
        \UUT/Mpath/the_alu/N91 ), .B2(n2050), .ZN(n2048) );
  AND2_X1 U3324 ( .A1(\UUT/Mpath/the_alu/N498 ), .A2(\UUT/Mpath/the_alu/N503 ), 
        .ZN(n2049) );
  AOI22_X1 U3325 ( .A1(\UUT/Mpath/the_alu/sum[0] ), .A2(n1211), .B1(n6351), 
        .B2(n6348), .ZN(n2044) );
  INV_X1 U3326 ( .A(n1025), .ZN(\UUT/d_mul_command [5]) );
  NAND2_X1 U3327 ( .A1(n2051), .A2(\UUT/Mcontrol/d_sampled_finstr [5]), .ZN(
        n1025) );
  INV_X1 U3328 ( .A(n1022), .ZN(\UUT/d_mul_command [4]) );
  NAND2_X1 U3329 ( .A1(n2051), .A2(\UUT/Mcontrol/d_sampled_finstr [4]), .ZN(
        n1022) );
  NAND2_X1 U3330 ( .A1(n2051), .A2(n5425), .ZN(\UUT/d_mul_command [3]) );
  NAND2_X1 U3331 ( .A1(n2051), .A2(n5426), .ZN(\UUT/d_mul_command [2]) );
  NAND2_X1 U3332 ( .A1(n2051), .A2(n5427), .ZN(\UUT/d_mul_command [1]) );
  NAND2_X1 U3333 ( .A1(n2051), .A2(n5428), .ZN(\UUT/d_mul_command [0]) );
  AND2_X1 U3334 ( .A1(n927), .A2(\UUT/Mcontrol/Operation_decoding32/N2043 ), 
        .ZN(n2051) );
  INV_X1 U3335 ( .A(\UUT/Mcontrol/st_logic/N42 ), .ZN(\UUT/byp_controlB[0] )
         );
  INV_X1 U3336 ( .A(n117), .ZN(\UUT/break_code[23] ) );
  AOI221_X1 U3337 ( .B1(n6093), .B2(n2052), .C1(\UUT/Mcontrol/d_instr [7]), 
        .C2(n2053), .A(n2054), .ZN(n117) );
  INV_X1 U3338 ( .A(n292), .ZN(\UUT/break_code[22] ) );
  AOI221_X1 U3339 ( .B1(n6101), .B2(n2052), .C1(n2053), .C2(
        \UUT/Mcontrol/d_instr [6]), .A(n2054), .ZN(n292) );
  INV_X1 U3340 ( .A(n327), .ZN(\UUT/break_code[21] ) );
  AOI221_X1 U3341 ( .B1(n6108), .B2(n2052), .C1(\UUT/Mcontrol/d_instr [5]), 
        .C2(n2053), .A(n2054), .ZN(n327) );
  INV_X1 U3342 ( .A(n348), .ZN(\UUT/break_code[20] ) );
  AOI221_X1 U3343 ( .B1(n6115), .B2(n2052), .C1(\UUT/Mcontrol/d_instr [4]), 
        .C2(n2053), .A(n2054), .ZN(n348) );
  OAI21_X1 U3344 ( .B1(n1169), .B2(n855), .A(n2055), .ZN(n2054) );
  INV_X1 U3345 ( .A(n448), .ZN(n2055) );
  NAND3_X1 U3346 ( .A1(\UUT/Mcontrol/d_sampled_finstr [15]), .A2(n1216), .A3(
        n857), .ZN(n855) );
  NOR2_X1 U3347 ( .A1(n1168), .A2(n1169), .ZN(n2052) );
  INV_X1 U3348 ( .A(n1167), .ZN(n1168) );
  NOR2_X1 U3349 ( .A1(n1216), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .ZN(n1167) );
  NAND4_X1 U3350 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1987 ), .A2(n1061), 
        .A3(n6042), .A4(\UUT/Mcontrol/Operation_decoding32/N1994 ), .ZN(n1216)
         );
  INV_X1 U3351 ( .A(n1064), .ZN(n6042) );
  NOR3_X1 U3352 ( .A1(\UUT/Mcontrol/d_instr [27]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2010 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .ZN(n1064) );
  OAI21_X1 U3353 ( .B1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .B2(n2056), 
        .A(n2057), .ZN(n1061) );
  NAND3_X1 U3354 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2005 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N2017 ), .ZN(n2057) );
  INV_X1 U3355 ( .A(\UUT/Mcontrol/Operation_decoding32/N1999 ), .ZN(n2056) );
  NAND2_X1 U3356 ( .A1(n2058), .A2(n2059), .ZN(\UUT/break_code[1] ) );
  NAND3_X1 U3357 ( .A1(n6086), .A2(n935), .A3(\UUT/Mcontrol/d_instr [7]), .ZN(
        n2059) );
  NAND2_X1 U3358 ( .A1(\UUT/Mcontrol/d_instr [1]), .A2(n2060), .ZN(n2058) );
  INV_X1 U3359 ( .A(n2061), .ZN(n2060) );
  OAI221_X1 U3360 ( .B1(n2062), .B2(n2063), .C1(n5425), .C2(n2064), .A(n2065), 
        .ZN(\UUT/break_code[19] ) );
  INV_X1 U3361 ( .A(\UUT/Mcontrol/d_sampled_finstr [3]), .ZN(n5425) );
  INV_X1 U3362 ( .A(n6126), .ZN(n2063) );
  OAI221_X1 U3363 ( .B1(n2062), .B2(n2066), .C1(n5426), .C2(n2064), .A(n2065), 
        .ZN(\UUT/break_code[18] ) );
  INV_X1 U3364 ( .A(\UUT/Mcontrol/d_sampled_finstr [2]), .ZN(n5426) );
  INV_X1 U3365 ( .A(n6135), .ZN(n2066) );
  OAI221_X1 U3366 ( .B1(n2062), .B2(n2067), .C1(n5427), .C2(n2064), .A(n2065), 
        .ZN(\UUT/break_code[17] ) );
  INV_X1 U3367 ( .A(\UUT/Mcontrol/d_sampled_finstr [1]), .ZN(n5427) );
  INV_X1 U3368 ( .A(n6153), .ZN(n2067) );
  OAI221_X1 U3369 ( .B1(n2062), .B2(n2068), .C1(n5428), .C2(n2064), .A(n2065), 
        .ZN(\UUT/break_code[16] ) );
  AOI21_X1 U3370 ( .B1(n6050), .B2(n6127), .A(n448), .ZN(n2065) );
  NOR3_X1 U3371 ( .A1(n933), .A2(n5831), .A3(n929), .ZN(n448) );
  INV_X1 U3372 ( .A(n2053), .ZN(n2064) );
  NOR2_X1 U3373 ( .A1(n857), .A2(n1169), .ZN(n2053) );
  INV_X1 U3374 ( .A(\UUT/Mcontrol/Operation_decoding32/N2025 ), .ZN(n857) );
  INV_X1 U3375 ( .A(\UUT/Mcontrol/d_sampled_finstr [0]), .ZN(n5428) );
  INV_X1 U3376 ( .A(n6162), .ZN(n2068) );
  NAND2_X1 U3377 ( .A1(n6050), .A2(n445), .ZN(n2062) );
  NOR2_X1 U3378 ( .A1(n1169), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .ZN(n6050) );
  NAND2_X1 U3379 ( .A1(n927), .A2(n931), .ZN(n1169) );
  INV_X1 U3381 ( .A(\UUT/Mcontrol/Operation_decoding32/N2030 ), .ZN(n943) );
  NOR2_X1 U3382 ( .A1(n933), .A2(n6170), .ZN(n927) );
  INV_X1 U3383 ( .A(n466), .ZN(\UUT/break_code[15] ) );
  NAND2_X1 U3384 ( .A1(n2069), .A2(n6030), .ZN(n466) );
  OAI22_X1 U3385 ( .A1(n6173), .A2(n2070), .B1(n5831), .B2(n2071), .ZN(n2069)
         );
  INV_X1 U3386 ( .A(n6170), .ZN(n2071) );
  INV_X1 U3387 ( .A(\UUT/Mcontrol/d_sampled_finstr [15]), .ZN(n5831) );
  OAI21_X1 U3388 ( .B1(n6032), .B2(n2072), .A(n2073), .ZN(\UUT/break_code[14] ) );
  NAND2_X1 U3389 ( .A1(n6181), .A2(n2074), .ZN(n2073) );
  INV_X1 U3390 ( .A(\UUT/Mcontrol/d_sampled_finstr [14]), .ZN(n6032) );
  OAI21_X1 U3391 ( .B1(n6033), .B2(n2072), .A(n2075), .ZN(\UUT/break_code[13] ) );
  NAND2_X1 U3392 ( .A1(n6188), .A2(n2074), .ZN(n2075) );
  INV_X1 U3393 ( .A(\UUT/Mcontrol/d_sampled_finstr [13]), .ZN(n6033) );
  OAI21_X1 U3394 ( .B1(n2061), .B2(\UUT/Mcontrol/Operation_decoding32/N1901 ), 
        .A(n2076), .ZN(\UUT/break_code[0] ) );
  NOR2_X1 U3397 ( .A1(n2077), .A2(n933), .ZN(n935) );
  AOI222_X1 U3399 ( .A1(n6092), .A2(n5564), .B1(n878), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[23] ), .C2(n5612), .ZN(n5480) );
  NAND2_X1 U3400 ( .A1(n2079), .A2(n2080), .ZN(n878) );
  AOI222_X1 U3401 ( .A1(\UUT/Mpath/the_shift/sh_ror [23]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [23]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [23]), .C2(n6199), .ZN(n2080) );
  AOI22_X1 U3402 ( .A1(\UUT/Mpath/the_shift/sh_sll [23]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [23]), .B2(n6198), .ZN(n2079) );
  NAND3_X1 U3403 ( .A1(n2081), .A2(n2082), .A3(n2083), .ZN(n6092) );
  AOI222_X1 U3404 ( .A1(n1208), .A2(n2084), .B1(\UUT/Mpath/the_alu/diff[23] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[23] ), .C2(n1211), .ZN(n2083)
         );
  INV_X1 U3405 ( .A(\UUT/Mpath/the_alu/N37 ), .ZN(n2084) );
  AOI22_X1 U3406 ( .A1(\UUT/Mpath/the_alu/N134 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N102 ), .B2(n1213), .ZN(n2082) );
  AOI22_X1 U3407 ( .A1(\UUT/Mpath/the_alu/N166 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N198 ), .B2(n1215), .ZN(n2081) );
  INV_X1 U3408 ( .A(n811), .ZN(n2078) );
  NAND4_X1 U3409 ( .A1(n2085), .A2(n2086), .A3(n2087), .A4(n2088), .ZN(n811)
         );
  NOR4_X1 U3410 ( .A1(n2089), .A2(n2090), .A3(n2091), .A4(n2092), .ZN(n2088)
         );
  NAND3_X1 U3411 ( .A1(n6090), .A2(n6089), .A3(n6091), .ZN(n2092) );
  OAI211_X1 U3412 ( .C1(n5560), .C2(n5397), .A(n6087), .B(n6088), .ZN(n2091)
         );
  OAI222_X1 U3413 ( .A1(n5558), .A2(n5269), .B1(n5559), .B2(n5237), .C1(n5561), 
        .C2(n5365), .ZN(n2090) );
  OAI221_X1 U3414 ( .B1(n5531), .B2(n5173), .C1(n5532), .C2(n5205), .A(n2093), 
        .ZN(n2089) );
  AOI22_X1 U3415 ( .A1(n1584), .A2(n1925), .B1(n1585), .B2(n1926), .ZN(n2093)
         );
  INV_X1 U3416 ( .A(n4981), .ZN(n1585) );
  INV_X1 U3417 ( .A(n4949), .ZN(n1584) );
  AOI211_X1 U3418 ( .C1(n1586), .C2(n1927), .A(n2094), .B(n2095), .ZN(n2087)
         );
  OAI22_X1 U3419 ( .A1(n5541), .A2(n4821), .B1(n5551), .B2(n4725), .ZN(n2095)
         );
  OAI222_X1 U3420 ( .A1(n5546), .A2(n4661), .B1(n5552), .B2(n4629), .C1(n5547), 
        .C2(n4693), .ZN(n2094) );
  INV_X1 U3421 ( .A(n4853), .ZN(n1586) );
  AOI221_X1 U3422 ( .B1(n1930), .B2(n1590), .C1(n1931), .C2(n2096), .A(n2097), 
        .ZN(n2086) );
  OAI22_X1 U3423 ( .A1(n4469), .A2(n1934), .B1(n5077), .B2(n6373), .ZN(n2097)
         );
  INV_X1 U3424 ( .A(n5301), .ZN(n2096) );
  INV_X1 U3425 ( .A(n5333), .ZN(n1590) );
  AOI222_X1 U3426 ( .A1(n1592), .A2(n1936), .B1(n1937), .B2(n1593), .C1(n1594), 
        .C2(n1938), .ZN(n2085) );
  INV_X1 U3427 ( .A(n4501), .ZN(n1594) );
  INV_X1 U3428 ( .A(n4437), .ZN(n1593) );
  INV_X1 U3429 ( .A(n4533), .ZN(n1592) );
  AOI222_X1 U3431 ( .A1(n6100), .A2(n5564), .B1(n324), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[22] ), .C2(n5612), .ZN(n5483) );
  NAND2_X1 U3432 ( .A1(n2099), .A2(n2100), .ZN(n324) );
  AOI222_X1 U3433 ( .A1(\UUT/Mpath/the_shift/sh_ror [22]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [22]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [22]), .C2(n6199), .ZN(n2100) );
  AOI22_X1 U3434 ( .A1(\UUT/Mpath/the_shift/sh_sll [22]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [22]), .B2(n6198), .ZN(n2099) );
  NAND3_X1 U3435 ( .A1(n2101), .A2(n2102), .A3(n2103), .ZN(n6100) );
  AOI222_X1 U3436 ( .A1(n1208), .A2(n2104), .B1(\UUT/Mpath/the_alu/diff[22] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[22] ), .C2(n1211), .ZN(n2103)
         );
  INV_X1 U3437 ( .A(\UUT/Mpath/the_alu/N39 ), .ZN(n2104) );
  AOI22_X1 U3438 ( .A1(\UUT/Mpath/the_alu/N135 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N103 ), .B2(n1213), .ZN(n2102) );
  AOI22_X1 U3439 ( .A1(\UUT/Mpath/the_alu/N167 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N199 ), .B2(n1215), .ZN(n2101) );
  INV_X1 U3440 ( .A(n313), .ZN(n2098) );
  NAND4_X1 U3441 ( .A1(n2105), .A2(n2106), .A3(n2107), .A4(n2108), .ZN(n313)
         );
  NOR4_X1 U3442 ( .A1(n2109), .A2(n2110), .A3(n2111), .A4(n2112), .ZN(n2108)
         );
  NAND3_X1 U3443 ( .A1(n6098), .A2(n6097), .A3(n6099), .ZN(n2112) );
  OAI211_X1 U3444 ( .C1(n5560), .C2(n5398), .A(n6095), .B(n6096), .ZN(n2111)
         );
  OAI222_X1 U3445 ( .A1(n5558), .A2(n5270), .B1(n5559), .B2(n5238), .C1(n5561), 
        .C2(n5366), .ZN(n2110) );
  OAI221_X1 U3446 ( .B1(n5531), .B2(n5174), .C1(n5532), .C2(n5206), .A(n2113), 
        .ZN(n2109) );
  AOI22_X1 U3447 ( .A1(n1564), .A2(n1925), .B1(n1565), .B2(n1926), .ZN(n2113)
         );
  INV_X1 U3448 ( .A(n4982), .ZN(n1565) );
  INV_X1 U3449 ( .A(n4950), .ZN(n1564) );
  AOI211_X1 U3450 ( .C1(n1566), .C2(n1927), .A(n2114), .B(n2115), .ZN(n2107)
         );
  OAI22_X1 U3451 ( .A1(n5541), .A2(n4822), .B1(n5551), .B2(n4726), .ZN(n2115)
         );
  OAI222_X1 U3452 ( .A1(n5546), .A2(n4662), .B1(n5552), .B2(n4630), .C1(n5547), 
        .C2(n4694), .ZN(n2114) );
  INV_X1 U3453 ( .A(n4854), .ZN(n1566) );
  AOI221_X1 U3454 ( .B1(n1930), .B2(n1570), .C1(n1931), .C2(n2116), .A(n2117), 
        .ZN(n2106) );
  OAI22_X1 U3455 ( .A1(n4470), .A2(n1934), .B1(n5078), .B2(n6373), .ZN(n2117)
         );
  INV_X1 U3456 ( .A(n5302), .ZN(n2116) );
  INV_X1 U3457 ( .A(n5334), .ZN(n1570) );
  AOI222_X1 U3458 ( .A1(n1572), .A2(n1936), .B1(n1937), .B2(n1573), .C1(n1574), 
        .C2(n1938), .ZN(n2105) );
  INV_X1 U3459 ( .A(n4502), .ZN(n1574) );
  INV_X1 U3460 ( .A(n4438), .ZN(n1573) );
  INV_X1 U3461 ( .A(n4534), .ZN(n1572) );
  OAI222_X1 U3462 ( .A1(n5488), .A2(n5530), .B1(n6364), .B2(n2118), .C1(n5528), 
        .C2(n5486), .ZN(\UUT/branch_rega [21]) );
  NAND2_X1 U3464 ( .A1(n2119), .A2(n2120), .ZN(n346) );
  AOI222_X1 U3465 ( .A1(\UUT/Mpath/the_shift/sh_ror [21]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [21]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [21]), .C2(n6199), .ZN(n2120) );
  AOI22_X1 U3466 ( .A1(\UUT/Mpath/the_shift/sh_sll [21]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [21]), .B2(n6198), .ZN(n2119) );
  NAND3_X1 U3467 ( .A1(n2121), .A2(n2122), .A3(n2123), .ZN(n6107) );
  AOI222_X1 U3468 ( .A1(n1208), .A2(n2124), .B1(\UUT/Mpath/the_alu/diff[21] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[21] ), .C2(n1211), .ZN(n2123)
         );
  INV_X1 U3469 ( .A(\UUT/Mpath/the_alu/N41 ), .ZN(n2124) );
  AOI22_X1 U3470 ( .A1(\UUT/Mpath/the_alu/N136 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N104 ), .B2(n1213), .ZN(n2122) );
  AOI22_X1 U3471 ( .A1(\UUT/Mpath/the_alu/N168 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N200 ), .B2(n1215), .ZN(n2121) );
  INV_X1 U3472 ( .A(n340), .ZN(n2118) );
  NAND4_X1 U3473 ( .A1(n2125), .A2(n2126), .A3(n2127), .A4(n2128), .ZN(n340)
         );
  NOR4_X1 U3474 ( .A1(n2129), .A2(n2130), .A3(n2131), .A4(n2132), .ZN(n2128)
         );
  NAND3_X1 U3475 ( .A1(n6105), .A2(n6104), .A3(n6106), .ZN(n2132) );
  OAI211_X1 U3476 ( .C1(n5560), .C2(n5399), .A(n6102), .B(n6103), .ZN(n2131)
         );
  OAI222_X1 U3477 ( .A1(n5558), .A2(n5271), .B1(n5559), .B2(n5239), .C1(n5561), 
        .C2(n5367), .ZN(n2130) );
  OAI221_X1 U3478 ( .B1(n5531), .B2(n5175), .C1(n5532), .C2(n5207), .A(n2133), 
        .ZN(n2129) );
  AOI22_X1 U3479 ( .A1(n1544), .A2(n1925), .B1(n1545), .B2(n1926), .ZN(n2133)
         );
  INV_X1 U3480 ( .A(n4983), .ZN(n1545) );
  INV_X1 U3481 ( .A(n4951), .ZN(n1544) );
  AOI211_X1 U3482 ( .C1(n1546), .C2(n1927), .A(n2134), .B(n2135), .ZN(n2127)
         );
  OAI22_X1 U3483 ( .A1(n5541), .A2(n4823), .B1(n5551), .B2(n4727), .ZN(n2135)
         );
  OAI222_X1 U3484 ( .A1(n5546), .A2(n4663), .B1(n5552), .B2(n4631), .C1(n5547), 
        .C2(n4695), .ZN(n2134) );
  INV_X1 U3485 ( .A(n4855), .ZN(n1546) );
  AOI221_X1 U3486 ( .B1(n1930), .B2(n1550), .C1(n1931), .C2(n2136), .A(n2137), 
        .ZN(n2126) );
  OAI22_X1 U3487 ( .A1(n4471), .A2(n1934), .B1(n5079), .B2(n6373), .ZN(n2137)
         );
  INV_X1 U3488 ( .A(n5303), .ZN(n2136) );
  INV_X1 U3489 ( .A(n5335), .ZN(n1550) );
  AOI222_X1 U3490 ( .A1(n1552), .A2(n1936), .B1(n1937), .B2(n1553), .C1(n1554), 
        .C2(n1938), .ZN(n2125) );
  INV_X1 U3491 ( .A(n4503), .ZN(n1554) );
  INV_X1 U3492 ( .A(n4439), .ZN(n1553) );
  INV_X1 U3493 ( .A(n4535), .ZN(n1552) );
  OAI222_X1 U3494 ( .A1(n5491), .A2(n5530), .B1(n6364), .B2(n2138), .C1(n5528), 
        .C2(n5489), .ZN(\UUT/branch_rega [20]) );
  AOI222_X1 U3495 ( .A1(n6114), .A2(n5564), .B1(n367), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[20] ), .C2(n5612), .ZN(n5489) );
  NAND2_X1 U3496 ( .A1(n2139), .A2(n2140), .ZN(n367) );
  AOI222_X1 U3497 ( .A1(\UUT/Mpath/the_shift/sh_ror [20]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [20]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [20]), .C2(n6199), .ZN(n2140) );
  AOI22_X1 U3498 ( .A1(\UUT/Mpath/the_shift/sh_sll [20]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [20]), .B2(n6198), .ZN(n2139) );
  NAND3_X1 U3499 ( .A1(n2141), .A2(n2142), .A3(n2143), .ZN(n6114) );
  AOI222_X1 U3500 ( .A1(n1208), .A2(n2144), .B1(\UUT/Mpath/the_alu/diff[20] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[20] ), .C2(n1211), .ZN(n2143)
         );
  INV_X1 U3501 ( .A(\UUT/Mpath/the_alu/N43 ), .ZN(n2144) );
  AOI22_X1 U3502 ( .A1(\UUT/Mpath/the_alu/N137 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N105 ), .B2(n1213), .ZN(n2142) );
  AOI22_X1 U3503 ( .A1(\UUT/Mpath/the_alu/N169 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N201 ), .B2(n1215), .ZN(n2141) );
  INV_X1 U3504 ( .A(n361), .ZN(n2138) );
  NAND4_X1 U3505 ( .A1(n2145), .A2(n2146), .A3(n2147), .A4(n2148), .ZN(n361)
         );
  NOR4_X1 U3506 ( .A1(n2149), .A2(n2150), .A3(n2151), .A4(n2152), .ZN(n2148)
         );
  NAND3_X1 U3507 ( .A1(n6112), .A2(n6111), .A3(n6113), .ZN(n2152) );
  OAI211_X1 U3508 ( .C1(n5560), .C2(n5400), .A(n6109), .B(n6110), .ZN(n2151)
         );
  OAI222_X1 U3509 ( .A1(n5558), .A2(n5272), .B1(n5559), .B2(n5240), .C1(n5561), 
        .C2(n5368), .ZN(n2150) );
  OAI221_X1 U3510 ( .B1(n5531), .B2(n5176), .C1(n5532), .C2(n5208), .A(n2153), 
        .ZN(n2149) );
  AOI22_X1 U3511 ( .A1(n1524), .A2(n1925), .B1(n1525), .B2(n1926), .ZN(n2153)
         );
  INV_X1 U3512 ( .A(n4984), .ZN(n1525) );
  INV_X1 U3513 ( .A(n4952), .ZN(n1524) );
  AOI211_X1 U3514 ( .C1(n1526), .C2(n1927), .A(n2154), .B(n2155), .ZN(n2147)
         );
  OAI22_X1 U3515 ( .A1(n5541), .A2(n4824), .B1(n5551), .B2(n4728), .ZN(n2155)
         );
  OAI222_X1 U3516 ( .A1(n5546), .A2(n4664), .B1(n5552), .B2(n4632), .C1(n5547), 
        .C2(n4696), .ZN(n2154) );
  INV_X1 U3517 ( .A(n4856), .ZN(n1526) );
  AOI221_X1 U3518 ( .B1(n1930), .B2(n1530), .C1(n1931), .C2(n2156), .A(n2157), 
        .ZN(n2146) );
  OAI22_X1 U3519 ( .A1(n4472), .A2(n1934), .B1(n5080), .B2(n6373), .ZN(n2157)
         );
  INV_X1 U3520 ( .A(n5304), .ZN(n2156) );
  INV_X1 U3521 ( .A(n5336), .ZN(n1530) );
  AOI222_X1 U3522 ( .A1(n1532), .A2(n1936), .B1(n1937), .B2(n1533), .C1(n1534), 
        .C2(n1938), .ZN(n2145) );
  INV_X1 U3523 ( .A(n4504), .ZN(n1534) );
  INV_X1 U3524 ( .A(n4440), .ZN(n1533) );
  INV_X1 U3525 ( .A(n4536), .ZN(n1532) );
  OAI222_X1 U3526 ( .A1(n5494), .A2(n5530), .B1(n5529), .B2(n2158), .C1(n5528), 
        .C2(n5492), .ZN(\UUT/branch_rega [1]) );
  AOI222_X1 U3527 ( .A1(\UUT/daddr_out [1]), .A2(n5564), .B1(n822), .B2(
        \UUT/Mpath/N119 ), .C1(\UUT/Mpath/out_jar[1] ), .C2(n5612), .ZN(n5492)
         );
  NAND2_X1 U3528 ( .A1(n2159), .A2(n2160), .ZN(n822) );
  AOI222_X1 U3529 ( .A1(\UUT/Mpath/the_shift/sh_ror [1]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [1]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [1]), .C2(n6199), .ZN(n2160) );
  AOI22_X1 U3530 ( .A1(\UUT/Mpath/the_shift/sh_sll [1]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [1]), .B2(n6198), .ZN(n2159) );
  OAI211_X1 U3531 ( .C1(\UUT/Mpath/the_alu/N81 ), .C2(n2161), .A(n2162), .B(
        n2163), .ZN(\UUT/daddr_out [1]) );
  AOI22_X1 U3532 ( .A1(\UUT/Mpath/the_alu/diff[1] ), .A2(n1210), .B1(
        \UUT/Mpath/the_alu/sum[1] ), .B2(n1211), .ZN(n2163) );
  AOI22_X1 U3533 ( .A1(n2164), .A2(\UUT/Mpath/the_alu/N82 ), .B1(n2165), .B2(
        n2166), .ZN(n2162) );
  INV_X1 U3534 ( .A(n2167), .ZN(n2165) );
  AOI21_X1 U3535 ( .B1(n6365), .B2(\UUT/Mpath/the_alu/N81 ), .A(n1212), .ZN(
        n2167) );
  AND2_X1 U3536 ( .A1(n1215), .A2(\UUT/Mpath/the_alu/N81 ), .ZN(n2164) );
  NOR3_X1 U3537 ( .A1(n2168), .A2(n1208), .A3(n1212), .ZN(n2161) );
  INV_X1 U3538 ( .A(n2169), .ZN(n2168) );
  AOI22_X1 U3539 ( .A1(n6365), .A2(\UUT/Mpath/the_alu/N82 ), .B1(n2166), .B2(
        n1213), .ZN(n2169) );
  INV_X1 U3540 ( .A(\UUT/Mpath/the_alu/N82 ), .ZN(n2166) );
  INV_X1 U3541 ( .A(n799), .ZN(n2158) );
  NAND4_X1 U3542 ( .A1(n2170), .A2(n2171), .A3(n2172), .A4(n2173), .ZN(n799)
         );
  NOR4_X1 U3543 ( .A1(n2174), .A2(n2175), .A3(n2176), .A4(n2177), .ZN(n2173)
         );
  NAND3_X1 U3544 ( .A1(n6083), .A2(n6082), .A3(n6084), .ZN(n2177) );
  OAI211_X1 U3545 ( .C1(n5560), .C2(n5401), .A(n6080), .B(n6081), .ZN(n2176)
         );
  OAI222_X1 U3546 ( .A1(n5558), .A2(n5273), .B1(n5559), .B2(n5241), .C1(n5561), 
        .C2(n5369), .ZN(n2175) );
  OAI221_X1 U3547 ( .B1(n5531), .B2(n5177), .C1(n5532), .C2(n5209), .A(n2178), 
        .ZN(n2174) );
  AOI22_X1 U3548 ( .A1(n1504), .A2(n1925), .B1(n1505), .B2(n1926), .ZN(n2178)
         );
  INV_X1 U3549 ( .A(n4985), .ZN(n1505) );
  INV_X1 U3550 ( .A(n4953), .ZN(n1504) );
  AOI211_X1 U3551 ( .C1(n1506), .C2(n1927), .A(n2179), .B(n2180), .ZN(n2172)
         );
  OAI22_X1 U3552 ( .A1(n5541), .A2(n4825), .B1(n5551), .B2(n4729), .ZN(n2180)
         );
  OAI222_X1 U3553 ( .A1(n5546), .A2(n4665), .B1(n5552), .B2(n4633), .C1(n5547), 
        .C2(n4697), .ZN(n2179) );
  INV_X1 U3554 ( .A(n4857), .ZN(n1506) );
  AOI221_X1 U3555 ( .B1(n1930), .B2(n1510), .C1(n1931), .C2(n2181), .A(n2182), 
        .ZN(n2171) );
  OAI22_X1 U3556 ( .A1(n4473), .A2(n1934), .B1(n5081), .B2(n1935), .ZN(n2182)
         );
  INV_X1 U3557 ( .A(n5305), .ZN(n2181) );
  INV_X1 U3558 ( .A(n5337), .ZN(n1510) );
  AOI222_X1 U3559 ( .A1(n1512), .A2(n1936), .B1(n1937), .B2(n1513), .C1(n1514), 
        .C2(n1938), .ZN(n2170) );
  INV_X1 U3560 ( .A(n4505), .ZN(n1514) );
  INV_X1 U3561 ( .A(n4441), .ZN(n1513) );
  INV_X1 U3562 ( .A(n4537), .ZN(n1512) );
  OAI222_X1 U3563 ( .A1(n5497), .A2(n5530), .B1(n5529), .B2(n2183), .C1(n5528), 
        .C2(n5495), .ZN(\UUT/branch_rega [19]) );
  AOI222_X1 U3564 ( .A1(n6124), .A2(n5564), .B1(n393), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[19] ), .C2(n5612), .ZN(n5495) );
  NAND2_X1 U3565 ( .A1(n2184), .A2(n2185), .ZN(n393) );
  AOI222_X1 U3566 ( .A1(\UUT/Mpath/the_shift/sh_ror [19]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [19]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [19]), .C2(n6199), .ZN(n2185) );
  AOI22_X1 U3567 ( .A1(\UUT/Mpath/the_shift/sh_sll [19]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [19]), .B2(n6198), .ZN(n2184) );
  NAND3_X1 U3568 ( .A1(n2186), .A2(n2187), .A3(n2188), .ZN(n6124) );
  AOI222_X1 U3569 ( .A1(n1208), .A2(n2189), .B1(\UUT/Mpath/the_alu/diff[19] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[19] ), .C2(n1211), .ZN(n2188)
         );
  INV_X1 U3570 ( .A(\UUT/Mpath/the_alu/N45 ), .ZN(n2189) );
  AOI22_X1 U3571 ( .A1(\UUT/Mpath/the_alu/N138 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N106 ), .B2(n1213), .ZN(n2187) );
  AOI22_X1 U3572 ( .A1(\UUT/Mpath/the_alu/N170 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N202 ), .B2(n1215), .ZN(n2186) );
  INV_X1 U3573 ( .A(n387), .ZN(n2183) );
  NAND4_X1 U3574 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n387)
         );
  NOR4_X1 U3575 ( .A1(n2194), .A2(n2195), .A3(n2196), .A4(n2197), .ZN(n2193)
         );
  NAND3_X1 U3576 ( .A1(n6122), .A2(n6121), .A3(n6123), .ZN(n2197) );
  OAI211_X1 U3577 ( .C1(n5560), .C2(n5402), .A(n6119), .B(n6120), .ZN(n2196)
         );
  OAI222_X1 U3578 ( .A1(n5558), .A2(n5274), .B1(n5559), .B2(n5242), .C1(n5561), 
        .C2(n5370), .ZN(n2195) );
  OAI221_X1 U3579 ( .B1(n5531), .B2(n5178), .C1(n5532), .C2(n5210), .A(n2198), 
        .ZN(n2194) );
  AOI22_X1 U3580 ( .A1(n1484), .A2(n1925), .B1(n1485), .B2(n1926), .ZN(n2198)
         );
  INV_X1 U3581 ( .A(n4986), .ZN(n1485) );
  INV_X1 U3582 ( .A(n4954), .ZN(n1484) );
  AOI211_X1 U3583 ( .C1(n1486), .C2(n1927), .A(n2199), .B(n2200), .ZN(n2192)
         );
  OAI22_X1 U3584 ( .A1(n5541), .A2(n4826), .B1(n5551), .B2(n4730), .ZN(n2200)
         );
  OAI222_X1 U3585 ( .A1(n5546), .A2(n4666), .B1(n5552), .B2(n4634), .C1(n5547), 
        .C2(n4698), .ZN(n2199) );
  INV_X1 U3586 ( .A(n4858), .ZN(n1486) );
  AOI221_X1 U3587 ( .B1(n1930), .B2(n1490), .C1(n1931), .C2(n2201), .A(n2202), 
        .ZN(n2191) );
  OAI22_X1 U3588 ( .A1(n4474), .A2(n1934), .B1(n5082), .B2(n6373), .ZN(n2202)
         );
  INV_X1 U3589 ( .A(n5306), .ZN(n2201) );
  INV_X1 U3590 ( .A(n5338), .ZN(n1490) );
  AOI222_X1 U3591 ( .A1(n1492), .A2(n1936), .B1(n1937), .B2(n1493), .C1(n1494), 
        .C2(n1938), .ZN(n2190) );
  INV_X1 U3592 ( .A(n4506), .ZN(n1494) );
  INV_X1 U3593 ( .A(n4442), .ZN(n1493) );
  INV_X1 U3594 ( .A(n4538), .ZN(n1492) );
  NAND2_X1 U3597 ( .A1(n2204), .A2(n2205), .ZN(n415) );
  AOI222_X1 U3598 ( .A1(\UUT/Mpath/the_shift/sh_ror [18]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [18]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [18]), .C2(n6199), .ZN(n2205) );
  AOI22_X1 U3599 ( .A1(\UUT/Mpath/the_shift/sh_sll [18]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [18]), .B2(n6198), .ZN(n2204) );
  NAND3_X1 U3600 ( .A1(n2206), .A2(n2207), .A3(n2208), .ZN(n6134) );
  AOI222_X1 U3601 ( .A1(n1208), .A2(n2209), .B1(\UUT/Mpath/the_alu/diff[18] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[18] ), .C2(n1211), .ZN(n2208)
         );
  INV_X1 U3602 ( .A(\UUT/Mpath/the_alu/N47 ), .ZN(n2209) );
  AOI22_X1 U3603 ( .A1(\UUT/Mpath/the_alu/N139 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N107 ), .B2(n1213), .ZN(n2207) );
  AOI22_X1 U3604 ( .A1(\UUT/Mpath/the_alu/N171 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N203 ), .B2(n1215), .ZN(n2206) );
  INV_X1 U3605 ( .A(n409), .ZN(n2203) );
  NAND4_X1 U3606 ( .A1(n2210), .A2(n2211), .A3(n2212), .A4(n2213), .ZN(n409)
         );
  NOR4_X1 U3607 ( .A1(n2214), .A2(n2215), .A3(n2216), .A4(n2217), .ZN(n2213)
         );
  NAND3_X1 U3608 ( .A1(n6132), .A2(n6131), .A3(n6133), .ZN(n2217) );
  OAI211_X1 U3609 ( .C1(n5560), .C2(n5403), .A(n6129), .B(n6130), .ZN(n2216)
         );
  OAI222_X1 U3610 ( .A1(n5558), .A2(n5275), .B1(n5559), .B2(n5243), .C1(n5561), 
        .C2(n5371), .ZN(n2215) );
  OAI221_X1 U3611 ( .B1(n5531), .B2(n5179), .C1(n5532), .C2(n5211), .A(n2218), 
        .ZN(n2214) );
  AOI22_X1 U3612 ( .A1(n1464), .A2(n1925), .B1(n1465), .B2(n1926), .ZN(n2218)
         );
  INV_X1 U3613 ( .A(n4987), .ZN(n1465) );
  INV_X1 U3614 ( .A(n4955), .ZN(n1464) );
  AOI211_X1 U3615 ( .C1(n1466), .C2(n1927), .A(n2219), .B(n2220), .ZN(n2212)
         );
  OAI22_X1 U3616 ( .A1(n5541), .A2(n4827), .B1(n5551), .B2(n4731), .ZN(n2220)
         );
  OAI222_X1 U3617 ( .A1(n5546), .A2(n4667), .B1(n5552), .B2(n4635), .C1(n5547), 
        .C2(n4699), .ZN(n2219) );
  INV_X1 U3618 ( .A(n4859), .ZN(n1466) );
  AOI221_X1 U3619 ( .B1(n1930), .B2(n1470), .C1(n1931), .C2(n2221), .A(n2222), 
        .ZN(n2211) );
  OAI22_X1 U3620 ( .A1(n4475), .A2(n1934), .B1(n5083), .B2(n1935), .ZN(n2222)
         );
  INV_X1 U3621 ( .A(n5307), .ZN(n2221) );
  INV_X1 U3622 ( .A(n5339), .ZN(n1470) );
  AOI222_X1 U3623 ( .A1(n1472), .A2(n1936), .B1(n1937), .B2(n1473), .C1(n1474), 
        .C2(n1938), .ZN(n2210) );
  INV_X1 U3624 ( .A(n4507), .ZN(n1474) );
  INV_X1 U3625 ( .A(n4443), .ZN(n1473) );
  INV_X1 U3626 ( .A(n4539), .ZN(n1472) );
  AOI222_X1 U3628 ( .A1(n6152), .A2(n5564), .B1(n437), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[17] ), .C2(n5612), .ZN(n5501) );
  NAND2_X1 U3629 ( .A1(n2224), .A2(n2225), .ZN(n437) );
  AOI222_X1 U3630 ( .A1(\UUT/Mpath/the_shift/sh_ror [17]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [17]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [17]), .C2(n6199), .ZN(n2225) );
  AOI22_X1 U3631 ( .A1(\UUT/Mpath/the_shift/sh_sll [17]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [17]), .B2(n6198), .ZN(n2224) );
  NAND3_X1 U3632 ( .A1(n2226), .A2(n2227), .A3(n2228), .ZN(n6152) );
  AOI222_X1 U3633 ( .A1(n1208), .A2(n2229), .B1(\UUT/Mpath/the_alu/diff[17] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[17] ), .C2(n1211), .ZN(n2228)
         );
  INV_X1 U3634 ( .A(\UUT/Mpath/the_alu/N49 ), .ZN(n2229) );
  AOI22_X1 U3635 ( .A1(\UUT/Mpath/the_alu/N140 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N108 ), .B2(n1213), .ZN(n2227) );
  AOI22_X1 U3636 ( .A1(\UUT/Mpath/the_alu/N172 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N204 ), .B2(n1215), .ZN(n2226) );
  INV_X1 U3637 ( .A(n431), .ZN(n2223) );
  NAND4_X1 U3638 ( .A1(n2230), .A2(n2231), .A3(n2232), .A4(n2233), .ZN(n431)
         );
  NOR4_X1 U3639 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2233)
         );
  NAND3_X1 U3640 ( .A1(n6150), .A2(n6149), .A3(n6151), .ZN(n2237) );
  OAI211_X1 U3641 ( .C1(n5560), .C2(n5404), .A(n6147), .B(n6148), .ZN(n2236)
         );
  OAI222_X1 U3642 ( .A1(n5558), .A2(n5276), .B1(n5559), .B2(n5244), .C1(n5561), 
        .C2(n5372), .ZN(n2235) );
  OAI221_X1 U3643 ( .B1(n5531), .B2(n5180), .C1(n5532), .C2(n5212), .A(n2238), 
        .ZN(n2234) );
  AOI22_X1 U3644 ( .A1(n1444), .A2(n1925), .B1(n1445), .B2(n1926), .ZN(n2238)
         );
  INV_X1 U3645 ( .A(n4988), .ZN(n1445) );
  INV_X1 U3646 ( .A(n4956), .ZN(n1444) );
  AOI211_X1 U3647 ( .C1(n1446), .C2(n1927), .A(n2239), .B(n2240), .ZN(n2232)
         );
  OAI22_X1 U3648 ( .A1(n5541), .A2(n4828), .B1(n5551), .B2(n4732), .ZN(n2240)
         );
  OAI222_X1 U3649 ( .A1(n5546), .A2(n4668), .B1(n5552), .B2(n4636), .C1(n5547), 
        .C2(n4700), .ZN(n2239) );
  INV_X1 U3650 ( .A(n4860), .ZN(n1446) );
  AOI221_X1 U3651 ( .B1(n1930), .B2(n1450), .C1(n1931), .C2(n2241), .A(n2242), 
        .ZN(n2231) );
  OAI22_X1 U3652 ( .A1(n4476), .A2(n1934), .B1(n5084), .B2(n6373), .ZN(n2242)
         );
  INV_X1 U3653 ( .A(n5308), .ZN(n2241) );
  INV_X1 U3654 ( .A(n5340), .ZN(n1450) );
  AOI222_X1 U3655 ( .A1(n1452), .A2(n1936), .B1(n1937), .B2(n1453), .C1(n1454), 
        .C2(n1938), .ZN(n2230) );
  INV_X1 U3656 ( .A(n4508), .ZN(n1454) );
  INV_X1 U3657 ( .A(n4444), .ZN(n1453) );
  INV_X1 U3658 ( .A(n4540), .ZN(n1452) );
  AOI222_X1 U3660 ( .A1(n6161), .A2(n5564), .B1(n464), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[16] ), .C2(n5612), .ZN(n5504) );
  NAND2_X1 U3661 ( .A1(n2244), .A2(n2245), .ZN(n464) );
  AOI222_X1 U3662 ( .A1(\UUT/Mpath/the_shift/sh_ror [16]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [16]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [16]), .C2(n6199), .ZN(n2245) );
  AOI22_X1 U3663 ( .A1(\UUT/Mpath/the_shift/sh_sll [16]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [16]), .B2(n6198), .ZN(n2244) );
  NAND3_X1 U3664 ( .A1(n2246), .A2(n2247), .A3(n2248), .ZN(n6161) );
  AOI222_X1 U3665 ( .A1(n1208), .A2(n2249), .B1(\UUT/Mpath/the_alu/diff[16] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[16] ), .C2(n1211), .ZN(n2248)
         );
  INV_X1 U3666 ( .A(\UUT/Mpath/the_alu/N51 ), .ZN(n2249) );
  AOI22_X1 U3667 ( .A1(\UUT/Mpath/the_alu/N141 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N109 ), .B2(n1213), .ZN(n2247) );
  AOI22_X1 U3668 ( .A1(\UUT/Mpath/the_alu/N173 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N205 ), .B2(n1215), .ZN(n2246) );
  INV_X1 U3669 ( .A(n458), .ZN(n2243) );
  NAND4_X1 U3670 ( .A1(n2250), .A2(n2251), .A3(n2252), .A4(n2253), .ZN(n458)
         );
  NOR4_X1 U3671 ( .A1(n2254), .A2(n2255), .A3(n2256), .A4(n2257), .ZN(n2253)
         );
  NAND3_X1 U3672 ( .A1(n6159), .A2(n6158), .A3(n6160), .ZN(n2257) );
  OAI211_X1 U3673 ( .C1(n5560), .C2(n5405), .A(n6156), .B(n6157), .ZN(n2256)
         );
  OAI222_X1 U3674 ( .A1(n5558), .A2(n5277), .B1(n5559), .B2(n5245), .C1(n5561), 
        .C2(n5373), .ZN(n2255) );
  OAI221_X1 U3675 ( .B1(n5531), .B2(n5181), .C1(n5532), .C2(n5213), .A(n2258), 
        .ZN(n2254) );
  AOI22_X1 U3676 ( .A1(n1424), .A2(n1925), .B1(n1425), .B2(n1926), .ZN(n2258)
         );
  INV_X1 U3677 ( .A(n4989), .ZN(n1425) );
  INV_X1 U3678 ( .A(n4957), .ZN(n1424) );
  AOI211_X1 U3679 ( .C1(n1426), .C2(n1927), .A(n2259), .B(n2260), .ZN(n2252)
         );
  OAI22_X1 U3680 ( .A1(n5541), .A2(n4829), .B1(n5551), .B2(n4733), .ZN(n2260)
         );
  OAI222_X1 U3681 ( .A1(n5546), .A2(n4669), .B1(n5552), .B2(n4637), .C1(n5547), 
        .C2(n4701), .ZN(n2259) );
  INV_X1 U3682 ( .A(n4861), .ZN(n1426) );
  AOI221_X1 U3683 ( .B1(n1930), .B2(n1430), .C1(n1931), .C2(n2261), .A(n2262), 
        .ZN(n2251) );
  OAI22_X1 U3684 ( .A1(n4477), .A2(n1934), .B1(n5085), .B2(n6373), .ZN(n2262)
         );
  INV_X1 U3685 ( .A(n5309), .ZN(n2261) );
  INV_X1 U3686 ( .A(n5341), .ZN(n1430) );
  AOI222_X1 U3687 ( .A1(n1432), .A2(n1936), .B1(n1937), .B2(n1433), .C1(n1434), 
        .C2(n1938), .ZN(n2250) );
  INV_X1 U3688 ( .A(n4509), .ZN(n1434) );
  INV_X1 U3689 ( .A(n4445), .ZN(n1433) );
  INV_X1 U3690 ( .A(n4541), .ZN(n1432) );
  AOI222_X1 U3692 ( .A1(n6169), .A2(n5564), .B1(n493), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[15] ), .C2(n5612), .ZN(n5507) );
  NAND2_X1 U3693 ( .A1(n2264), .A2(n2265), .ZN(n493) );
  AOI222_X1 U3694 ( .A1(\UUT/Mpath/the_shift/sh_ror [15]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [15]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [15]), .C2(n6199), .ZN(n2265) );
  AOI22_X1 U3695 ( .A1(\UUT/Mpath/the_shift/sh_sll [15]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [15]), .B2(n6198), .ZN(n2264) );
  NAND3_X1 U3696 ( .A1(n2266), .A2(n2267), .A3(n2268), .ZN(n6169) );
  AOI222_X1 U3697 ( .A1(n1208), .A2(n2269), .B1(\UUT/Mpath/the_alu/diff[15] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[15] ), .C2(n1211), .ZN(n2268)
         );
  INV_X1 U3698 ( .A(\UUT/Mpath/the_alu/N53 ), .ZN(n2269) );
  AOI22_X1 U3699 ( .A1(\UUT/Mpath/the_alu/N142 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N110 ), .B2(n1213), .ZN(n2267) );
  AOI22_X1 U3700 ( .A1(\UUT/Mpath/the_alu/N174 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N206 ), .B2(n1215), .ZN(n2266) );
  INV_X1 U3701 ( .A(n479), .ZN(n2263) );
  NAND4_X1 U3702 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n479)
         );
  NOR4_X1 U3703 ( .A1(n2274), .A2(n2275), .A3(n2276), .A4(n2277), .ZN(n2273)
         );
  NAND3_X1 U3704 ( .A1(n6167), .A2(n6166), .A3(n6168), .ZN(n2277) );
  OAI211_X1 U3705 ( .C1(n5560), .C2(n5406), .A(n6164), .B(n6165), .ZN(n2276)
         );
  OAI222_X1 U3706 ( .A1(n5558), .A2(n5278), .B1(n5559), .B2(n5246), .C1(n5561), 
        .C2(n5374), .ZN(n2275) );
  OAI221_X1 U3707 ( .B1(n5531), .B2(n5182), .C1(n5532), .C2(n5214), .A(n2278), 
        .ZN(n2274) );
  AOI22_X1 U3708 ( .A1(n1404), .A2(n1925), .B1(n1405), .B2(n1926), .ZN(n2278)
         );
  INV_X1 U3709 ( .A(n4990), .ZN(n1405) );
  INV_X1 U3710 ( .A(n4958), .ZN(n1404) );
  AOI211_X1 U3711 ( .C1(n1406), .C2(n1927), .A(n2279), .B(n2280), .ZN(n2272)
         );
  OAI22_X1 U3712 ( .A1(n5541), .A2(n4830), .B1(n5551), .B2(n4734), .ZN(n2280)
         );
  OAI222_X1 U3713 ( .A1(n5546), .A2(n4670), .B1(n5552), .B2(n4638), .C1(n5547), 
        .C2(n4702), .ZN(n2279) );
  INV_X1 U3714 ( .A(n4862), .ZN(n1406) );
  AOI221_X1 U3715 ( .B1(n1930), .B2(n1410), .C1(n1931), .C2(n2281), .A(n2282), 
        .ZN(n2271) );
  OAI22_X1 U3716 ( .A1(n4478), .A2(n1934), .B1(n5086), .B2(n6373), .ZN(n2282)
         );
  INV_X1 U3717 ( .A(n5310), .ZN(n2281) );
  INV_X1 U3718 ( .A(n5342), .ZN(n1410) );
  AOI222_X1 U3719 ( .A1(n1412), .A2(n1936), .B1(n1937), .B2(n1413), .C1(n1414), 
        .C2(n1938), .ZN(n2270) );
  INV_X1 U3720 ( .A(n4510), .ZN(n1414) );
  INV_X1 U3721 ( .A(n4446), .ZN(n1413) );
  INV_X1 U3722 ( .A(n4542), .ZN(n1412) );
  AOI222_X1 U3724 ( .A1(n6180), .A2(n5564), .B1(n518), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[14] ), .C2(n5612), .ZN(n5510) );
  NAND2_X1 U3725 ( .A1(n2284), .A2(n2285), .ZN(n518) );
  AOI222_X1 U3726 ( .A1(\UUT/Mpath/the_shift/sh_ror [14]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [14]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [14]), .C2(n6199), .ZN(n2285) );
  AOI22_X1 U3727 ( .A1(\UUT/Mpath/the_shift/sh_sll [14]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [14]), .B2(n6198), .ZN(n2284) );
  NAND3_X1 U3728 ( .A1(n2286), .A2(n2287), .A3(n2288), .ZN(n6180) );
  AOI222_X1 U3729 ( .A1(n1208), .A2(n2289), .B1(\UUT/Mpath/the_alu/diff[14] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[14] ), .C2(n1211), .ZN(n2288)
         );
  INV_X1 U3730 ( .A(\UUT/Mpath/the_alu/N55 ), .ZN(n2289) );
  AOI22_X1 U3731 ( .A1(\UUT/Mpath/the_alu/N143 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N111 ), .B2(n1213), .ZN(n2287) );
  AOI22_X1 U3732 ( .A1(\UUT/Mpath/the_alu/N175 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N207 ), .B2(n1215), .ZN(n2286) );
  INV_X1 U3733 ( .A(n508), .ZN(n2283) );
  NAND4_X1 U3734 ( .A1(n2290), .A2(n2291), .A3(n2292), .A4(n2293), .ZN(n508)
         );
  NOR4_X1 U3735 ( .A1(n2294), .A2(n2295), .A3(n2296), .A4(n2297), .ZN(n2293)
         );
  NAND3_X1 U3736 ( .A1(n6178), .A2(n6177), .A3(n6179), .ZN(n2297) );
  OAI211_X1 U3737 ( .C1(n5560), .C2(n5407), .A(n6175), .B(n6176), .ZN(n2296)
         );
  OAI222_X1 U3738 ( .A1(n5558), .A2(n5279), .B1(n5559), .B2(n5247), .C1(n5561), 
        .C2(n5375), .ZN(n2295) );
  OAI221_X1 U3739 ( .B1(n5531), .B2(n5183), .C1(n5532), .C2(n5215), .A(n2298), 
        .ZN(n2294) );
  AOI22_X1 U3740 ( .A1(n1384), .A2(n1925), .B1(n1385), .B2(n1926), .ZN(n2298)
         );
  INV_X1 U3741 ( .A(n4991), .ZN(n1385) );
  INV_X1 U3742 ( .A(n4959), .ZN(n1384) );
  AOI211_X1 U3743 ( .C1(n1386), .C2(n1927), .A(n2299), .B(n2300), .ZN(n2292)
         );
  OAI22_X1 U3744 ( .A1(n5541), .A2(n4831), .B1(n5551), .B2(n4735), .ZN(n2300)
         );
  OAI222_X1 U3745 ( .A1(n5546), .A2(n4671), .B1(n5552), .B2(n4639), .C1(n5547), 
        .C2(n4703), .ZN(n2299) );
  INV_X1 U3746 ( .A(n4863), .ZN(n1386) );
  AOI221_X1 U3747 ( .B1(n1930), .B2(n1390), .C1(n1931), .C2(n2301), .A(n2302), 
        .ZN(n2291) );
  OAI22_X1 U3748 ( .A1(n4479), .A2(n1934), .B1(n5087), .B2(n6373), .ZN(n2302)
         );
  INV_X1 U3749 ( .A(n5311), .ZN(n2301) );
  INV_X1 U3750 ( .A(n5343), .ZN(n1390) );
  AOI222_X1 U3751 ( .A1(n1392), .A2(n1936), .B1(n1937), .B2(n1393), .C1(n1394), 
        .C2(n1938), .ZN(n2290) );
  INV_X1 U3752 ( .A(n4511), .ZN(n1394) );
  INV_X1 U3753 ( .A(n4447), .ZN(n1393) );
  INV_X1 U3754 ( .A(n4543), .ZN(n1392) );
  AOI222_X1 U3756 ( .A1(n6187), .A2(n5564), .B1(n543), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[13] ), .C2(n5612), .ZN(n5513) );
  NAND2_X1 U3757 ( .A1(n2304), .A2(n2305), .ZN(n543) );
  AOI222_X1 U3758 ( .A1(\UUT/Mpath/the_shift/sh_ror [13]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [13]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [13]), .C2(n6199), .ZN(n2305) );
  AOI22_X1 U3759 ( .A1(\UUT/Mpath/the_shift/sh_sll [13]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [13]), .B2(n6198), .ZN(n2304) );
  NAND3_X1 U3760 ( .A1(n2306), .A2(n2307), .A3(n2308), .ZN(n6187) );
  AOI222_X1 U3761 ( .A1(n1208), .A2(n2309), .B1(\UUT/Mpath/the_alu/diff[13] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[13] ), .C2(n1211), .ZN(n2308)
         );
  INV_X1 U3762 ( .A(\UUT/Mpath/the_alu/N57 ), .ZN(n2309) );
  AOI22_X1 U3763 ( .A1(\UUT/Mpath/the_alu/N144 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N112 ), .B2(n1213), .ZN(n2307) );
  AOI22_X1 U3764 ( .A1(\UUT/Mpath/the_alu/N176 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N208 ), .B2(n1215), .ZN(n2306) );
  INV_X1 U3765 ( .A(n533), .ZN(n2303) );
  NAND4_X1 U3766 ( .A1(n2310), .A2(n2311), .A3(n2312), .A4(n2313), .ZN(n533)
         );
  NOR4_X1 U3767 ( .A1(n2314), .A2(n2315), .A3(n2316), .A4(n2317), .ZN(n2313)
         );
  NAND3_X1 U3768 ( .A1(n6185), .A2(n6184), .A3(n6186), .ZN(n2317) );
  OAI211_X1 U3769 ( .C1(n5560), .C2(n5408), .A(n6182), .B(n6183), .ZN(n2316)
         );
  OAI222_X1 U3770 ( .A1(n5558), .A2(n5280), .B1(n5559), .B2(n5248), .C1(n5561), 
        .C2(n5376), .ZN(n2315) );
  OAI221_X1 U3771 ( .B1(n5531), .B2(n5184), .C1(n5532), .C2(n5216), .A(n2318), 
        .ZN(n2314) );
  AOI22_X1 U3772 ( .A1(n1364), .A2(n1925), .B1(n1365), .B2(n1926), .ZN(n2318)
         );
  INV_X1 U3773 ( .A(n4992), .ZN(n1365) );
  INV_X1 U3774 ( .A(n4960), .ZN(n1364) );
  AOI211_X1 U3775 ( .C1(n1366), .C2(n1927), .A(n2319), .B(n2320), .ZN(n2312)
         );
  OAI22_X1 U3776 ( .A1(n5541), .A2(n4832), .B1(n5551), .B2(n4736), .ZN(n2320)
         );
  OAI222_X1 U3777 ( .A1(n5546), .A2(n4672), .B1(n5552), .B2(n4640), .C1(n5547), 
        .C2(n4704), .ZN(n2319) );
  INV_X1 U3778 ( .A(n4864), .ZN(n1366) );
  AOI221_X1 U3779 ( .B1(n1930), .B2(n1370), .C1(n1931), .C2(n2321), .A(n2322), 
        .ZN(n2311) );
  OAI22_X1 U3780 ( .A1(n4480), .A2(n1934), .B1(n5088), .B2(n6373), .ZN(n2322)
         );
  INV_X1 U3781 ( .A(n5312), .ZN(n2321) );
  INV_X1 U3782 ( .A(n5344), .ZN(n1370) );
  AOI222_X1 U3783 ( .A1(n1372), .A2(n1936), .B1(n1937), .B2(n1373), .C1(n1374), 
        .C2(n1938), .ZN(n2310) );
  INV_X1 U3784 ( .A(n4512), .ZN(n1374) );
  INV_X1 U3785 ( .A(n4448), .ZN(n1373) );
  INV_X1 U3786 ( .A(n4544), .ZN(n1372) );
  NAND2_X1 U3787 ( .A1(\UUT/Mcontrol/bp_logicB/memory_main ), .A2(n2323), .ZN(
        \UUT/Mcontrol/st_logic/N42 ) );
  INV_X1 U3788 ( .A(\UUT/Mcontrol/bp_logicB/exec_main ), .ZN(n2323) );
  INV_X1 U3789 ( .A(n763), .ZN(\UUT/Mcontrol/Program_counter/N8 ) );
  INV_X1 U3793 ( .A(n764), .ZN(\UUT/break_code[2] ) );
  AOI222_X1 U3796 ( .A1(n6202), .A2(n5564), .B1(n785), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[2] ), .C2(n5612), .ZN(n5459) );
  NAND2_X1 U3797 ( .A1(n2331), .A2(n2332), .ZN(n785) );
  AOI222_X1 U3798 ( .A1(\UUT/Mpath/the_shift/sh_ror [2]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [2]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [2]), .C2(n6199), .ZN(n2332) );
  AOI22_X1 U3799 ( .A1(\UUT/Mpath/the_shift/sh_sll [2]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [2]), .B2(n6198), .ZN(n2331) );
  NAND3_X1 U3800 ( .A1(n2333), .A2(n2334), .A3(n2335), .ZN(n6202) );
  AOI222_X1 U3801 ( .A1(n1208), .A2(n2336), .B1(\UUT/Mpath/the_alu/diff[2] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[2] ), .C2(n1211), .ZN(n2335) );
  INV_X1 U3802 ( .A(\UUT/Mpath/the_alu/N79 ), .ZN(n2336) );
  AOI22_X1 U3803 ( .A1(\UUT/Mpath/the_alu/N155 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N123 ), .B2(n1213), .ZN(n2334) );
  AOI22_X1 U3804 ( .A1(\UUT/Mpath/the_alu/N187 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N219 ), .B2(n1215), .ZN(n2333) );
  INV_X1 U3805 ( .A(n776), .ZN(n2330) );
  NAND4_X1 U3806 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n776)
         );
  NOR4_X1 U3807 ( .A1(n2341), .A2(n2342), .A3(n2343), .A4(n2344), .ZN(n2340)
         );
  NAND3_X1 U3808 ( .A1(n6261), .A2(n6260), .A3(n6262), .ZN(n2344) );
  OAI211_X1 U3809 ( .C1(n5560), .C2(n5390), .A(n6258), .B(n6259), .ZN(n2343)
         );
  OAI222_X1 U3810 ( .A1(n5558), .A2(n5262), .B1(n5559), .B2(n5230), .C1(n5561), 
        .C2(n5358), .ZN(n2342) );
  OAI221_X1 U3811 ( .B1(n5531), .B2(n5166), .C1(n5532), .C2(n5198), .A(n2345), 
        .ZN(n2341) );
  AOI22_X1 U3812 ( .A1(n1724), .A2(n1925), .B1(n1725), .B2(n1926), .ZN(n2345)
         );
  INV_X1 U3813 ( .A(n4974), .ZN(n1725) );
  INV_X1 U3814 ( .A(n4942), .ZN(n1724) );
  AOI211_X1 U3815 ( .C1(n1726), .C2(n1927), .A(n2346), .B(n2347), .ZN(n2339)
         );
  OAI22_X1 U3816 ( .A1(n5541), .A2(n4814), .B1(n5551), .B2(n4718), .ZN(n2347)
         );
  OAI222_X1 U3817 ( .A1(n5546), .A2(n4654), .B1(n5552), .B2(n4622), .C1(n5547), 
        .C2(n4686), .ZN(n2346) );
  INV_X1 U3818 ( .A(n4846), .ZN(n1726) );
  AOI221_X1 U3819 ( .B1(n1930), .B2(n1730), .C1(n1931), .C2(n2348), .A(n2349), 
        .ZN(n2338) );
  OAI22_X1 U3820 ( .A1(n4462), .A2(n1934), .B1(n5070), .B2(n1935), .ZN(n2349)
         );
  INV_X1 U3821 ( .A(n5294), .ZN(n2348) );
  INV_X1 U3822 ( .A(n5326), .ZN(n1730) );
  AOI222_X1 U3823 ( .A1(n1732), .A2(n1936), .B1(n1937), .B2(n1733), .C1(n1734), 
        .C2(n1938), .ZN(n2337) );
  INV_X1 U3824 ( .A(n4494), .ZN(n1734) );
  INV_X1 U3825 ( .A(n4430), .ZN(n1733) );
  INV_X1 U3826 ( .A(n4526), .ZN(n1732) );
  AOI22_X1 U3830 ( .A1(n908), .A2(\UUT/break_code[12] ), .B1(n6715), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [12]), .ZN(n2351) );
  OAI21_X1 U3831 ( .B1(n6035), .B2(n2072), .A(n2352), .ZN(\UUT/break_code[12] ) );
  NAND2_X1 U3832 ( .A1(n6272), .A2(n2074), .ZN(n2352) );
  INV_X1 U3833 ( .A(\UUT/Mcontrol/d_sampled_finstr [12]), .ZN(n6035) );
  AOI222_X1 U3835 ( .A1(n6203), .A2(n5564), .B1(n569), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[12] ), .C2(n5612), .ZN(n5516) );
  NAND2_X1 U3836 ( .A1(n2354), .A2(n2355), .ZN(n569) );
  AOI222_X1 U3837 ( .A1(\UUT/Mpath/the_shift/sh_ror [12]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [12]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [12]), .C2(n6199), .ZN(n2355) );
  AOI22_X1 U3838 ( .A1(\UUT/Mpath/the_shift/sh_sll [12]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [12]), .B2(n6198), .ZN(n2354) );
  NAND3_X1 U3839 ( .A1(n2356), .A2(n2357), .A3(n2358), .ZN(n6203) );
  AOI222_X1 U3840 ( .A1(n1208), .A2(n2359), .B1(\UUT/Mpath/the_alu/diff[12] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[12] ), .C2(n1211), .ZN(n2358)
         );
  INV_X1 U3841 ( .A(\UUT/Mpath/the_alu/N59 ), .ZN(n2359) );
  AOI22_X1 U3842 ( .A1(\UUT/Mpath/the_alu/N145 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N113 ), .B2(n1213), .ZN(n2357) );
  AOI22_X1 U3843 ( .A1(\UUT/Mpath/the_alu/N177 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N209 ), .B2(n1215), .ZN(n2356) );
  INV_X1 U3844 ( .A(n559), .ZN(n2353) );
  NAND4_X1 U3845 ( .A1(n2360), .A2(n2361), .A3(n2362), .A4(n2363), .ZN(n559)
         );
  NOR4_X1 U3846 ( .A1(n2364), .A2(n2365), .A3(n2366), .A4(n2367), .ZN(n2363)
         );
  NAND3_X1 U3847 ( .A1(n6270), .A2(n6269), .A3(n6271), .ZN(n2367) );
  OAI211_X1 U3848 ( .C1(n5560), .C2(n5409), .A(n6267), .B(n6268), .ZN(n2366)
         );
  OAI222_X1 U3849 ( .A1(n5558), .A2(n5281), .B1(n5559), .B2(n5249), .C1(n5561), 
        .C2(n5377), .ZN(n2365) );
  OAI221_X1 U3850 ( .B1(n5531), .B2(n5185), .C1(n5532), .C2(n5217), .A(n2368), 
        .ZN(n2364) );
  AOI22_X1 U3851 ( .A1(n1344), .A2(n1925), .B1(n1345), .B2(n1926), .ZN(n2368)
         );
  INV_X1 U3852 ( .A(n4993), .ZN(n1345) );
  INV_X1 U3853 ( .A(n4961), .ZN(n1344) );
  AOI211_X1 U3854 ( .C1(n1346), .C2(n1927), .A(n2369), .B(n2370), .ZN(n2362)
         );
  OAI22_X1 U3855 ( .A1(n5541), .A2(n4833), .B1(n5551), .B2(n4737), .ZN(n2370)
         );
  OAI222_X1 U3856 ( .A1(n5546), .A2(n4673), .B1(n5552), .B2(n4641), .C1(n5547), 
        .C2(n4705), .ZN(n2369) );
  INV_X1 U3857 ( .A(n4865), .ZN(n1346) );
  AOI221_X1 U3858 ( .B1(n1930), .B2(n1350), .C1(n1931), .C2(n2371), .A(n2372), 
        .ZN(n2361) );
  OAI22_X1 U3859 ( .A1(n4481), .A2(n1934), .B1(n5089), .B2(n6373), .ZN(n2372)
         );
  INV_X1 U3860 ( .A(n5313), .ZN(n2371) );
  INV_X1 U3861 ( .A(n5345), .ZN(n1350) );
  AOI222_X1 U3862 ( .A1(n1352), .A2(n1936), .B1(n1937), .B2(n1353), .C1(n1354), 
        .C2(n1938), .ZN(n2360) );
  INV_X1 U3863 ( .A(n4513), .ZN(n1354) );
  INV_X1 U3864 ( .A(n4449), .ZN(n1353) );
  INV_X1 U3865 ( .A(n4545), .ZN(n1352) );
  AOI22_X1 U3869 ( .A1(n908), .A2(\UUT/break_code[11] ), .B1(n6449), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [11]), .ZN(n2374) );
  OAI21_X1 U3870 ( .B1(n6036), .B2(n2072), .A(n2375), .ZN(\UUT/break_code[11] ) );
  NAND2_X1 U3871 ( .A1(n6278), .A2(n2074), .ZN(n2375) );
  INV_X1 U3872 ( .A(\UUT/Mcontrol/d_sampled_finstr [11]), .ZN(n6036) );
  AOI222_X1 U3874 ( .A1(n6204), .A2(n5564), .B1(n594), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[11] ), .C2(n5612), .ZN(n5519) );
  NAND2_X1 U3875 ( .A1(n2377), .A2(n2378), .ZN(n594) );
  AOI222_X1 U3876 ( .A1(\UUT/Mpath/the_shift/sh_ror [11]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [11]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [11]), .C2(n6199), .ZN(n2378) );
  AOI22_X1 U3877 ( .A1(\UUT/Mpath/the_shift/sh_sll [11]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [11]), .B2(n6198), .ZN(n2377) );
  NAND3_X1 U3878 ( .A1(n2379), .A2(n2380), .A3(n2381), .ZN(n6204) );
  AOI222_X1 U3879 ( .A1(n1208), .A2(n2382), .B1(\UUT/Mpath/the_alu/diff[11] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[11] ), .C2(n1211), .ZN(n2381)
         );
  INV_X1 U3880 ( .A(\UUT/Mpath/the_alu/N61 ), .ZN(n2382) );
  AOI22_X1 U3881 ( .A1(\UUT/Mpath/the_alu/N146 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N114 ), .B2(n1213), .ZN(n2380) );
  AOI22_X1 U3882 ( .A1(\UUT/Mpath/the_alu/N178 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N210 ), .B2(n1215), .ZN(n2379) );
  INV_X1 U3883 ( .A(n584), .ZN(n2376) );
  NAND4_X1 U3884 ( .A1(n2383), .A2(n2384), .A3(n2385), .A4(n2386), .ZN(n584)
         );
  NOR4_X1 U3885 ( .A1(n2387), .A2(n2388), .A3(n2389), .A4(n2390), .ZN(n2386)
         );
  NAND3_X1 U3886 ( .A1(n6276), .A2(n6275), .A3(n6277), .ZN(n2390) );
  OAI211_X1 U3887 ( .C1(n5560), .C2(n5410), .A(n6273), .B(n6274), .ZN(n2389)
         );
  OAI222_X1 U3888 ( .A1(n5558), .A2(n5282), .B1(n5559), .B2(n5250), .C1(n5561), 
        .C2(n5378), .ZN(n2388) );
  OAI221_X1 U3889 ( .B1(n5531), .B2(n5186), .C1(n5532), .C2(n5218), .A(n2391), 
        .ZN(n2387) );
  AOI22_X1 U3890 ( .A1(n1324), .A2(n1925), .B1(n1325), .B2(n1926), .ZN(n2391)
         );
  INV_X1 U3891 ( .A(n4994), .ZN(n1325) );
  INV_X1 U3892 ( .A(n4962), .ZN(n1324) );
  AOI211_X1 U3893 ( .C1(n1326), .C2(n1927), .A(n2392), .B(n2393), .ZN(n2385)
         );
  OAI22_X1 U3894 ( .A1(n5541), .A2(n4834), .B1(n5551), .B2(n4738), .ZN(n2393)
         );
  OAI222_X1 U3895 ( .A1(n5546), .A2(n4674), .B1(n5552), .B2(n4642), .C1(n5547), 
        .C2(n4706), .ZN(n2392) );
  INV_X1 U3896 ( .A(n4866), .ZN(n1326) );
  AOI221_X1 U3897 ( .B1(n1930), .B2(n1330), .C1(n1931), .C2(n2394), .A(n2395), 
        .ZN(n2384) );
  OAI22_X1 U3898 ( .A1(n4482), .A2(n1934), .B1(n5090), .B2(n6373), .ZN(n2395)
         );
  INV_X1 U3899 ( .A(n5314), .ZN(n2394) );
  INV_X1 U3900 ( .A(n5346), .ZN(n1330) );
  AOI222_X1 U3901 ( .A1(n1332), .A2(n1936), .B1(n1937), .B2(n1333), .C1(n1334), 
        .C2(n1938), .ZN(n2383) );
  INV_X1 U3902 ( .A(n4514), .ZN(n1334) );
  INV_X1 U3903 ( .A(n4450), .ZN(n1333) );
  INV_X1 U3904 ( .A(n4546), .ZN(n1332) );
  INV_X1 U3905 ( .A(n979), .ZN(\UUT/Mcontrol/Program_counter/N24 ) );
  OAI21_X1 U3909 ( .B1(n5881), .B2(n2072), .A(n2398), .ZN(\UUT/break_code[10] ) );
  NAND2_X1 U3910 ( .A1(n6327), .A2(n2074), .ZN(n2398) );
  INV_X1 U3911 ( .A(\UUT/Mcontrol/d_sampled_finstr [10]), .ZN(n5881) );
  AOI222_X1 U3913 ( .A1(n6205), .A2(n5564), .B1(n1162), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[10] ), .C2(n5612), .ZN(n5522) );
  NAND2_X1 U3914 ( .A1(n2400), .A2(n2401), .ZN(n1162) );
  AOI222_X1 U3915 ( .A1(\UUT/Mpath/the_shift/sh_ror [10]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [10]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [10]), .C2(n6199), .ZN(n2401) );
  AOI22_X1 U3916 ( .A1(\UUT/Mpath/the_shift/sh_sll [10]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [10]), .B2(n6198), .ZN(n2400) );
  NAND3_X1 U3917 ( .A1(n2402), .A2(n2403), .A3(n2404), .ZN(n6205) );
  AOI222_X1 U3918 ( .A1(n1208), .A2(n2405), .B1(\UUT/Mpath/the_alu/diff[10] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[10] ), .C2(n1211), .ZN(n2404)
         );
  INV_X1 U3919 ( .A(\UUT/Mpath/the_alu/N63 ), .ZN(n2405) );
  AOI22_X1 U3920 ( .A1(\UUT/Mpath/the_alu/N147 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N115 ), .B2(n1213), .ZN(n2403) );
  AOI22_X1 U3921 ( .A1(\UUT/Mpath/the_alu/N179 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N211 ), .B2(n1215), .ZN(n2402) );
  INV_X1 U3922 ( .A(n604), .ZN(n2399) );
  NAND4_X1 U3923 ( .A1(n2406), .A2(n2407), .A3(n2408), .A4(n2409), .ZN(n604)
         );
  NOR4_X1 U3924 ( .A1(n2410), .A2(n2411), .A3(n2412), .A4(n2413), .ZN(n2409)
         );
  NAND3_X1 U3925 ( .A1(n6282), .A2(n6281), .A3(n6283), .ZN(n2413) );
  OAI211_X1 U3926 ( .C1(n5560), .C2(n5411), .A(n6279), .B(n6280), .ZN(n2412)
         );
  OAI222_X1 U3927 ( .A1(n5558), .A2(n5283), .B1(n5559), .B2(n5251), .C1(n5561), 
        .C2(n5379), .ZN(n2411) );
  OAI221_X1 U3928 ( .B1(n5531), .B2(n5187), .C1(n5532), .C2(n5219), .A(n2414), 
        .ZN(n2410) );
  AOI22_X1 U3929 ( .A1(n1304), .A2(n1925), .B1(n1305), .B2(n1926), .ZN(n2414)
         );
  INV_X1 U3930 ( .A(n4995), .ZN(n1305) );
  INV_X1 U3931 ( .A(n4963), .ZN(n1304) );
  AOI211_X1 U3932 ( .C1(n1306), .C2(n1927), .A(n2415), .B(n2416), .ZN(n2408)
         );
  OAI22_X1 U3933 ( .A1(n5541), .A2(n4835), .B1(n5551), .B2(n4739), .ZN(n2416)
         );
  OAI222_X1 U3934 ( .A1(n5546), .A2(n4675), .B1(n5552), .B2(n4643), .C1(n5547), 
        .C2(n4707), .ZN(n2415) );
  INV_X1 U3935 ( .A(n4867), .ZN(n1306) );
  AOI221_X1 U3936 ( .B1(n1930), .B2(n1310), .C1(n1931), .C2(n2417), .A(n2418), 
        .ZN(n2407) );
  OAI22_X1 U3937 ( .A1(n4483), .A2(n1934), .B1(n5091), .B2(n6373), .ZN(n2418)
         );
  INV_X1 U3938 ( .A(n5315), .ZN(n2417) );
  INV_X1 U3939 ( .A(n5347), .ZN(n1310) );
  AOI222_X1 U3940 ( .A1(n1312), .A2(n1936), .B1(n1937), .B2(n1313), .C1(n1314), 
        .C2(n1938), .ZN(n2406) );
  INV_X1 U3941 ( .A(n4515), .ZN(n1314) );
  INV_X1 U3942 ( .A(n4451), .ZN(n1313) );
  INV_X1 U3943 ( .A(n4547), .ZN(n1312) );
  INV_X1 U3944 ( .A(n909), .ZN(\UUT/Mcontrol/Program_counter/N22 ) );
  OAI21_X1 U3948 ( .B1(n5889), .B2(n2072), .A(n2421), .ZN(\UUT/break_code[9] )
         );
  NAND2_X1 U3949 ( .A1(n6216), .A2(n2074), .ZN(n2421) );
  INV_X1 U3950 ( .A(\UUT/Mcontrol/d_sampled_finstr [9]), .ZN(n5889) );
  OAI222_X1 U3951 ( .A1(n5433), .A2(n5530), .B1(n5529), .B2(n2422), .C1(n5528), 
        .C2(n5429), .ZN(\UUT/branch_rega [9]) );
  AOI222_X1 U3952 ( .A1(n6189), .A2(n5564), .B1(n629), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[9] ), .C2(n5612), .ZN(n5429) );
  NAND2_X1 U3953 ( .A1(n2423), .A2(n2424), .ZN(n629) );
  AOI222_X1 U3954 ( .A1(\UUT/Mpath/the_shift/sh_ror [9]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [9]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [9]), .C2(n6199), .ZN(n2424) );
  AOI22_X1 U3955 ( .A1(\UUT/Mpath/the_shift/sh_sll [9]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [9]), .B2(n6198), .ZN(n2423) );
  NAND3_X1 U3956 ( .A1(n2425), .A2(n2426), .A3(n2427), .ZN(n6189) );
  AOI222_X1 U3957 ( .A1(n1208), .A2(n2428), .B1(\UUT/Mpath/the_alu/diff[9] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[9] ), .C2(n1211), .ZN(n2427) );
  INV_X1 U3958 ( .A(\UUT/Mpath/the_alu/N65 ), .ZN(n2428) );
  AOI22_X1 U3959 ( .A1(\UUT/Mpath/the_alu/N148 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N116 ), .B2(n1213), .ZN(n2426) );
  AOI22_X1 U3960 ( .A1(\UUT/Mpath/the_alu/N180 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N212 ), .B2(n1215), .ZN(n2425) );
  INV_X1 U3961 ( .A(n619), .ZN(n2422) );
  NAND4_X1 U3962 ( .A1(n2429), .A2(n2430), .A3(n2431), .A4(n2432), .ZN(n619)
         );
  NOR4_X1 U3963 ( .A1(n2433), .A2(n2434), .A3(n2435), .A4(n2436), .ZN(n2432)
         );
  NAND3_X1 U3964 ( .A1(n6214), .A2(n6213), .A3(n6215), .ZN(n2436) );
  OAI211_X1 U3965 ( .C1(n5560), .C2(n5381), .A(n6211), .B(n6212), .ZN(n2435)
         );
  OAI222_X1 U3966 ( .A1(n5558), .A2(n5253), .B1(n5559), .B2(n5221), .C1(n5561), 
        .C2(n5349), .ZN(n2434) );
  OAI221_X1 U3967 ( .B1(n5531), .B2(n5157), .C1(n5532), .C2(n5189), .A(n2437), 
        .ZN(n2433) );
  AOI22_X1 U3968 ( .A1(n1904), .A2(n1925), .B1(n1905), .B2(n1926), .ZN(n2437)
         );
  INV_X1 U3969 ( .A(n4965), .ZN(n1905) );
  INV_X1 U3970 ( .A(n4933), .ZN(n1904) );
  AOI211_X1 U3971 ( .C1(n1906), .C2(n1927), .A(n2438), .B(n2439), .ZN(n2431)
         );
  OAI22_X1 U3972 ( .A1(n5541), .A2(n4805), .B1(n5551), .B2(n4709), .ZN(n2439)
         );
  OAI222_X1 U3973 ( .A1(n5546), .A2(n4645), .B1(n5552), .B2(n4613), .C1(n5547), 
        .C2(n4677), .ZN(n2438) );
  INV_X1 U3974 ( .A(n4837), .ZN(n1906) );
  AOI221_X1 U3975 ( .B1(n1930), .B2(n1910), .C1(n1931), .C2(n2440), .A(n2441), 
        .ZN(n2430) );
  OAI22_X1 U3976 ( .A1(n4453), .A2(n1934), .B1(n5061), .B2(n6373), .ZN(n2441)
         );
  INV_X1 U3977 ( .A(n5285), .ZN(n2440) );
  INV_X1 U3978 ( .A(n5317), .ZN(n1910) );
  AOI222_X1 U3979 ( .A1(n1913), .A2(n1936), .B1(n1937), .B2(n1914), .C1(n1915), 
        .C2(n1938), .ZN(n2429) );
  INV_X1 U3980 ( .A(n4485), .ZN(n1915) );
  INV_X1 U3981 ( .A(n4421), .ZN(n1914) );
  INV_X1 U3982 ( .A(n4517), .ZN(n1913) );
  INV_X1 U3983 ( .A(n631), .ZN(\UUT/Mcontrol/Program_counter/N20 ) );
  AOI22_X1 U3986 ( .A1(n908), .A2(\UUT/break_code[8] ), .B1(n906), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [8]), .ZN(n2443) );
  OAI21_X1 U3987 ( .B1(n5897), .B2(n2072), .A(n2444), .ZN(\UUT/break_code[8] )
         );
  NAND2_X1 U3988 ( .A1(n6222), .A2(n2074), .ZN(n2444) );
  INV_X1 U3989 ( .A(\UUT/Mcontrol/d_sampled_finstr [8]), .ZN(n5897) );
  AOI222_X1 U3991 ( .A1(n6190), .A2(n5564), .B1(n1153), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[8] ), .C2(n5612), .ZN(n5435) );
  NAND2_X1 U3992 ( .A1(n2446), .A2(n2447), .ZN(n1153) );
  AOI222_X1 U3993 ( .A1(\UUT/Mpath/the_shift/sh_ror [8]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [8]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [8]), .C2(n6199), .ZN(n2447) );
  AOI22_X1 U3994 ( .A1(\UUT/Mpath/the_shift/sh_sll [8]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [8]), .B2(n6198), .ZN(n2446) );
  NAND3_X1 U3995 ( .A1(n2448), .A2(n2449), .A3(n2450), .ZN(n6190) );
  AOI222_X1 U3996 ( .A1(n1208), .A2(n2451), .B1(\UUT/Mpath/the_alu/diff[8] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[8] ), .C2(n1211), .ZN(n2450) );
  INV_X1 U3997 ( .A(\UUT/Mpath/the_alu/N67 ), .ZN(n2451) );
  AOI22_X1 U3998 ( .A1(\UUT/Mpath/the_alu/N149 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N117 ), .B2(n1213), .ZN(n2449) );
  AOI22_X1 U3999 ( .A1(\UUT/Mpath/the_alu/N181 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N213 ), .B2(n1215), .ZN(n2448) );
  INV_X1 U4000 ( .A(n640), .ZN(n2445) );
  NAND4_X1 U4001 ( .A1(n2452), .A2(n2453), .A3(n2454), .A4(n2455), .ZN(n640)
         );
  NOR4_X1 U4002 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  NAND3_X1 U4003 ( .A1(n6220), .A2(n6219), .A3(n6221), .ZN(n2459) );
  OAI211_X1 U4004 ( .C1(n5560), .C2(n5382), .A(n6217), .B(n6218), .ZN(n2458)
         );
  OAI222_X1 U4005 ( .A1(n5558), .A2(n5254), .B1(n5559), .B2(n5222), .C1(n5561), 
        .C2(n5350), .ZN(n2457) );
  OAI221_X1 U4006 ( .B1(n5531), .B2(n5158), .C1(n5532), .C2(n5190), .A(n2460), 
        .ZN(n2456) );
  AOI22_X1 U4007 ( .A1(n1884), .A2(n1925), .B1(n1885), .B2(n1926), .ZN(n2460)
         );
  INV_X1 U4008 ( .A(n4966), .ZN(n1885) );
  INV_X1 U4009 ( .A(n4934), .ZN(n1884) );
  AOI211_X1 U4010 ( .C1(n1886), .C2(n1927), .A(n2461), .B(n2462), .ZN(n2454)
         );
  OAI22_X1 U4011 ( .A1(n5541), .A2(n4806), .B1(n5551), .B2(n4710), .ZN(n2462)
         );
  OAI222_X1 U4012 ( .A1(n5546), .A2(n4646), .B1(n5552), .B2(n4614), .C1(n5547), 
        .C2(n4678), .ZN(n2461) );
  INV_X1 U4013 ( .A(n4838), .ZN(n1886) );
  AOI221_X1 U4014 ( .B1(n1930), .B2(n1890), .C1(n1931), .C2(n2463), .A(n2464), 
        .ZN(n2453) );
  OAI22_X1 U4015 ( .A1(n4454), .A2(n1934), .B1(n5062), .B2(n1935), .ZN(n2464)
         );
  INV_X1 U4016 ( .A(n5286), .ZN(n2463) );
  INV_X1 U4017 ( .A(n5318), .ZN(n1890) );
  AOI222_X1 U4018 ( .A1(n1892), .A2(n1936), .B1(n1937), .B2(n1893), .C1(n1894), 
        .C2(n1938), .ZN(n2452) );
  INV_X1 U4019 ( .A(n4486), .ZN(n1894) );
  INV_X1 U4020 ( .A(n4422), .ZN(n1893) );
  INV_X1 U4021 ( .A(n4518), .ZN(n1892) );
  AOI22_X1 U4025 ( .A1(n908), .A2(\UUT/break_code[7] ), .B1(n906), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [7]), .ZN(n2466) );
  OAI21_X1 U4026 ( .B1(n6094), .B2(n2072), .A(n2467), .ZN(\UUT/break_code[7] )
         );
  NAND2_X1 U4027 ( .A1(n6228), .A2(n2074), .ZN(n2467) );
  INV_X1 U4028 ( .A(\UUT/Mcontrol/d_sampled_finstr [7]), .ZN(n6094) );
  AOI222_X1 U4030 ( .A1(n6191), .A2(n5564), .B1(n664), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[7] ), .C2(n5612), .ZN(n5438) );
  NAND2_X1 U4031 ( .A1(n2469), .A2(n2470), .ZN(n664) );
  AOI222_X1 U4032 ( .A1(\UUT/Mpath/the_shift/sh_ror [7]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [7]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [7]), .C2(n6199), .ZN(n2470) );
  AOI22_X1 U4033 ( .A1(\UUT/Mpath/the_shift/sh_sll [7]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [7]), .B2(n6198), .ZN(n2469) );
  NAND3_X1 U4034 ( .A1(n2471), .A2(n2472), .A3(n2473), .ZN(n6191) );
  AOI222_X1 U4035 ( .A1(n1208), .A2(n2474), .B1(\UUT/Mpath/the_alu/diff[7] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[7] ), .C2(n1211), .ZN(n2473) );
  INV_X1 U4036 ( .A(\UUT/Mpath/the_alu/N69 ), .ZN(n2474) );
  AOI22_X1 U4037 ( .A1(\UUT/Mpath/the_alu/N150 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N118 ), .B2(n1213), .ZN(n2472) );
  AOI22_X1 U4038 ( .A1(\UUT/Mpath/the_alu/N182 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N214 ), .B2(n1215), .ZN(n2471) );
  INV_X1 U4039 ( .A(n656), .ZN(n2468) );
  NAND4_X1 U4040 ( .A1(n2475), .A2(n2476), .A3(n2477), .A4(n2478), .ZN(n656)
         );
  NOR4_X1 U4041 ( .A1(n2479), .A2(n2480), .A3(n2481), .A4(n2482), .ZN(n2478)
         );
  NAND3_X1 U4042 ( .A1(n6226), .A2(n6225), .A3(n6227), .ZN(n2482) );
  OAI211_X1 U4043 ( .C1(n5560), .C2(n5383), .A(n6223), .B(n6224), .ZN(n2481)
         );
  OAI222_X1 U4044 ( .A1(n5558), .A2(n5255), .B1(n5559), .B2(n5223), .C1(n5561), 
        .C2(n5351), .ZN(n2480) );
  OAI221_X1 U4045 ( .B1(n5531), .B2(n5159), .C1(n5532), .C2(n5191), .A(n2483), 
        .ZN(n2479) );
  AOI22_X1 U4046 ( .A1(n1864), .A2(n1925), .B1(n1865), .B2(n1926), .ZN(n2483)
         );
  INV_X1 U4047 ( .A(n4967), .ZN(n1865) );
  INV_X1 U4048 ( .A(n4935), .ZN(n1864) );
  AOI211_X1 U4049 ( .C1(n1866), .C2(n1927), .A(n2484), .B(n2485), .ZN(n2477)
         );
  OAI22_X1 U4050 ( .A1(n5541), .A2(n4807), .B1(n5551), .B2(n4711), .ZN(n2485)
         );
  OAI222_X1 U4051 ( .A1(n5546), .A2(n4647), .B1(n5552), .B2(n4615), .C1(n5547), 
        .C2(n4679), .ZN(n2484) );
  INV_X1 U4052 ( .A(n4839), .ZN(n1866) );
  AOI221_X1 U4053 ( .B1(n1930), .B2(n1870), .C1(n1931), .C2(n2486), .A(n2487), 
        .ZN(n2476) );
  OAI22_X1 U4054 ( .A1(n4455), .A2(n1934), .B1(n5063), .B2(n6373), .ZN(n2487)
         );
  INV_X1 U4055 ( .A(n5287), .ZN(n2486) );
  INV_X1 U4056 ( .A(n5319), .ZN(n1870) );
  AOI222_X1 U4057 ( .A1(n1872), .A2(n1936), .B1(n1937), .B2(n1873), .C1(n1874), 
        .C2(n1938), .ZN(n2475) );
  INV_X1 U4058 ( .A(n4487), .ZN(n1874) );
  INV_X1 U4059 ( .A(n4423), .ZN(n1873) );
  INV_X1 U4060 ( .A(n4519), .ZN(n1872) );
  AOI22_X1 U4064 ( .A1(n908), .A2(\UUT/break_code[6] ), .B1(n906), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [6]), .ZN(n2489) );
  OAI21_X1 U4065 ( .B1(n6143), .B2(n2072), .A(n2490), .ZN(\UUT/break_code[6] )
         );
  NAND2_X1 U4066 ( .A1(n6234), .A2(n2074), .ZN(n2490) );
  INV_X1 U4067 ( .A(\UUT/Mcontrol/d_sampled_finstr [6]), .ZN(n6143) );
  AOI222_X1 U4069 ( .A1(n6192), .A2(n5564), .B1(n692), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[6] ), .C2(n5612), .ZN(n5441) );
  NAND2_X1 U4070 ( .A1(n2492), .A2(n2493), .ZN(n692) );
  AOI222_X1 U4071 ( .A1(\UUT/Mpath/the_shift/sh_ror [6]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [6]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [6]), .C2(n6199), .ZN(n2493) );
  AOI22_X1 U4072 ( .A1(\UUT/Mpath/the_shift/sh_sll [6]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [6]), .B2(n6198), .ZN(n2492) );
  NAND3_X1 U4073 ( .A1(n2494), .A2(n2495), .A3(n2496), .ZN(n6192) );
  AOI222_X1 U4074 ( .A1(n1208), .A2(n2497), .B1(\UUT/Mpath/the_alu/diff[6] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[6] ), .C2(n1211), .ZN(n2496) );
  INV_X1 U4075 ( .A(\UUT/Mpath/the_alu/N71 ), .ZN(n2497) );
  AOI22_X1 U4076 ( .A1(\UUT/Mpath/the_alu/N151 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N119 ), .B2(n1213), .ZN(n2495) );
  AOI22_X1 U4077 ( .A1(\UUT/Mpath/the_alu/N183 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N215 ), .B2(n1215), .ZN(n2494) );
  INV_X1 U4078 ( .A(n679), .ZN(n2491) );
  NAND4_X1 U4079 ( .A1(n2498), .A2(n2499), .A3(n2500), .A4(n2501), .ZN(n679)
         );
  NOR4_X1 U4080 ( .A1(n2502), .A2(n2503), .A3(n2504), .A4(n2505), .ZN(n2501)
         );
  NAND3_X1 U4081 ( .A1(n6232), .A2(n6231), .A3(n6233), .ZN(n2505) );
  OAI211_X1 U4082 ( .C1(n5560), .C2(n5384), .A(n6229), .B(n6230), .ZN(n2504)
         );
  OAI222_X1 U4083 ( .A1(n5558), .A2(n5256), .B1(n5559), .B2(n5224), .C1(n5561), 
        .C2(n5352), .ZN(n2503) );
  OAI221_X1 U4084 ( .B1(n5531), .B2(n5160), .C1(n5532), .C2(n5192), .A(n2506), 
        .ZN(n2502) );
  AOI22_X1 U4085 ( .A1(n1844), .A2(n1925), .B1(n1845), .B2(n1926), .ZN(n2506)
         );
  INV_X1 U4086 ( .A(n4968), .ZN(n1845) );
  INV_X1 U4087 ( .A(n4936), .ZN(n1844) );
  AOI211_X1 U4088 ( .C1(n1846), .C2(n1927), .A(n2507), .B(n2508), .ZN(n2500)
         );
  OAI22_X1 U4089 ( .A1(n5541), .A2(n4808), .B1(n5551), .B2(n4712), .ZN(n2508)
         );
  OAI222_X1 U4090 ( .A1(n5546), .A2(n4648), .B1(n5552), .B2(n4616), .C1(n5547), 
        .C2(n4680), .ZN(n2507) );
  INV_X1 U4091 ( .A(n4840), .ZN(n1846) );
  AOI221_X1 U4092 ( .B1(n1930), .B2(n1850), .C1(n1931), .C2(n2509), .A(n2510), 
        .ZN(n2499) );
  OAI22_X1 U4093 ( .A1(n4456), .A2(n1934), .B1(n5064), .B2(n6373), .ZN(n2510)
         );
  INV_X1 U4094 ( .A(n5288), .ZN(n2509) );
  INV_X1 U4095 ( .A(n5320), .ZN(n1850) );
  AOI222_X1 U4096 ( .A1(n1852), .A2(n1936), .B1(n1937), .B2(n1853), .C1(n1854), 
        .C2(n1938), .ZN(n2498) );
  INV_X1 U4097 ( .A(n4488), .ZN(n1854) );
  INV_X1 U4098 ( .A(n4424), .ZN(n1853) );
  INV_X1 U4099 ( .A(n4520), .ZN(n1852) );
  OAI21_X1 U4104 ( .B1(n5423), .B2(n2072), .A(n2513), .ZN(\UUT/break_code[5] )
         );
  NAND2_X1 U4105 ( .A1(n6240), .A2(n2074), .ZN(n2513) );
  OAI21_X1 U4107 ( .B1(n6170), .B2(n2514), .A(n6030), .ZN(n2072) );
  NOR2_X1 U4108 ( .A1(n2070), .A2(n445), .ZN(n2514) );
  INV_X1 U4109 ( .A(n6209), .ZN(n445) );
  INV_X1 U4110 ( .A(n6172), .ZN(n2070) );
  NAND2_X1 U4111 ( .A1(n932), .A2(n929), .ZN(n6170) );
  NOR2_X1 U4112 ( .A1(n2077), .A2(n1219), .ZN(n929) );
  OAI21_X1 U4113 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2071 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A(
        \UUT/Mcontrol/Operation_decoding32/N2066 ), .ZN(n1219) );
  NAND2_X1 U4114 ( .A1(n915), .A2(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
        .ZN(n2077) );
  INV_X1 U4115 ( .A(\UUT/Mcontrol/Operation_decoding32/N2079 ), .ZN(n915) );
  NOR2_X1 U4116 ( .A1(n1004), .A2(\UUT/Mcontrol/Operation_decoding32/N2061 ), 
        .ZN(n932) );
  NAND2_X1 U4117 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2054 ), .A2(n924), 
        .ZN(n1004) );
  OR2_X1 U4118 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2047 ), .ZN(n924) );
  INV_X1 U4119 ( .A(\UUT/Mcontrol/d_sampled_finstr [5]), .ZN(n5423) );
  OAI222_X1 U4120 ( .A1(n5446), .A2(n5530), .B1(n5529), .B2(n2515), .C1(n5528), 
        .C2(n5444), .ZN(\UUT/branch_rega [5]) );
  AOI222_X1 U4121 ( .A1(n6193), .A2(n5564), .B1(n715), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[5] ), .C2(n5612), .ZN(n5444) );
  NAND2_X1 U4122 ( .A1(n2516), .A2(n2517), .ZN(n715) );
  AOI222_X1 U4123 ( .A1(\UUT/Mpath/the_shift/sh_ror [5]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [5]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [5]), .C2(n6199), .ZN(n2517) );
  AOI22_X1 U4124 ( .A1(\UUT/Mpath/the_shift/sh_sll [5]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [5]), .B2(n6198), .ZN(n2516) );
  NAND3_X1 U4125 ( .A1(n2518), .A2(n2519), .A3(n2520), .ZN(n6193) );
  AOI222_X1 U4126 ( .A1(n1208), .A2(n2521), .B1(\UUT/Mpath/the_alu/diff[5] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[5] ), .C2(n1211), .ZN(n2520) );
  INV_X1 U4127 ( .A(\UUT/Mpath/the_alu/N73 ), .ZN(n2521) );
  AOI22_X1 U4128 ( .A1(\UUT/Mpath/the_alu/N152 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N120 ), .B2(n1213), .ZN(n2519) );
  AOI22_X1 U4129 ( .A1(\UUT/Mpath/the_alu/N184 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N216 ), .B2(n1215), .ZN(n2518) );
  INV_X1 U4130 ( .A(n707), .ZN(n2515) );
  NAND4_X1 U4131 ( .A1(n2522), .A2(n2523), .A3(n2524), .A4(n2525), .ZN(n707)
         );
  NOR4_X1 U4132 ( .A1(n2526), .A2(n2527), .A3(n2528), .A4(n2529), .ZN(n2525)
         );
  NAND3_X1 U4133 ( .A1(n6238), .A2(n6237), .A3(n6239), .ZN(n2529) );
  OAI211_X1 U4134 ( .C1(n5560), .C2(n5385), .A(n6235), .B(n6236), .ZN(n2528)
         );
  OAI222_X1 U4135 ( .A1(n5558), .A2(n5257), .B1(n5559), .B2(n5225), .C1(n5561), 
        .C2(n5353), .ZN(n2527) );
  OAI221_X1 U4136 ( .B1(n5531), .B2(n5161), .C1(n5532), .C2(n5193), .A(n2530), 
        .ZN(n2526) );
  AOI22_X1 U4137 ( .A1(n1824), .A2(n1925), .B1(n1825), .B2(n1926), .ZN(n2530)
         );
  INV_X1 U4138 ( .A(n4969), .ZN(n1825) );
  INV_X1 U4139 ( .A(n4937), .ZN(n1824) );
  AOI211_X1 U4140 ( .C1(n1826), .C2(n1927), .A(n2531), .B(n2532), .ZN(n2524)
         );
  OAI22_X1 U4141 ( .A1(n5541), .A2(n4809), .B1(n5551), .B2(n4713), .ZN(n2532)
         );
  OAI222_X1 U4142 ( .A1(n5546), .A2(n4649), .B1(n5552), .B2(n4617), .C1(n5547), 
        .C2(n4681), .ZN(n2531) );
  INV_X1 U4143 ( .A(n4841), .ZN(n1826) );
  AOI221_X1 U4144 ( .B1(n1930), .B2(n1830), .C1(n1931), .C2(n2533), .A(n2534), 
        .ZN(n2523) );
  OAI22_X1 U4145 ( .A1(n4457), .A2(n1934), .B1(n5065), .B2(n1935), .ZN(n2534)
         );
  INV_X1 U4146 ( .A(n5289), .ZN(n2533) );
  INV_X1 U4147 ( .A(n5321), .ZN(n1830) );
  AOI222_X1 U4148 ( .A1(n1832), .A2(n1936), .B1(n1937), .B2(n1833), .C1(n1834), 
        .C2(n1938), .ZN(n2522) );
  INV_X1 U4149 ( .A(n4489), .ZN(n1834) );
  INV_X1 U4150 ( .A(n4425), .ZN(n1833) );
  INV_X1 U4151 ( .A(n4521), .ZN(n1832) );
  INV_X1 U4156 ( .A(n718), .ZN(\UUT/break_code[4] ) );
  AOI22_X1 U4157 ( .A1(n6247), .A2(n2328), .B1(n2329), .B2(
        \UUT/Mcontrol/d_sampled_finstr [4]), .ZN(n718) );
  OAI222_X1 U4158 ( .A1(n5449), .A2(n5530), .B1(n5529), .B2(n2537), .C1(n5528), 
        .C2(n5447), .ZN(\UUT/branch_rega [4]) );
  AOI222_X1 U4159 ( .A1(n6194), .A2(n5564), .B1(n738), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[4] ), .C2(n5612), .ZN(n5447) );
  NAND2_X1 U4160 ( .A1(n2538), .A2(n2539), .ZN(n738) );
  AOI222_X1 U4161 ( .A1(\UUT/Mpath/the_shift/sh_ror [4]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [4]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [4]), .C2(n6199), .ZN(n2539) );
  AOI22_X1 U4162 ( .A1(\UUT/Mpath/the_shift/sh_sll [4]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [4]), .B2(n6198), .ZN(n2538) );
  NAND3_X1 U4163 ( .A1(n2540), .A2(n2541), .A3(n2542), .ZN(n6194) );
  AOI222_X1 U4164 ( .A1(n1208), .A2(n2543), .B1(\UUT/Mpath/the_alu/diff[4] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[4] ), .C2(n1211), .ZN(n2542) );
  INV_X1 U4165 ( .A(\UUT/Mpath/the_alu/N75 ), .ZN(n2543) );
  AOI22_X1 U4166 ( .A1(\UUT/Mpath/the_alu/N153 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N121 ), .B2(n1213), .ZN(n2541) );
  AOI22_X1 U4167 ( .A1(\UUT/Mpath/the_alu/N185 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N217 ), .B2(n1215), .ZN(n2540) );
  INV_X1 U4168 ( .A(n730), .ZN(n2537) );
  NAND4_X1 U4169 ( .A1(n2544), .A2(n2545), .A3(n2546), .A4(n2547), .ZN(n730)
         );
  NOR4_X1 U4170 ( .A1(n2548), .A2(n2549), .A3(n2550), .A4(n2551), .ZN(n2547)
         );
  NAND3_X1 U4171 ( .A1(n6244), .A2(n6243), .A3(n6245), .ZN(n2551) );
  OAI211_X1 U4172 ( .C1(n5560), .C2(n5386), .A(n6241), .B(n6242), .ZN(n2550)
         );
  OAI222_X1 U4173 ( .A1(n5558), .A2(n5258), .B1(n5559), .B2(n5226), .C1(n5561), 
        .C2(n5354), .ZN(n2549) );
  OAI221_X1 U4174 ( .B1(n5531), .B2(n5162), .C1(n5532), .C2(n5194), .A(n2552), 
        .ZN(n2548) );
  AOI22_X1 U4175 ( .A1(n1804), .A2(n1925), .B1(n1805), .B2(n1926), .ZN(n2552)
         );
  INV_X1 U4176 ( .A(n4970), .ZN(n1805) );
  INV_X1 U4177 ( .A(n4938), .ZN(n1804) );
  AOI211_X1 U4178 ( .C1(n1806), .C2(n1927), .A(n2553), .B(n2554), .ZN(n2546)
         );
  OAI22_X1 U4179 ( .A1(n5541), .A2(n4810), .B1(n5551), .B2(n4714), .ZN(n2554)
         );
  OAI222_X1 U4180 ( .A1(n5546), .A2(n4650), .B1(n5552), .B2(n4618), .C1(n5547), 
        .C2(n4682), .ZN(n2553) );
  INV_X1 U4181 ( .A(n4842), .ZN(n1806) );
  AOI221_X1 U4182 ( .B1(n1930), .B2(n1810), .C1(n1931), .C2(n2555), .A(n2556), 
        .ZN(n2545) );
  OAI22_X1 U4183 ( .A1(n4458), .A2(n1934), .B1(n5066), .B2(n1935), .ZN(n2556)
         );
  INV_X1 U4184 ( .A(n5290), .ZN(n2555) );
  INV_X1 U4185 ( .A(n5322), .ZN(n1810) );
  AOI222_X1 U4186 ( .A1(n1812), .A2(n1936), .B1(n1937), .B2(n1813), .C1(n1814), 
        .C2(n1938), .ZN(n2544) );
  INV_X1 U4187 ( .A(n4490), .ZN(n1814) );
  INV_X1 U4188 ( .A(n4426), .ZN(n1813) );
  INV_X1 U4189 ( .A(n4522), .ZN(n1812) );
  AOI22_X1 U4193 ( .A1(n908), .A2(\UUT/break_code[3] ), .B1(n906), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [3]), .ZN(n2558) );
  INV_X1 U4195 ( .A(n2561), .ZN(n2559) );
  INV_X1 U4196 ( .A(n741), .ZN(\UUT/break_code[3] ) );
  AOI22_X1 U4197 ( .A1(n6255), .A2(n2328), .B1(n2329), .B2(
        \UUT/Mcontrol/d_sampled_finstr [3]), .ZN(n741) );
  OAI21_X1 U4198 ( .B1(n6246), .B2(n2562), .A(n2563), .ZN(n2329) );
  INV_X1 U4199 ( .A(n6266), .ZN(n2563) );
  AND2_X1 U4200 ( .A1(n6246), .A2(n913), .ZN(n2328) );
  INV_X1 U4201 ( .A(n2562), .ZN(n913) );
  NAND2_X1 U4202 ( .A1(n6030), .A2(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
        .ZN(n2562) );
  INV_X1 U4203 ( .A(n933), .ZN(n6030) );
  NOR2_X1 U4204 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2089 ), .ZN(n933) );
  AND3_X1 U4205 ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(n2564), .A3(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(n908) );
  AOI222_X1 U4207 ( .A1(n6195), .A2(n5564), .B1(n761), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[3] ), .C2(n5612), .ZN(n5450) );
  NAND2_X1 U4208 ( .A1(n2566), .A2(n2567), .ZN(n761) );
  AOI222_X1 U4209 ( .A1(\UUT/Mpath/the_shift/sh_ror [3]), .A2(n6378), .B1(
        \UUT/Mpath/the_shift/sh_srl [3]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .C1(\UUT/Mpath/the_shift/sh_rol [3]), .C2(n6199), .ZN(n2567) );
  AOI22_X1 U4210 ( .A1(\UUT/Mpath/the_shift/sh_sll [3]), .A2(n6200), .B1(
        \UUT/Mpath/the_shift/sh_sra [3]), .B2(n6198), .ZN(n2566) );
  NAND3_X1 U4211 ( .A1(n2568), .A2(n2569), .A3(n2570), .ZN(n6195) );
  AOI222_X1 U4212 ( .A1(n1208), .A2(n2571), .B1(\UUT/Mpath/the_alu/diff[3] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[3] ), .C2(n1211), .ZN(n2570) );
  INV_X1 U4214 ( .A(n2047), .ZN(n2572) );
  INV_X1 U4215 ( .A(\UUT/Mpath/the_alu/N77 ), .ZN(n2571) );
  INV_X1 U4217 ( .A(n2574), .ZN(n2573) );
  AOI22_X1 U4218 ( .A1(\UUT/Mpath/the_alu/N154 ), .A2(n1212), .B1(
        \UUT/Mpath/the_alu/N122 ), .B2(n1213), .ZN(n2569) );
  INV_X1 U4220 ( .A(\UUT/Mpath/the_alu/N491 ), .ZN(\UUT/Mpath/the_alu/N492 )
         );
  NOR4_X1 U4221 ( .A1(n2047), .A2(n1211), .A3(n2050), .A4(
        \UUT/Mpath/the_alu/N498 ), .ZN(n6348) );
  INV_X1 U4222 ( .A(\UUT/Mpath/the_alu/N503 ), .ZN(n2050) );
  INV_X1 U4224 ( .A(\UUT/Mpath/the_alu/N468 ), .ZN(n2575) );
  NAND2_X1 U4225 ( .A1(\UUT/Mpath/the_alu/N515 ), .A2(\UUT/Mpath/the_alu/N509 ), .ZN(n2047) );
  INV_X1 U4227 ( .A(\UUT/Mpath/the_alu/N486 ), .ZN(n2576) );
  AOI22_X1 U4228 ( .A1(\UUT/Mpath/the_alu/N186 ), .A2(n6365), .B1(
        \UUT/Mpath/the_alu/N218 ), .B2(n1215), .ZN(n2568) );
  NOR3_X1 U4230 ( .A1(\UUT/Mpath/the_alu/N486 ), .A2(n6349), .A3(
        \UUT/Mpath/the_alu/N480 ), .ZN(n2574) );
  INV_X1 U4232 ( .A(\UUT/Mpath/the_alu/N480 ), .ZN(n2577) );
  INV_X1 U4234 ( .A(n753), .ZN(n2565) );
  NAND4_X1 U4235 ( .A1(n2578), .A2(n2579), .A3(n2580), .A4(n2581), .ZN(n753)
         );
  NOR4_X1 U4236 ( .A1(n2582), .A2(n2583), .A3(n2584), .A4(n2585), .ZN(n2581)
         );
  NAND3_X1 U4237 ( .A1(n6253), .A2(n6252), .A3(n6254), .ZN(n2585) );
  OAI211_X1 U4238 ( .C1(n5560), .C2(n5387), .A(n6250), .B(n6251), .ZN(n2584)
         );
  OAI222_X1 U4239 ( .A1(n5558), .A2(n5259), .B1(n5559), .B2(n5227), .C1(n5561), 
        .C2(n5355), .ZN(n2583) );
  OAI221_X1 U4240 ( .B1(n5531), .B2(n5163), .C1(n5532), .C2(n5195), .A(n2586), 
        .ZN(n2582) );
  AOI22_X1 U4241 ( .A1(n1784), .A2(n1925), .B1(n1785), .B2(n1926), .ZN(n2586)
         );
  INV_X1 U4243 ( .A(n4971), .ZN(n1785) );
  INV_X1 U4245 ( .A(n4939), .ZN(n1784) );
  AOI211_X1 U4246 ( .C1(n1786), .C2(n1927), .A(n2587), .B(n2588), .ZN(n2580)
         );
  OAI22_X1 U4247 ( .A1(n5541), .A2(n4811), .B1(n5551), .B2(n4715), .ZN(n2588)
         );
  OAI222_X1 U4248 ( .A1(n5546), .A2(n4651), .B1(n5552), .B2(n4619), .C1(n5547), 
        .C2(n4683), .ZN(n2587) );
  INV_X1 U4250 ( .A(n4843), .ZN(n1786) );
  AOI221_X1 U4251 ( .B1(n1930), .B2(n1790), .C1(n1931), .C2(n2589), .A(n2590), 
        .ZN(n2579) );
  OAI22_X1 U4252 ( .A1(n4459), .A2(n1934), .B1(n5067), .B2(n1935), .ZN(n2590)
         );
  NAND3_X1 U4253 ( .A1(n6306), .A2(n6304), .A3(n6317), .ZN(n1935) );
  INV_X1 U4255 ( .A(n5291), .ZN(n2589) );
  INV_X1 U4257 ( .A(n5323), .ZN(n1790) );
  INV_X1 U4259 ( .A(n6318), .ZN(n2591) );
  AOI222_X1 U4260 ( .A1(n1792), .A2(n1936), .B1(n1937), .B2(n1793), .C1(n1794), 
        .C2(n1938), .ZN(n2578) );
  INV_X1 U4262 ( .A(n4491), .ZN(n1794) );
  INV_X1 U4263 ( .A(n4427), .ZN(n1793) );
  INV_X1 U4266 ( .A(n4523), .ZN(n1792) );
  INV_X1 U4268 ( .A(\UUT/byp_controlA[2] ), .ZN(n2593) );
  INV_X1 U4269 ( .A(n6303), .ZN(n2592) );
  INV_X1 U4271 ( .A(\UUT/Mcontrol/st_logic/N47 ), .ZN(\UUT/byp_controlA[0] )
         );
  NAND2_X1 U4272 ( .A1(\UUT/Mcontrol/bp_logicA/memory_main ), .A2(n2594), .ZN(
        \UUT/Mcontrol/st_logic/N47 ) );
  INV_X1 U4273 ( .A(\UUT/Mcontrol/bp_logicA/exec_main ), .ZN(n2594) );
  AOI21_X1 U4276 ( .B1(n2564), .B2(\UUT/Mcontrol/st_logic/N65 ), .A(n2325), 
        .ZN(n2561) );
  INV_X1 U4277 ( .A(\UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(n2325) );
  INV_X1 U4278 ( .A(\UUT/Mcontrol/Nextpc_decoding/N116 ), .ZN(n2564) );
  INV_X1 U4279 ( .A(\UUT/Mcontrol/st_logic/N103 ), .ZN(n2560) );
  INV_X1 U4280 ( .A(\UUT/Mcontrol/Operation_decoding32/N2084 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2085 ) );
  NOR2_X1 U4281 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2077 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2079 ) );
  INV_X1 U4282 ( .A(\UUT/Mcontrol/Operation_decoding32/N2060 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2061 ) );
  NOR2_X1 U4283 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2041 ), .A2(
        \UUT/Mcontrol/d_instr [26]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2043 ) );
  NOR2_X1 U4284 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2023 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2025 ) );
  NOR2_X1 U4285 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2017 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2019 ) );
  NOR2_X1 U4286 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2005 ), .A2(
        \UUT/Mcontrol/d_instr [26]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2007 ) );
  NOR2_X1 U4287 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1999 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2001 ) );
  INV_X1 U4288 ( .A(\UUT/Mcontrol/Operation_decoding32/N1994 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1995 ) );
  INV_X1 U4289 ( .A(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1976 ) );
  INV_X1 U4290 ( .A(\UUT/Mcontrol/d_instr [26]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1922 ) );
  INV_X1 U4300 ( .A(\localbus/N338 ), .ZN(n4339) );
  INV_X1 U4303 ( .A(\localbus/N62 ), .ZN(n4340) );
  NOR2_X1 U4304 ( .A1(\localbus/c1_op[OP][0] ), .A2(n4343), .ZN(
        \localbus/c1_op[OP][1] ) );
  INV_X1 U4305 ( .A(\localbus/N46 ), .ZN(n4343) );
  NOR2_X1 U4306 ( .A1(\localbus/c1_op[OP][0] ), .A2(\localbus/N46 ), .ZN(
        \localbus/c1_op[MASTER] ) );
  INV_X1 U4315 ( .A(n4352), .ZN(\localbus/c1_addr_outbus[30] ) );
  INV_X1 U4317 ( .A(n4354), .ZN(\localbus/c1_addr_outbus[29] ) );
  INV_X1 U4318 ( .A(n4355), .ZN(\localbus/c1_addr_outbus[28] ) );
  INV_X1 U4319 ( .A(n4356), .ZN(\localbus/c1_addr_outbus[27] ) );
  INV_X1 U4320 ( .A(n4357), .ZN(\localbus/c1_addr_outbus[26] ) );
  INV_X1 U4321 ( .A(n4358), .ZN(\localbus/c1_addr_outbus[25] ) );
  INV_X1 U4322 ( .A(n4359), .ZN(\localbus/c1_addr_outbus[24] ) );
  INV_X1 U4323 ( .A(n4360), .ZN(\localbus/c1_addr_outbus[23] ) );
  INV_X1 U4324 ( .A(n4361), .ZN(\localbus/c1_addr_outbus[22] ) );
  INV_X1 U4325 ( .A(n4362), .ZN(\localbus/c1_addr_outbus[21] ) );
  INV_X1 U4326 ( .A(n4363), .ZN(\localbus/c1_addr_outbus[20] ) );
  INV_X1 U4328 ( .A(n4365), .ZN(\localbus/c1_addr_outbus[19] ) );
  INV_X1 U4329 ( .A(n4366), .ZN(\localbus/c1_addr_outbus[18] ) );
  INV_X1 U4330 ( .A(n4367), .ZN(\localbus/c1_addr_outbus[17] ) );
  INV_X1 U4331 ( .A(n4368), .ZN(\localbus/c1_addr_outbus[16] ) );
  INV_X1 U4332 ( .A(n4369), .ZN(\localbus/c1_addr_outbus[15] ) );
  INV_X1 U4333 ( .A(n4370), .ZN(\localbus/c1_addr_outbus[14] ) );
  INV_X1 U4334 ( .A(n4371), .ZN(\localbus/c1_addr_outbus[13] ) );
  INV_X1 U4339 ( .A(\localbus/N89 ), .ZN(dram_mw) );
  INV_X1 U4340 ( .A(\localbus/N85 ), .ZN(dram_mr) );
  NOR2_X1 U4341 ( .A1(n4376), .A2(n4377), .ZN(dram_data_outbus[9]) );
  NOR2_X1 U4342 ( .A1(n4378), .A2(n4377), .ZN(dram_data_outbus[8]) );
  NOR2_X1 U4343 ( .A1(n4379), .A2(n4380), .ZN(dram_data_outbus[7]) );
  NOR2_X1 U4344 ( .A1(n4379), .A2(n4381), .ZN(dram_data_outbus[6]) );
  NOR2_X1 U4345 ( .A1(n4379), .A2(n4382), .ZN(dram_data_outbus[5]) );
  NOR2_X1 U4346 ( .A1(n4379), .A2(n4383), .ZN(dram_data_outbus[4]) );
  NOR2_X1 U4347 ( .A1(n4379), .A2(n4384), .ZN(dram_data_outbus[3]) );
  NOR2_X1 U4348 ( .A1(n4385), .A2(n4377), .ZN(dram_data_outbus[31]) );
  NOR2_X1 U4349 ( .A1(n4386), .A2(n4377), .ZN(dram_data_outbus[30]) );
  NOR2_X1 U4350 ( .A1(n4379), .A2(n4387), .ZN(dram_data_outbus[2]) );
  NOR2_X1 U4351 ( .A1(n4388), .A2(n4377), .ZN(dram_data_outbus[29]) );
  NOR2_X1 U4352 ( .A1(n4389), .A2(n4377), .ZN(dram_data_outbus[28]) );
  NOR2_X1 U4353 ( .A1(n4390), .A2(n4377), .ZN(dram_data_outbus[27]) );
  NOR2_X1 U4354 ( .A1(n4391), .A2(n4377), .ZN(dram_data_outbus[26]) );
  NOR2_X1 U4355 ( .A1(n4392), .A2(n4377), .ZN(dram_data_outbus[25]) );
  NOR2_X1 U4356 ( .A1(n4393), .A2(n4377), .ZN(dram_data_outbus[24]) );
  NOR2_X1 U4357 ( .A1(n4394), .A2(n4377), .ZN(dram_data_outbus[23]) );
  NOR2_X1 U4358 ( .A1(n4395), .A2(n4377), .ZN(dram_data_outbus[22]) );
  NOR2_X1 U4359 ( .A1(n4396), .A2(n4377), .ZN(dram_data_outbus[21]) );
  NOR2_X1 U4360 ( .A1(n4397), .A2(n4377), .ZN(dram_data_outbus[20]) );
  NOR2_X1 U4361 ( .A1(n4398), .A2(n4379), .ZN(dram_data_outbus[1]) );
  NOR2_X1 U4362 ( .A1(n4399), .A2(n4377), .ZN(dram_data_outbus[19]) );
  NOR2_X1 U4363 ( .A1(n4400), .A2(n4377), .ZN(dram_data_outbus[18]) );
  NOR2_X1 U4364 ( .A1(n4401), .A2(n4377), .ZN(dram_data_outbus[17]) );
  NOR2_X1 U4365 ( .A1(n4402), .A2(n4377), .ZN(dram_data_outbus[16]) );
  NOR2_X1 U4366 ( .A1(n4403), .A2(n4377), .ZN(dram_data_outbus[15]) );
  NOR2_X1 U4367 ( .A1(n4404), .A2(n4377), .ZN(dram_data_outbus[14]) );
  NOR2_X1 U4368 ( .A1(n4405), .A2(n4377), .ZN(dram_data_outbus[13]) );
  NOR2_X1 U4369 ( .A1(n4406), .A2(n4377), .ZN(dram_data_outbus[12]) );
  NOR2_X1 U4370 ( .A1(n4407), .A2(n4377), .ZN(dram_data_outbus[11]) );
  NOR2_X1 U4371 ( .A1(n4408), .A2(n4377), .ZN(dram_data_outbus[10]) );
  INV_X1 U4372 ( .A(\localbus/N218 ), .ZN(n4377) );
  NOR2_X1 U4373 ( .A1(n4409), .A2(n4379), .ZN(dram_data_outbus[0]) );
  NAND2_X1 U4374 ( .A1(\localbus/N218 ), .A2(\localbus/N51 ), .ZN(n4379) );
  NOR2_X1 U4375 ( .A1(n4344), .A2(n4410), .ZN(dram_addr_outbus[9]) );
  NOR2_X1 U4376 ( .A1(n4410), .A2(n4345), .ZN(dram_addr_outbus[8]) );
  NOR2_X1 U4377 ( .A1(n4410), .A2(n4346), .ZN(dram_addr_outbus[7]) );
  NOR2_X1 U4378 ( .A1(n4410), .A2(n4347), .ZN(dram_addr_outbus[6]) );
  NOR2_X1 U4379 ( .A1(n4410), .A2(n4348), .ZN(dram_addr_outbus[5]) );
  NOR2_X1 U4380 ( .A1(n4410), .A2(n4349), .ZN(dram_addr_outbus[4]) );
  NOR2_X1 U4381 ( .A1(n4410), .A2(n4350), .ZN(dram_addr_outbus[3]) );
  NOR2_X1 U4382 ( .A1(n4410), .A2(n4353), .ZN(dram_addr_outbus[2]) );
  NOR2_X1 U4383 ( .A1(n4410), .A2(n4372), .ZN(dram_addr_outbus[12]) );
  NOR2_X1 U4384 ( .A1(n4410), .A2(n4373), .ZN(dram_addr_outbus[11]) );
  NOR2_X1 U4385 ( .A1(n4410), .A2(n4374), .ZN(dram_addr_outbus[10]) );
  INV_X1 U4386 ( .A(\localbus/N215 ), .ZN(n4410) );
  AND4_X1 U4387 ( .A1(n4411), .A2(n4412), .A3(n4413), .A4(n4414), .ZN(
        d_select[31]) );
  NAND2_X1 U4388 ( .A1(n4415), .A2(n4416), .ZN(n4411) );
  INV_X1 U4389 ( .A(N35), .ZN(n4416) );
  AND3_X1 U4390 ( .A1(n4412), .A2(n4413), .A3(n4417), .ZN(d_select[23]) );
  OAI21_X1 U4391 ( .B1(N35), .B2(n4415), .A(n4414), .ZN(n4417) );
  INV_X1 U4392 ( .A(N31), .ZN(n4414) );
  NOR2_X1 U4393 ( .A1(N43), .A2(N42), .ZN(n4415) );
  INV_X1 U4394 ( .A(N27), .ZN(n4413) );
  INV_X1 U4395 ( .A(N22), .ZN(n4412) );
  OAI21_X1 U4396 ( .B1(N43), .B2(n4418), .A(n4419), .ZN(d_select[9]) );
  INV_X1 U4397 ( .A(N42), .ZN(n4418) );
  NAND2_X1 U4398 ( .A1(n4419), .A2(n4420), .ZN(d_select[7]) );
  INV_X1 U4399 ( .A(N43), .ZN(n4420) );
  NOR4_X1 U4400 ( .A1(N22), .A2(N27), .A3(N31), .A4(N35), .ZN(n4419) );
  OR2_X1 U4401 ( .A1(\UUT/Mcontrol/x_sampled_dmem_command[MW] ), .A2(
        \UUT/x_we ), .ZN(dmem_write) );
  AND2_X1 U4402 ( .A1(\UUT/Mcontrol/m_sampled_xrd[4] ), .A2(n5413), .ZN(
        \UUT/regfile/N358 ) );
  AND2_X1 U4403 ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), .A2(n5413), .ZN(
        \UUT/rd_addr [3]) );
  AND2_X1 U4404 ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), .A2(n5413), .ZN(
        \UUT/rd_addr [2]) );
  AND2_X1 U4405 ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), .A2(n5413), .ZN(
        \UUT/rd_addr [1]) );
  OR2_X1 U4406 ( .A1(\UUT/Mcontrol/bp_logicB/memory_main ), .A2(
        \UUT/Mcontrol/bp_logicB/exec_main ), .ZN(\UUT/byp_controlB[2] ) );
  OR2_X1 U4407 ( .A1(\UUT/Mcontrol/bp_logicA/memory_main ), .A2(
        \UUT/Mcontrol/bp_logicA/exec_main ), .ZN(\UUT/byp_controlA[2] ) );
  OAI222_X1 U4408 ( .A1(n5429), .A2(n5430), .B1(n5431), .B2(n5432), .C1(n5433), 
        .C2(n5434), .ZN(\UUT/branch_regb [9]) );
  OAI222_X1 U4409 ( .A1(n5435), .A2(n5430), .B1(n5436), .B2(n5432), .C1(n5437), 
        .C2(n5434), .ZN(\UUT/branch_regb [8]) );
  OAI222_X1 U4410 ( .A1(n5438), .A2(n5430), .B1(n5439), .B2(n5432), .C1(n5440), 
        .C2(n5434), .ZN(\UUT/branch_regb [7]) );
  OAI222_X1 U4411 ( .A1(n5441), .A2(n5430), .B1(n5442), .B2(n5432), .C1(n5443), 
        .C2(n5434), .ZN(\UUT/branch_regb [6]) );
  OAI222_X1 U4412 ( .A1(n5444), .A2(n5430), .B1(n5445), .B2(n5432), .C1(n5446), 
        .C2(n5434), .ZN(\UUT/branch_regb [5]) );
  OAI222_X1 U4413 ( .A1(n5447), .A2(n5430), .B1(n5448), .B2(n5432), .C1(n5449), 
        .C2(n5434), .ZN(\UUT/branch_regb [4]) );
  OAI222_X1 U4414 ( .A1(n5450), .A2(n5430), .B1(n5451), .B2(n5432), .C1(n5452), 
        .C2(n5434), .ZN(\UUT/branch_regb [3]) );
  OAI222_X1 U4416 ( .A1(n6625), .A2(n5430), .B1(n5457), .B2(n5432), .C1(n5458), 
        .C2(n5434), .ZN(\UUT/branch_regb [30]) );
  OAI222_X1 U4417 ( .A1(n5459), .A2(n5430), .B1(n5460), .B2(n5432), .C1(n5461), 
        .C2(n5434), .ZN(\UUT/branch_regb [2]) );
  OAI222_X1 U4419 ( .A1(n5465), .A2(n5430), .B1(n5466), .B2(n5432), .C1(n5467), 
        .C2(n5434), .ZN(\UUT/branch_regb [28]) );
  OAI222_X1 U4422 ( .A1(n5474), .A2(n5430), .B1(n5475), .B2(n5432), .C1(n5476), 
        .C2(n5434), .ZN(\UUT/branch_regb [25]) );
  OAI222_X1 U4423 ( .A1(n5477), .A2(n5430), .B1(n5478), .B2(n5432), .C1(n5479), 
        .C2(n5434), .ZN(\UUT/branch_regb [24]) );
  OAI222_X1 U4424 ( .A1(n5480), .A2(n5430), .B1(n5481), .B2(n5432), .C1(n5482), 
        .C2(n5434), .ZN(\UUT/branch_regb [23]) );
  OAI222_X1 U4425 ( .A1(n5483), .A2(n5430), .B1(n5484), .B2(n5432), .C1(n5485), 
        .C2(n5434), .ZN(\UUT/branch_regb [22]) );
  OAI222_X1 U4426 ( .A1(n5486), .A2(n5430), .B1(n5487), .B2(n5432), .C1(n5488), 
        .C2(n5434), .ZN(\UUT/branch_regb [21]) );
  OAI222_X1 U4427 ( .A1(n5489), .A2(n5430), .B1(n5490), .B2(n5432), .C1(n5491), 
        .C2(n5434), .ZN(\UUT/branch_regb [20]) );
  OAI222_X1 U4428 ( .A1(n5492), .A2(n5430), .B1(n5493), .B2(n5432), .C1(n5494), 
        .C2(n5434), .ZN(\UUT/branch_regb [1]) );
  OAI222_X1 U4429 ( .A1(n5495), .A2(n5430), .B1(n5496), .B2(n5432), .C1(n5497), 
        .C2(n5434), .ZN(\UUT/branch_regb [19]) );
  OAI222_X1 U4430 ( .A1(n5498), .A2(n5430), .B1(n5499), .B2(n5432), .C1(n5500), 
        .C2(n5434), .ZN(\UUT/branch_regb [18]) );
  OAI222_X1 U4431 ( .A1(n5501), .A2(n5430), .B1(n5502), .B2(n5432), .C1(n5503), 
        .C2(n5434), .ZN(\UUT/branch_regb [17]) );
  OAI222_X1 U4432 ( .A1(n5504), .A2(n5430), .B1(n5505), .B2(n5432), .C1(n5506), 
        .C2(n5434), .ZN(\UUT/branch_regb [16]) );
  OAI222_X1 U4433 ( .A1(n5507), .A2(n5430), .B1(n5508), .B2(n5432), .C1(n5509), 
        .C2(n5434), .ZN(\UUT/branch_regb [15]) );
  OAI222_X1 U4434 ( .A1(n5510), .A2(n5430), .B1(n5511), .B2(n5432), .C1(n5512), 
        .C2(n5434), .ZN(\UUT/branch_regb [14]) );
  OAI222_X1 U4435 ( .A1(n5513), .A2(n5430), .B1(n5514), .B2(n5432), .C1(n5515), 
        .C2(n5434), .ZN(\UUT/branch_regb [13]) );
  OAI222_X1 U4436 ( .A1(n5516), .A2(n5430), .B1(n5517), .B2(n5432), .C1(n5518), 
        .C2(n5434), .ZN(\UUT/branch_regb [12]) );
  OAI222_X1 U4437 ( .A1(n5519), .A2(n5430), .B1(n5520), .B2(n5432), .C1(n5521), 
        .C2(n5434), .ZN(\UUT/branch_regb [11]) );
  OAI222_X1 U4438 ( .A1(n5522), .A2(n5430), .B1(n5523), .B2(n5432), .C1(n5524), 
        .C2(n5434), .ZN(\UUT/branch_regb [10]) );
  OAI222_X1 U4439 ( .A1(n5525), .A2(n5430), .B1(n5526), .B2(n5432), .C1(n5527), 
        .C2(n5434), .ZN(\UUT/branch_regb [0]) );
  AOI22_X1 U4444 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][30] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][30] ), .ZN(n5533) );
  AOI22_X1 U4445 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][30] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][30] ), .ZN(n5538) );
  AOI22_X1 U4446 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][30] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][30] ), .ZN(n5543) );
  AOI22_X1 U4447 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][30] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][30] ), .ZN(n5548) );
  AOI22_X1 U4448 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][30] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][30] ), .ZN(n5555) );
  AOI22_X1 U4451 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][29] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][29] ), .ZN(n5565) );
  AOI22_X1 U4452 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][29] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][29] ), .ZN(n5566) );
  AOI22_X1 U4453 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][29] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][29] ), .ZN(n5567) );
  AOI22_X1 U4454 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][29] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][29] ), .ZN(n5568) );
  AOI22_X1 U4455 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][29] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][29] ), .ZN(n5569) );
  AOI22_X1 U4458 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][28] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][28] ), .ZN(n5572) );
  AOI22_X1 U4459 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][28] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][28] ), .ZN(n5573) );
  AOI22_X1 U4460 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][28] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][28] ), .ZN(n5574) );
  AOI22_X1 U4461 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][28] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][28] ), .ZN(n5575) );
  AOI22_X1 U4462 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][28] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][28] ), .ZN(n5576) );
  AOI22_X1 U4465 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][27] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][27] ), .ZN(n5579) );
  AOI22_X1 U4466 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][27] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][27] ), .ZN(n5580) );
  AOI22_X1 U4467 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][27] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][27] ), .ZN(n5581) );
  AOI22_X1 U4468 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][27] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][27] ), .ZN(n5582) );
  AOI22_X1 U4469 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][27] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][27] ), .ZN(n5583) );
  AOI22_X1 U4472 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][26] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][26] ), .ZN(n5586) );
  AOI22_X1 U4473 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][26] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][26] ), .ZN(n5587) );
  AOI22_X1 U4474 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][26] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][26] ), .ZN(n5588) );
  AOI22_X1 U4475 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][26] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][26] ), .ZN(n5589) );
  AOI22_X1 U4476 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][26] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][26] ), .ZN(n5590) );
  AOI22_X1 U4479 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][25] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][25] ), .ZN(n5593) );
  AOI22_X1 U4480 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][25] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][25] ), .ZN(n5594) );
  AOI22_X1 U4481 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][25] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][25] ), .ZN(n5595) );
  AOI22_X1 U4482 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][25] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][25] ), .ZN(n5596) );
  AOI22_X1 U4483 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][25] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][25] ), .ZN(n5597) );
  AOI22_X1 U4484 ( .A1(n5598), .A2(\UUT/Mpath/N119 ), .B1(n5599), .B2(n5564), 
        .ZN(n5474) );
  AOI22_X1 U4486 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][24] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][24] ), .ZN(n5600) );
  AOI22_X1 U4487 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][24] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][24] ), .ZN(n5601) );
  AOI22_X1 U4488 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][24] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][24] ), .ZN(n5602) );
  AOI22_X1 U4489 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][24] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][24] ), .ZN(n5603) );
  AOI22_X1 U4490 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][24] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][24] ), .ZN(n5604) );
  AOI22_X1 U4491 ( .A1(n5605), .A2(\UUT/Mpath/N119 ), .B1(n5606), .B2(n5564), 
        .ZN(n5477) );
  OAI222_X1 U4492 ( .A1(n5525), .A2(n5528), .B1(n5422), .B2(n5529), .C1(n5527), 
        .C2(n5530), .ZN(\UUT/branch_rega [0]) );
  AOI22_X1 U4493 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][0] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][0] ), .ZN(n5607) );
  AOI22_X1 U4494 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][0] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][0] ), .ZN(n5608) );
  AOI22_X1 U4495 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][0] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][0] ), .ZN(n5609) );
  AOI22_X1 U4496 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][0] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][0] ), .ZN(n5610) );
  AOI22_X1 U4497 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][0] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][0] ), .ZN(n5611) );
  AOI222_X1 U4498 ( .A1(\UUT/daddr_out [0]), .A2(n5564), .B1(
        \UUT/Mpath/out_jar[0] ), .B2(n5612), .C1(n5613), .C2(\UUT/Mpath/N119 ), 
        .ZN(n5525) );
  AOI22_X1 U4499 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][9] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][9] ), .ZN(n5718) );
  AOI22_X1 U4500 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][9] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][9] ), .ZN(n5723) );
  AOI22_X1 U4501 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][9] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][9] ), .ZN(n5728) );
  AOI22_X1 U4502 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][9] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][9] ), .ZN(n5733) );
  AOI22_X1 U4503 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][9] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][9] ), .ZN(n5740) );
  AOI22_X1 U4504 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][8] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][8] ), .ZN(n5749) );
  AOI22_X1 U4505 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][8] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][8] ), .ZN(n5750) );
  AOI22_X1 U4506 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][8] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][8] ), .ZN(n5751) );
  AOI22_X1 U4507 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][8] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][8] ), .ZN(n5752) );
  AOI22_X1 U4508 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][8] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][8] ), .ZN(n5753) );
  OAI22_X1 U4509 ( .A1(n5760), .A2(n5761), .B1(n5762), .B2(n5763), .ZN(n5759)
         );
  AOI22_X1 U4510 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][7] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][7] ), .ZN(n5764) );
  AOI22_X1 U4511 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][7] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][7] ), .ZN(n5765) );
  AOI22_X1 U4512 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][7] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][7] ), .ZN(n5766) );
  AOI22_X1 U4513 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][7] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][7] ), .ZN(n5767) );
  AOI22_X1 U4514 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][7] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][7] ), .ZN(n5768) );
  OAI22_X1 U4515 ( .A1(n5761), .A2(n5772), .B1(n5763), .B2(n5773), .ZN(n5771)
         );
  OAI22_X1 U4516 ( .A1(n5776), .A2(n5777), .B1(n5773), .B2(n5778), .ZN(n5775)
         );
  AOI22_X1 U4517 ( .A1(dram_data_inbus[6]), .A2(n5779), .B1(BUS_DATA_INBUS[6]), 
        .B2(n6377), .ZN(n5773) );
  INV_X1 U4518 ( .A(n5772), .ZN(n5774) );
  AOI22_X1 U4519 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][6] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][6] ), .ZN(n5781) );
  AOI22_X1 U4520 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][6] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][6] ), .ZN(n5782) );
  AOI22_X1 U4521 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][6] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][6] ), .ZN(n5783) );
  AOI22_X1 U4522 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][6] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][6] ), .ZN(n5784) );
  AOI22_X1 U4523 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][6] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][6] ), .ZN(n5785) );
  OAI22_X1 U4524 ( .A1(n5761), .A2(n5789), .B1(n5763), .B2(n5790), .ZN(n5788)
         );
  OAI22_X1 U4525 ( .A1(n5793), .A2(n5777), .B1(n5790), .B2(n5778), .ZN(n5792)
         );
  AOI22_X1 U4526 ( .A1(dram_data_inbus[5]), .A2(n5779), .B1(BUS_DATA_INBUS[5]), 
        .B2(n6377), .ZN(n5790) );
  INV_X1 U4527 ( .A(n5789), .ZN(n5791) );
  AOI22_X1 U4528 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][5] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][5] ), .ZN(n5794) );
  AOI22_X1 U4529 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][5] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][5] ), .ZN(n5795) );
  AOI22_X1 U4530 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][5] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][5] ), .ZN(n5796) );
  AOI22_X1 U4531 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][5] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][5] ), .ZN(n5797) );
  AOI22_X1 U4532 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][5] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][5] ), .ZN(n5798) );
  OAI22_X1 U4533 ( .A1(n5761), .A2(n5802), .B1(n5763), .B2(n5803), .ZN(n5801)
         );
  OAI22_X1 U4534 ( .A1(n5806), .A2(n5777), .B1(n5803), .B2(n5778), .ZN(n5805)
         );
  AOI22_X1 U4535 ( .A1(dram_data_inbus[4]), .A2(n5779), .B1(BUS_DATA_INBUS[4]), 
        .B2(n6377), .ZN(n5803) );
  INV_X1 U4536 ( .A(n5802), .ZN(n5804) );
  AOI22_X1 U4537 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][4] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][4] ), .ZN(n5807) );
  AOI22_X1 U4538 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][4] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][4] ), .ZN(n5808) );
  AOI22_X1 U4539 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][4] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][4] ), .ZN(n5809) );
  AOI22_X1 U4540 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][4] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][4] ), .ZN(n5810) );
  AOI22_X1 U4541 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][4] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][4] ), .ZN(n5811) );
  OAI22_X1 U4542 ( .A1(n5761), .A2(n5815), .B1(n5763), .B2(n5816), .ZN(n5814)
         );
  OAI22_X1 U4543 ( .A1(n5819), .A2(n5777), .B1(n5816), .B2(n5778), .ZN(n5818)
         );
  AOI22_X1 U4544 ( .A1(dram_data_inbus[3]), .A2(n5779), .B1(BUS_DATA_INBUS[3]), 
        .B2(n6377), .ZN(n5816) );
  INV_X1 U4545 ( .A(n5815), .ZN(n5817) );
  AOI22_X1 U4546 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][3] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][3] ), .ZN(n5820) );
  AOI22_X1 U4547 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][3] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][3] ), .ZN(n5821) );
  AOI22_X1 U4548 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][3] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][3] ), .ZN(n5822) );
  AOI22_X1 U4549 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][3] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][3] ), .ZN(n5823) );
  AOI22_X1 U4550 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][3] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][3] ), .ZN(n5824) );
  AOI22_X1 U4551 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][31] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][31] ), .ZN(n5826) );
  AOI22_X1 U4552 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][31] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][31] ), .ZN(n5827) );
  AOI22_X1 U4553 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][31] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][31] ), .ZN(n5828) );
  AOI22_X1 U4554 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][31] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][31] ), .ZN(n5829) );
  AOI22_X1 U4555 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][31] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][31] ), .ZN(n5830) );
  AOI22_X1 U4556 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][30] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][30] ), .ZN(n5833) );
  AOI22_X1 U4557 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][30] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][30] ), .ZN(n5834) );
  AOI22_X1 U4558 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][30] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][30] ), .ZN(n5835) );
  AOI22_X1 U4559 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][30] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][30] ), .ZN(n5836) );
  AOI22_X1 U4560 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][30] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][30] ), .ZN(n5837) );
  OAI22_X1 U4561 ( .A1(n5761), .A2(n5841), .B1(n5763), .B2(n5842), .ZN(n5840)
         );
  OAI22_X1 U4562 ( .A1(n5845), .A2(n5777), .B1(n5842), .B2(n5778), .ZN(n5844)
         );
  AOI22_X1 U4563 ( .A1(dram_data_inbus[2]), .A2(n5779), .B1(BUS_DATA_INBUS[2]), 
        .B2(n6377), .ZN(n5842) );
  INV_X1 U4564 ( .A(n5841), .ZN(n5843) );
  AOI22_X1 U4565 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][2] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][2] ), .ZN(n5846) );
  AOI22_X1 U4566 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][2] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][2] ), .ZN(n5847) );
  AOI22_X1 U4567 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][2] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][2] ), .ZN(n5848) );
  AOI22_X1 U4568 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][2] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][2] ), .ZN(n5849) );
  AOI22_X1 U4569 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][2] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][2] ), .ZN(n5850) );
  AOI22_X1 U4570 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][29] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][29] ), .ZN(n5852) );
  AOI22_X1 U4571 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][29] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][29] ), .ZN(n5853) );
  AOI22_X1 U4572 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][29] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][29] ), .ZN(n5854) );
  AOI22_X1 U4573 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][29] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][29] ), .ZN(n5855) );
  AOI22_X1 U4574 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][29] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][29] ), .ZN(n5856) );
  AOI22_X1 U4575 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][28] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][28] ), .ZN(n5858) );
  AOI22_X1 U4576 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][28] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][28] ), .ZN(n5859) );
  AOI22_X1 U4577 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][28] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][28] ), .ZN(n5860) );
  AOI22_X1 U4578 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][28] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][28] ), .ZN(n5861) );
  AOI22_X1 U4579 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][28] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][28] ), .ZN(n5862) );
  AOI22_X1 U4580 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][27] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][27] ), .ZN(n5864) );
  AOI22_X1 U4581 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][27] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][27] ), .ZN(n5865) );
  AOI22_X1 U4582 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][27] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][27] ), .ZN(n5866) );
  AOI22_X1 U4583 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][27] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][27] ), .ZN(n5867) );
  AOI22_X1 U4584 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][27] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][27] ), .ZN(n5868) );
  NOR2_X1 U4585 ( .A1(n5871), .A2(n5872), .ZN(n5869) );
  AOI22_X1 U4586 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][26] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][26] ), .ZN(n5874) );
  AOI22_X1 U4587 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][26] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][26] ), .ZN(n5875) );
  AOI22_X1 U4588 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][26] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][26] ), .ZN(n5876) );
  AOI22_X1 U4589 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][26] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][26] ), .ZN(n5877) );
  AOI22_X1 U4590 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][26] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][26] ), .ZN(n5878) );
  AOI22_X1 U4591 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][25] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][25] ), .ZN(n5883) );
  AOI22_X1 U4592 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][25] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][25] ), .ZN(n5884) );
  AOI22_X1 U4593 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][25] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][25] ), .ZN(n5885) );
  AOI22_X1 U4594 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][25] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][25] ), .ZN(n5886) );
  AOI22_X1 U4595 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][25] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][25] ), .ZN(n5887) );
  AOI22_X1 U4596 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][24] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][24] ), .ZN(n5891) );
  AOI22_X1 U4597 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][24] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][24] ), .ZN(n5892) );
  AOI22_X1 U4598 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][24] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][24] ), .ZN(n5893) );
  AOI22_X1 U4599 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][24] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][24] ), .ZN(n5894) );
  AOI22_X1 U4600 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][24] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][24] ), .ZN(n5895) );
  AOI22_X1 U4601 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][23] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][23] ), .ZN(n5898) );
  AOI22_X1 U4602 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][23] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][23] ), .ZN(n5899) );
  AOI22_X1 U4603 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][23] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][23] ), .ZN(n5900) );
  AOI22_X1 U4604 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][23] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][23] ), .ZN(n5901) );
  AOI22_X1 U4605 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][23] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][23] ), .ZN(n5902) );
  AOI22_X1 U4606 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][22] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][22] ), .ZN(n5903) );
  AOI22_X1 U4607 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][22] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][22] ), .ZN(n5904) );
  AOI22_X1 U4608 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][22] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][22] ), .ZN(n5905) );
  AOI22_X1 U4609 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][22] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][22] ), .ZN(n5906) );
  AOI22_X1 U4610 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][22] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][22] ), .ZN(n5907) );
  AOI22_X1 U4611 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][21] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][21] ), .ZN(n5908) );
  AOI22_X1 U4612 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][21] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][21] ), .ZN(n5909) );
  AOI22_X1 U4613 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][21] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][21] ), .ZN(n5910) );
  AOI22_X1 U4614 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][21] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][21] ), .ZN(n5911) );
  AOI22_X1 U4615 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][21] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][21] ), .ZN(n5912) );
  AOI22_X1 U4616 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][20] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][20] ), .ZN(n5913) );
  AOI22_X1 U4617 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][20] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][20] ), .ZN(n5914) );
  AOI22_X1 U4618 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][20] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][20] ), .ZN(n5915) );
  AOI22_X1 U4619 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][20] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][20] ), .ZN(n5916) );
  AOI22_X1 U4620 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][20] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][20] ), .ZN(n5917) );
  OAI22_X1 U4621 ( .A1(n5761), .A2(n5919), .B1(n5763), .B2(n5920), .ZN(n5918)
         );
  OAI22_X1 U4623 ( .A1(n5921), .A2(n5777), .B1(n5920), .B2(n5778), .ZN(n5923)
         );
  AOI22_X1 U4624 ( .A1(dram_data_inbus[1]), .A2(n5779), .B1(BUS_DATA_INBUS[1]), 
        .B2(n6377), .ZN(n5920) );
  AOI22_X1 U4625 ( .A1(dram_data_inbus[9]), .A2(n5779), .B1(BUS_DATA_INBUS[9]), 
        .B2(n6377), .ZN(n5921) );
  INV_X1 U4626 ( .A(n5882), .ZN(n5712) );
  INV_X1 U4627 ( .A(n5919), .ZN(n5922) );
  AOI22_X1 U4628 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][1] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][1] ), .ZN(n5924) );
  AOI22_X1 U4629 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][1] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][1] ), .ZN(n5925) );
  AOI22_X1 U4630 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][1] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][1] ), .ZN(n5926) );
  AOI22_X1 U4631 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][1] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][1] ), .ZN(n5927) );
  AOI22_X1 U4632 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][1] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][1] ), .ZN(n5928) );
  AOI22_X1 U4633 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][19] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][19] ), .ZN(n5929) );
  AOI22_X1 U4634 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][19] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][19] ), .ZN(n5930) );
  AOI22_X1 U4635 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][19] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][19] ), .ZN(n5931) );
  AOI22_X1 U4636 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][19] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][19] ), .ZN(n5932) );
  AOI22_X1 U4637 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][19] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][19] ), .ZN(n5933) );
  AOI22_X1 U4638 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][18] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][18] ), .ZN(n5934) );
  AOI22_X1 U4639 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][18] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][18] ), .ZN(n5935) );
  AOI22_X1 U4640 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][18] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][18] ), .ZN(n5936) );
  AOI22_X1 U4641 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][18] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][18] ), .ZN(n5937) );
  AOI22_X1 U4642 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][18] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][18] ), .ZN(n5938) );
  AOI22_X1 U4643 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][17] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][17] ), .ZN(n5939) );
  AOI22_X1 U4644 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][17] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][17] ), .ZN(n5940) );
  AOI22_X1 U4645 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][17] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][17] ), .ZN(n5941) );
  AOI22_X1 U4646 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][17] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][17] ), .ZN(n5942) );
  AOI22_X1 U4647 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][17] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][17] ), .ZN(n5943) );
  NOR3_X1 U4648 ( .A1(n5946), .A2(n5947), .A3(n5948), .ZN(n5945) );
  AOI22_X1 U4649 ( .A1(n5758), .A2(n5949), .B1(\UUT/Mpath/the_memhandle/N239 ), 
        .B2(n5756), .ZN(n5947) );
  INV_X1 U4650 ( .A(\UUT/Mpath/the_memhandle/N86 ), .ZN(n5946) );
  AOI22_X1 U4651 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][16] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][16] ), .ZN(n5952) );
  AOI22_X1 U4652 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][16] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][16] ), .ZN(n5953) );
  AOI22_X1 U4653 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][16] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][16] ), .ZN(n5954) );
  AOI22_X1 U4654 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][16] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][16] ), .ZN(n5955) );
  AOI22_X1 U4655 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][16] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][16] ), .ZN(n5956) );
  INV_X1 U4656 ( .A(n5957), .ZN(n5758) );
  INV_X1 U4657 ( .A(n5825), .ZN(n5756) );
  AOI22_X1 U4658 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][15] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][15] ), .ZN(n5958) );
  AOI22_X1 U4659 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][15] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][15] ), .ZN(n5959) );
  AOI22_X1 U4660 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][15] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][15] ), .ZN(n5960) );
  AOI22_X1 U4661 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][15] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][15] ), .ZN(n5961) );
  AOI22_X1 U4662 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][15] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][15] ), .ZN(n5962) );
  AOI22_X1 U4664 ( .A1(dram_data_inbus[14]), .A2(n5779), .B1(
        BUS_DATA_INBUS[14]), .B2(n6377), .ZN(n5776) );
  INV_X1 U4665 ( .A(n5832), .ZN(n5769) );
  AOI22_X1 U4666 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][14] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][14] ), .ZN(n5963) );
  AOI22_X1 U4667 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][14] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][14] ), .ZN(n5964) );
  AOI22_X1 U4668 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][14] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][14] ), .ZN(n5965) );
  AOI22_X1 U4669 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][14] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][14] ), .ZN(n5966) );
  AOI22_X1 U4670 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][14] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][14] ), .ZN(n5967) );
  AOI22_X1 U4672 ( .A1(dram_data_inbus[13]), .A2(n5779), .B1(
        BUS_DATA_INBUS[13]), .B2(n6377), .ZN(n5793) );
  INV_X1 U4673 ( .A(n5851), .ZN(n5786) );
  AOI22_X1 U4674 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][13] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][13] ), .ZN(n5968) );
  AOI22_X1 U4675 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][13] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][13] ), .ZN(n5969) );
  AOI22_X1 U4676 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][13] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][13] ), .ZN(n5970) );
  AOI22_X1 U4677 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][13] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][13] ), .ZN(n5971) );
  AOI22_X1 U4678 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][13] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][13] ), .ZN(n5972) );
  AOI22_X1 U4680 ( .A1(dram_data_inbus[12]), .A2(n5779), .B1(
        BUS_DATA_INBUS[12]), .B2(n6377), .ZN(n5806) );
  INV_X1 U4681 ( .A(n5857), .ZN(n5799) );
  AOI22_X1 U4682 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][12] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][12] ), .ZN(n5973) );
  AOI22_X1 U4683 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][12] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][12] ), .ZN(n5974) );
  AOI22_X1 U4684 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][12] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][12] ), .ZN(n5975) );
  AOI22_X1 U4685 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][12] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][12] ), .ZN(n5976) );
  AOI22_X1 U4686 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][12] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][12] ), .ZN(n5977) );
  AOI22_X1 U4688 ( .A1(dram_data_inbus[11]), .A2(n5779), .B1(
        BUS_DATA_INBUS[11]), .B2(n6377), .ZN(n5819) );
  INV_X1 U4689 ( .A(n5863), .ZN(n5812) );
  AOI22_X1 U4690 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][11] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][11] ), .ZN(n5978) );
  AOI22_X1 U4691 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][11] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][11] ), .ZN(n5979) );
  AOI22_X1 U4692 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][11] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][11] ), .ZN(n5980) );
  AOI22_X1 U4693 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][11] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][11] ), .ZN(n5981) );
  AOI22_X1 U4694 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][11] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][11] ), .ZN(n5982) );
  INV_X1 U4695 ( .A(n5754), .ZN(n5715) );
  OAI22_X1 U4696 ( .A1(n5825), .A2(n5985), .B1(n5760), .B2(n5986), .ZN(n5984)
         );
  INV_X1 U4697 ( .A(\UUT/Mpath/the_memhandle/N37 ), .ZN(n5986) );
  INV_X1 U4698 ( .A(\UUT/Mpath/the_memhandle/N36 ), .ZN(n5985) );
  OAI22_X1 U4699 ( .A1(n5957), .A2(n5777), .B1(n5762), .B2(n5778), .ZN(n5983)
         );
  AOI22_X1 U4700 ( .A1(dram_data_inbus[7]), .A2(n5779), .B1(BUS_DATA_INBUS[7]), 
        .B2(n6377), .ZN(n5762) );
  AOI22_X1 U4701 ( .A1(dram_data_inbus[15]), .A2(n5779), .B1(
        BUS_DATA_INBUS[15]), .B2(n6377), .ZN(n5957) );
  AOI22_X1 U4703 ( .A1(dram_data_inbus[10]), .A2(n5779), .B1(
        BUS_DATA_INBUS[10]), .B2(n6377), .ZN(n5845) );
  NOR2_X1 U4704 ( .A1(n5948), .A2(n5987), .ZN(n5713) );
  INV_X1 U4705 ( .A(n5873), .ZN(n5838) );
  NOR2_X1 U4706 ( .A1(n5988), .A2(n5948), .ZN(n5711) );
  INV_X1 U4707 ( .A(n5950), .ZN(n5948) );
  NOR2_X1 U4708 ( .A1(\UUT/Mpath/the_memhandle/N34 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5950) );
  AOI22_X1 U4709 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][10] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][10] ), .ZN(n5989) );
  AOI22_X1 U4710 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][10] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][10] ), .ZN(n5990) );
  AOI22_X1 U4711 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][10] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][10] ), .ZN(n5991) );
  AOI22_X1 U4712 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][10] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][10] ), .ZN(n5992) );
  AOI22_X1 U4713 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][10] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][10] ), .ZN(n5993) );
  OAI22_X1 U4714 ( .A1(n5761), .A2(n5944), .B1(n5763), .B2(n5995), .ZN(n5994)
         );
  AOI21_X1 U4715 ( .B1(n5996), .B2(n5988), .A(n5997), .ZN(n5763) );
  AND2_X1 U4716 ( .A1(\UUT/Mpath/the_memhandle/N77 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5997) );
  INV_X1 U4717 ( .A(n5998), .ZN(n5761) );
  OAI22_X1 U4718 ( .A1(n5996), .A2(\UUT/Mpath/the_memhandle/N243 ), .B1(
        \UUT/Mpath/the_memhandle/N72 ), .B2(n5988), .ZN(n5998) );
  INV_X1 U4719 ( .A(n5987), .ZN(n5988) );
  NOR2_X1 U4720 ( .A1(n5949), .A2(n5951), .ZN(n5987) );
  NOR2_X1 U4721 ( .A1(\UUT/Mpath/the_memhandle/N120 ), .A2(
        \UUT/Mpath/the_memhandle/N86 ), .ZN(n5951) );
  INV_X1 U4722 ( .A(\UUT/Mpath/the_memhandle/N239 ), .ZN(n5949) );
  INV_X1 U4723 ( .A(\UUT/Mpath/the_memhandle/N72 ), .ZN(n5996) );
  AND2_X1 U4725 ( .A1(\UUT/Mpath/the_memhandle/N76 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5757) );
  AND2_X1 U4726 ( .A1(\UUT/Mpath/the_memhandle/N74 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5755) );
  OAI22_X1 U4727 ( .A1(n5999), .A2(n5777), .B1(n5995), .B2(n5778), .ZN(n6001)
         );
  INV_X1 U4728 ( .A(\UUT/Mpath/the_memhandle/N39 ), .ZN(n5778) );
  AOI22_X1 U4729 ( .A1(dram_data_inbus[0]), .A2(n5779), .B1(BUS_DATA_INBUS[0]), 
        .B2(n6377), .ZN(n5995) );
  INV_X1 U4730 ( .A(\UUT/Mpath/the_memhandle/N38 ), .ZN(n5777) );
  AOI22_X1 U4731 ( .A1(dram_data_inbus[8]), .A2(n5779), .B1(BUS_DATA_INBUS[8]), 
        .B2(n6377), .ZN(n5999) );
  INV_X1 U4732 ( .A(n5890), .ZN(n5747) );
  INV_X1 U4733 ( .A(n5944), .ZN(n6000) );
  NOR3_X1 U4734 ( .A1(\localbus/N93 ), .A2(\localbus/c2_op[MASTER] ), .A3(
        n6002), .ZN(n5780) );
  INV_X1 U4735 ( .A(\localbus/N95 ), .ZN(n6002) );
  INV_X1 U4737 ( .A(\localbus/N93 ), .ZN(n6003) );
  AOI22_X1 U4738 ( .A1(n5719), .A2(\UUT/regfile/reg_out[19][0] ), .B1(n5720), 
        .B2(\UUT/regfile/reg_out[18][0] ), .ZN(n6004) );
  AND2_X1 U4743 ( .A1(n6009), .A2(n6010), .ZN(n6005) );
  AOI22_X1 U4744 ( .A1(n5724), .A2(\UUT/regfile/reg_out[21][0] ), .B1(n5725), 
        .B2(\UUT/regfile/reg_out[20][0] ), .ZN(n6011) );
  NAND3_X1 U4747 ( .A1(n6006), .A2(\UUT/rs2_addr [2]), .A3(n6009), .ZN(n5722)
         );
  NAND4_X1 U4748 ( .A1(n6009), .A2(\UUT/rs2_addr [1]), .A3(\UUT/rs2_addr [0]), 
        .A4(\UUT/rs2_addr [2]), .ZN(n5721) );
  NOR2_X1 U4749 ( .A1(n6014), .A2(\UUT/rs2_addr [3]), .ZN(n6009) );
  AOI22_X1 U4750 ( .A1(n5729), .A2(\UUT/regfile/reg_out[25][0] ), .B1(n5730), 
        .B2(\UUT/regfile/reg_out[24][0] ), .ZN(n6015) );
  NAND3_X1 U4753 ( .A1(n6006), .A2(\UUT/rs2_addr [4]), .A3(n6018), .ZN(n5727)
         );
  AOI22_X1 U4755 ( .A1(n5734), .A2(\UUT/regfile/reg_out[29][0] ), .B1(n5735), 
        .B2(\UUT/regfile/reg_out[28][0] ), .ZN(n6019) );
  NOR2_X1 U4760 ( .A1(n6014), .A2(n6007), .ZN(n6017) );
  AOI22_X1 U4763 ( .A1(n5741), .A2(\UUT/regfile/reg_out[5][0] ), .B1(n5742), 
        .B2(\UUT/regfile/reg_out[4][0] ), .ZN(n6024) );
  NAND3_X1 U4766 ( .A1(\UUT/rs2_addr [2]), .A2(n6022), .A3(n6023), .ZN(n5739)
         );
  NAND3_X1 U4767 ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/rs2_addr [2]), .A3(n6021), 
        .ZN(n5738) );
  AND2_X1 U4768 ( .A1(n6025), .A2(n6022), .ZN(n6021) );
  NOR2_X1 U4771 ( .A1(n6022), .A2(n6010), .ZN(n6020) );
  AND2_X1 U4772 ( .A1(n6013), .A2(n6007), .ZN(n6012) );
  INV_X1 U4773 ( .A(n6022), .ZN(\UUT/rs2_addr [3]) );
  NOR2_X1 U4774 ( .A1(n6010), .A2(\UUT/rs2_addr [1]), .ZN(n6013) );
  INV_X1 U4775 ( .A(\UUT/rs2_addr [2]), .ZN(n6010) );
  INV_X1 U4777 ( .A(n6008), .ZN(\UUT/rs2_addr [1]) );
  AND2_X1 U4779 ( .A1(n6006), .A2(n6014), .ZN(n6023) );
  NOR2_X1 U4780 ( .A1(n6008), .A2(\UUT/rs2_addr [0]), .ZN(n6006) );
  AND2_X1 U4781 ( .A1(n6018), .A2(n6008), .ZN(n6016) );
  NAND2_X1 U4782 ( .A1(\UUT/Mcontrol/d_sampled_finstr [17]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1873 ), .ZN(n6008) );
  NOR2_X1 U4783 ( .A1(n6022), .A2(\UUT/rs2_addr [2]), .ZN(n6018) );
  NAND2_X1 U4784 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(n6026), 
        .ZN(\UUT/rs2_addr [2]) );
  NAND2_X1 U4785 ( .A1(\UUT/Mcontrol/d_sampled_finstr [19]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1873 ), .ZN(n6022) );
  NOR2_X1 U4786 ( .A1(n6007), .A2(\UUT/rs2_addr [4]), .ZN(n6025) );
  INV_X1 U4787 ( .A(n6014), .ZN(\UUT/rs2_addr [4]) );
  NAND2_X1 U4788 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [20]), .ZN(n6014) );
  INV_X1 U4789 ( .A(\UUT/rs2_addr [0]), .ZN(n6007) );
  NAND2_X1 U4790 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(n6027), 
        .ZN(\UUT/rs2_addr [0]) );
  INV_X1 U4791 ( .A(\UUT/Mcontrol/st_logic/N2 ), .ZN(
        \UUT/Mcontrol/st_logic/load_stall ) );
  INV_X1 U4792 ( .A(\UUT/Mcontrol/st_logic/N8 ), .ZN(
        \UUT/Mcontrol/st_logic/branchmul_stall ) );
  INV_X1 U4793 ( .A(\UUT/Mcontrol/st_logic/N6 ), .ZN(
        \UUT/Mcontrol/st_logic/branchlw_stall ) );
  INV_X1 U4794 ( .A(\UUT/Mcontrol/st_logic/N4 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_regb ) );
  INV_X1 U4795 ( .A(\UUT/Mcontrol/st_logic/N3 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_rega ) );
  INV_X1 U4796 ( .A(\UUT/Mcontrol/st_logic/N5 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_main_mem_result ) );
  INV_X1 U4797 ( .A(\UUT/Mcontrol/st_logic/N7 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_main_exe_result ) );
  INV_X1 U4798 ( .A(\UUT/Mcontrol/st_logic/N10 ), .ZN(\UUT/Mcontrol/N19 ) );
  AOI21_X1 U4799 ( .B1(n6040), .B2(\UUT/Mcontrol/Operation_decoding32/N1952 ), 
        .A(\UUT/Mcontrol/Operation_decoding32/N1964 ), .ZN(n6038) );
  NAND4_X1 U4800 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1907 ), .A2(n6044), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N89 ), .A4(n6045), .ZN(n6041)
         );
  NOR3_X1 U4801 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1958 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1970 ), .A3(n6039), .ZN(n6044) );
  NOR4_X1 U4802 ( .A1(n6052), .A2(n6029), .A3(n6053), .A4(n6054), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N255 ) );
  AOI21_X1 U4803 ( .B1(\UUT/Mcontrol/Operation_decoding32/N1928 ), .B2(n6046), 
        .A(\UUT/Mcontrol/Operation_decoding32/N1946 ), .ZN(n6052) );
  OAI21_X1 U4804 ( .B1(n6055), .B2(n6053), .A(n6056), .ZN(
        \UUT/Mcontrol/d_jump_type[2] ) );
  AOI21_X1 U4805 ( .B1(\UUT/Mcontrol/d_sampled_finstr [18]), .B2(n6057), .A(
        n6058), .ZN(n6055) );
  AOI21_X1 U4806 ( .B1(n6059), .B2(n6060), .A(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .ZN(n6058) );
  OAI21_X1 U4807 ( .B1(n6061), .B2(n6053), .A(n6056), .ZN(
        \UUT/Mcontrol/d_jump_type[1] ) );
  AOI21_X1 U4808 ( .B1(\UUT/Mcontrol/d_sampled_finstr [17]), .B2(n6062), .A(
        n6045), .ZN(n6061) );
  OAI21_X1 U4809 ( .B1(n6063), .B2(n6064), .A(n6056), .ZN(
        \UUT/Mcontrol/d_jump_type[0] ) );
  AOI221_X1 U4810 ( .B1(n6065), .B2(n6060), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .C2(
        \UUT/Mcontrol/d_sampled_finstr [16]), .A(n6066), .ZN(n6063) );
  INV_X1 U4811 ( .A(\UUT/Mcontrol/Operation_decoding32/N1940 ), .ZN(n6060) );
  OAI22_X1 U4812 ( .A1(n6027), .A2(n6067), .B1(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .B2(n6059), .ZN(n6065) );
  NOR2_X1 U4813 ( .A1(n6068), .A2(\UUT/Mcontrol/Operation_decoding32/N1934 ), 
        .ZN(n6059) );
  AOI21_X1 U4814 ( .B1(\UUT/Mcontrol/Operation_decoding32/N62 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N89 ), .A(
        \UUT/Mcontrol/Operation_decoding32/N1928 ), .ZN(n6068) );
  INV_X1 U4821 ( .A(\UUT/Mcontrol/Operation_decoding32/N2061 ), .ZN(n6075) );
  OAI211_X1 U4822 ( .C1(n6076), .C2(n6039), .A(n6051), .B(n6078), .ZN(n6077)
         );
  AOI22_X1 U4823 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][1] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][1] ), .ZN(n6080) );
  AOI22_X1 U4824 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][1] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][1] ), .ZN(n6081) );
  AOI22_X1 U4825 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][1] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][1] ), .ZN(n6082) );
  AOI22_X1 U4826 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][1] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][1] ), .ZN(n6083) );
  AOI22_X1 U4827 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][1] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][1] ), .ZN(n6084) );
  INV_X1 U4828 ( .A(n5427), .ZN(\UUT/Mcontrol/d_instr [1]) );
  AOI22_X1 U4829 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][23] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][23] ), .ZN(n6087) );
  AOI22_X1 U4830 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][23] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][23] ), .ZN(n6088) );
  AOI22_X1 U4831 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][23] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][23] ), .ZN(n6089) );
  AOI22_X1 U4832 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][23] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][23] ), .ZN(n6090) );
  AOI22_X1 U4833 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][23] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][23] ), .ZN(n6091) );
  OAI21_X1 U4834 ( .B1(n6037), .B2(n5872), .A(n5880), .ZN(n6093) );
  INV_X1 U4835 ( .A(n6094), .ZN(\UUT/Mcontrol/d_instr [7]) );
  AOI22_X1 U4836 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][22] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][22] ), .ZN(n6095) );
  AOI22_X1 U4837 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][22] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][22] ), .ZN(n6096) );
  AOI22_X1 U4838 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][22] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][22] ), .ZN(n6097) );
  AOI22_X1 U4839 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][22] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][22] ), .ZN(n6098) );
  AOI22_X1 U4840 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][22] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][22] ), .ZN(n6099) );
  OAI21_X1 U4841 ( .B1(n6029), .B2(n5872), .A(n5880), .ZN(n6101) );
  AOI22_X1 U4842 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][21] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][21] ), .ZN(n6102) );
  AOI22_X1 U4843 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][21] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][21] ), .ZN(n6103) );
  AOI22_X1 U4844 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][21] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][21] ), .ZN(n6104) );
  AOI22_X1 U4845 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][21] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][21] ), .ZN(n6105) );
  AOI22_X1 U4846 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][21] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][21] ), .ZN(n6106) );
  OAI21_X1 U4847 ( .B1(n6031), .B2(n5872), .A(n5880), .ZN(n6108) );
  INV_X1 U4848 ( .A(n5423), .ZN(\UUT/Mcontrol/d_instr [5]) );
  AOI22_X1 U4849 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][20] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][20] ), .ZN(n6109) );
  AOI22_X1 U4850 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][20] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][20] ), .ZN(n6110) );
  AOI22_X1 U4851 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][20] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][20] ), .ZN(n6111) );
  AOI22_X1 U4852 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][20] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][20] ), .ZN(n6112) );
  AOI22_X1 U4853 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][20] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][20] ), .ZN(n6113) );
  OAI21_X1 U4854 ( .B1(n5872), .B2(n6026), .A(n5880), .ZN(n6115) );
  OAI21_X1 U4855 ( .B1(n5831), .B2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A(n6117), .ZN(n5870) );
  AOI22_X1 U4856 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][19] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][19] ), .ZN(n6119) );
  AOI22_X1 U4857 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][19] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][19] ), .ZN(n6120) );
  AOI22_X1 U4858 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][19] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][19] ), .ZN(n6121) );
  AOI22_X1 U4859 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][19] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][19] ), .ZN(n6122) );
  AOI22_X1 U4860 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][19] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][19] ), .ZN(n6123) );
  OAI221_X1 U4861 ( .B1(n6034), .B2(n6118), .C1(n5871), .C2(n6446), .A(n6117), 
        .ZN(n6126) );
  AOI22_X1 U4862 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][18] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][18] ), .ZN(n6129) );
  AOI22_X1 U4863 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][18] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][18] ), .ZN(n6130) );
  AOI22_X1 U4864 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][18] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][18] ), .ZN(n6131) );
  AOI22_X1 U4865 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][18] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][18] ), .ZN(n6132) );
  AOI22_X1 U4866 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][18] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][18] ), .ZN(n6133) );
  OAI221_X1 U4867 ( .B1(n6118), .B2(n6027), .C1(n5879), .C2(n6446), .A(n6117), 
        .ZN(n6135) );
  AND2_X1 U4868 ( .A1(n6136), .A2(n6137), .ZN(n6117) );
  OR3_X1 U4869 ( .A1(n6053), .A2(n6045), .A3(n5831), .ZN(n6137) );
  NAND2_X1 U4870 ( .A1(n6064), .A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n6118) );
  OAI21_X1 U4871 ( .B1(n6073), .B2(n6138), .A(n6139), .ZN(n6086) );
  NAND3_X1 U4872 ( .A1(n6140), .A2(n6141), .A3(n6142), .ZN(n6139) );
  INV_X1 U4873 ( .A(n6128), .ZN(n6141) );
  INV_X1 U4874 ( .A(n6143), .ZN(\UUT/Mcontrol/d_instr [6]) );
  OAI21_X1 U4875 ( .B1(n6144), .B2(n6145), .A(n6146), .ZN(n6085) );
  AOI21_X1 U4876 ( .B1(n6078), .B2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
        .A(n6073), .ZN(n6146) );
  INV_X1 U4877 ( .A(n6142), .ZN(n6145) );
  NOR3_X1 U4878 ( .A1(n6048), .A2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
        .A3(n6073), .ZN(n6142) );
  INV_X1 U4879 ( .A(n6039), .ZN(n6144) );
  NAND2_X1 U4880 ( .A1(n6140), .A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n6039) );
  AND4_X1 U4881 ( .A1(n6043), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N1987 ), .A4(n6042), .ZN(n6140)
         );
  NOR3_X1 U4882 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2001 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2007 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1995 ), .ZN(n6043) );
  INV_X1 U4883 ( .A(n5428), .ZN(\UUT/Mcontrol/d_instr [0]) );
  AOI22_X1 U4884 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][17] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][17] ), .ZN(n6147) );
  AOI22_X1 U4885 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][17] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][17] ), .ZN(n6148) );
  AOI22_X1 U4886 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][17] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][17] ), .ZN(n6149) );
  AOI22_X1 U4887 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][17] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][17] ), .ZN(n6150) );
  AOI22_X1 U4888 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][17] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][17] ), .ZN(n6151) );
  OAI221_X1 U4889 ( .B1(n6446), .B2(n5888), .C1(n6154), .C2(n5831), .A(n6136), 
        .ZN(n6153) );
  INV_X1 U4890 ( .A(n6155), .ZN(n6154) );
  AOI22_X1 U4891 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][16] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][16] ), .ZN(n6156) );
  AOI22_X1 U4892 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][16] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][16] ), .ZN(n6157) );
  AOI22_X1 U4893 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][16] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][16] ), .ZN(n6158) );
  AOI22_X1 U4894 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][16] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][16] ), .ZN(n6159) );
  AOI22_X1 U4895 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][16] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][16] ), .ZN(n6160) );
  OAI221_X1 U4896 ( .B1(n6163), .B2(n6032), .C1(n5896), .C2(n6446), .A(n6136), 
        .ZN(n6162) );
  AOI22_X1 U4897 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][15] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][15] ), .ZN(n6164) );
  AOI22_X1 U4898 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][15] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][15] ), .ZN(n6165) );
  AOI22_X1 U4899 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][15] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][15] ), .ZN(n6166) );
  AOI22_X1 U4900 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][15] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][15] ), .ZN(n6167) );
  AOI22_X1 U4901 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][15] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][15] ), .ZN(n6168) );
  AOI21_X1 U4903 ( .B1(n6125), .B2(n6174), .A(n6127), .ZN(n6173) );
  NOR2_X1 U4904 ( .A1(n5831), .A2(n6125), .ZN(n6127) );
  OAI221_X1 U4905 ( .B1(n6163), .B2(n6033), .C1(n6037), .C2(n6446), .A(n6136), 
        .ZN(n6174) );
  NAND2_X1 U4906 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1976 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [15]), .ZN(n6136) );
  AOI22_X1 U4907 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][14] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][14] ), .ZN(n6175) );
  AOI22_X1 U4908 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][14] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][14] ), .ZN(n6176) );
  AOI22_X1 U4909 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][14] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][14] ), .ZN(n6177) );
  AOI22_X1 U4910 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][14] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][14] ), .ZN(n6178) );
  AOI22_X1 U4911 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][14] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][14] ), .ZN(n6179) );
  AOI22_X1 U4913 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][13] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][13] ), .ZN(n6182) );
  AOI22_X1 U4914 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][13] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][13] ), .ZN(n6183) );
  AOI22_X1 U4915 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][13] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][13] ), .ZN(n6184) );
  AOI22_X1 U4916 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][13] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][13] ), .ZN(n6185) );
  AOI22_X1 U4917 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][13] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][13] ), .ZN(n6186) );
  AOI21_X1 U4919 ( .B1(n6207), .B2(\UUT/Mcontrol/Operation_decoding32/N2036 ), 
        .A(\UUT/Mcontrol/Operation_decoding32/N2043 ), .ZN(n6206) );
  OAI21_X1 U4920 ( .B1(n6208), .B2(n6074), .A(
        \UUT/Mcontrol/Operation_decoding32/N2030 ), .ZN(n6207) );
  AOI211_X1 U4921 ( .C1(n6046), .C2(\UUT/Mcontrol/Operation_decoding32/N1945 ), 
        .A(n6066), .B(n6064), .ZN(n6208) );
  INV_X1 U4922 ( .A(n6210), .ZN(n6064) );
  AOI22_X1 U4923 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][9] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][9] ), .ZN(n6211) );
  AOI22_X1 U4924 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][9] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][9] ), .ZN(n6212) );
  AOI22_X1 U4925 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][9] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][9] ), .ZN(n6213) );
  AOI22_X1 U4926 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][9] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][9] ), .ZN(n6214) );
  AOI22_X1 U4927 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][9] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][9] ), .ZN(n6215) );
  OAI222_X1 U4928 ( .A1(n6128), .A2(n5831), .B1(n6163), .B2(n6094), .C1(n5889), 
        .C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(n6216) );
  AOI22_X1 U4929 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][8] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][8] ), .ZN(n6217) );
  AOI22_X1 U4930 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][8] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][8] ), .ZN(n6218) );
  AOI22_X1 U4931 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][8] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][8] ), .ZN(n6219) );
  AOI22_X1 U4932 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][8] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][8] ), .ZN(n6220) );
  AOI22_X1 U4933 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][8] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][8] ), .ZN(n6221) );
  OAI222_X1 U4934 ( .A1(n6128), .A2(n6032), .B1(n6163), .B2(n6143), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n5897), .ZN(n6222) );
  AOI22_X1 U4935 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][7] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][7] ), .ZN(n6223) );
  AOI22_X1 U4936 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][7] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][7] ), .ZN(n6224) );
  AOI22_X1 U4937 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][7] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][7] ), .ZN(n6225) );
  AOI22_X1 U4938 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][7] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][7] ), .ZN(n6226) );
  AOI22_X1 U4939 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][7] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][7] ), .ZN(n6227) );
  OAI222_X1 U4940 ( .A1(n6128), .A2(n6033), .B1(n5423), .B2(n6163), .C1(n6094), 
        .C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(n6228) );
  AOI22_X1 U4941 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][6] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][6] ), .ZN(n6229) );
  AOI22_X1 U4942 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][6] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][6] ), .ZN(n6230) );
  AOI22_X1 U4943 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][6] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][6] ), .ZN(n6231) );
  AOI22_X1 U4944 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][6] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][6] ), .ZN(n6232) );
  AOI22_X1 U4945 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][6] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][6] ), .ZN(n6233) );
  OAI222_X1 U4946 ( .A1(n6128), .A2(n6035), .B1(n5424), .B2(n6163), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n6143), .ZN(n6234) );
  AOI22_X1 U4947 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][5] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][5] ), .ZN(n6235) );
  AOI22_X1 U4948 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][5] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][5] ), .ZN(n6236) );
  AOI22_X1 U4949 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][5] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][5] ), .ZN(n6237) );
  AOI22_X1 U4950 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][5] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][5] ), .ZN(n6238) );
  AOI22_X1 U4951 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][5] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][5] ), .ZN(n6239) );
  OAI222_X1 U4952 ( .A1(n6128), .A2(n6036), .B1(n6163), .B2(n5425), .C1(n5423), 
        .C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(n6240) );
  AOI22_X1 U4953 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][4] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][4] ), .ZN(n6241) );
  AOI22_X1 U4954 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][4] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][4] ), .ZN(n6242) );
  AOI22_X1 U4955 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][4] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][4] ), .ZN(n6243) );
  AOI22_X1 U4956 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][4] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][4] ), .ZN(n6244) );
  AOI22_X1 U4957 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][4] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][4] ), .ZN(n6245) );
  OAI22_X1 U4958 ( .A1(n5881), .A2(n6138), .B1(n6248), .B2(n6048), .ZN(n6247)
         );
  AOI22_X1 U4959 ( .A1(n6125), .A2(n6249), .B1(\UUT/Mcontrol/d_instr [4]), 
        .B2(n6209), .ZN(n6248) );
  INV_X1 U4960 ( .A(n5424), .ZN(\UUT/Mcontrol/d_instr [4]) );
  OAI222_X1 U4961 ( .A1(n6128), .A2(n5881), .B1(n6163), .B2(n5426), .C1(n5424), 
        .C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(n6249) );
  AOI22_X1 U4962 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][3] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][3] ), .ZN(n6250) );
  AOI22_X1 U4963 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][3] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][3] ), .ZN(n6251) );
  AOI22_X1 U4964 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][3] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][3] ), .ZN(n6252) );
  AOI22_X1 U4965 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][3] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][3] ), .ZN(n6253) );
  AOI22_X1 U4966 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][3] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][3] ), .ZN(n6254) );
  OAI22_X1 U4967 ( .A1(n5889), .A2(n6138), .B1(n6256), .B2(n6048), .ZN(n6255)
         );
  AOI22_X1 U4968 ( .A1(n6125), .A2(n6257), .B1(\UUT/Mcontrol/d_instr [3]), 
        .B2(n6209), .ZN(n6256) );
  INV_X1 U4969 ( .A(n5425), .ZN(\UUT/Mcontrol/d_instr [3]) );
  OAI222_X1 U4970 ( .A1(n6128), .A2(n5889), .B1(n6163), .B2(n5427), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n5425), .ZN(n6257) );
  AOI22_X1 U4971 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][2] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][2] ), .ZN(n6258) );
  AOI22_X1 U4972 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][2] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][2] ), .ZN(n6259) );
  AOI22_X1 U4973 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][2] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][2] ), .ZN(n6260) );
  AOI22_X1 U4974 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][2] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][2] ), .ZN(n6261) );
  AOI22_X1 U4975 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][2] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][2] ), .ZN(n6262) );
  OAI22_X1 U4976 ( .A1(n5897), .A2(n6138), .B1(n6264), .B2(n6048), .ZN(n6263)
         );
  AOI22_X1 U4977 ( .A1(n6125), .A2(n6265), .B1(\UUT/Mcontrol/d_instr [2]), 
        .B2(n6209), .ZN(n6264) );
  INV_X1 U4978 ( .A(n5426), .ZN(\UUT/Mcontrol/d_instr [2]) );
  OAI222_X1 U4979 ( .A1(n6128), .A2(n5897), .B1(n6163), .B2(n5428), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n5426), .ZN(n6265) );
  NAND2_X1 U4980 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2037 ), .A2(n6028), 
        .ZN(n6138) );
  AND2_X1 U4981 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2085 ), .A2(n6030), 
        .ZN(n6266) );
  NOR2_X1 U4982 ( .A1(n6073), .A2(\UUT/Mcontrol/Operation_decoding32/N2079 ), 
        .ZN(n6246) );
  AOI22_X1 U4983 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][12] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][12] ), .ZN(n6267) );
  AOI22_X1 U4984 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][12] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][12] ), .ZN(n6268) );
  AOI22_X1 U4985 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][12] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][12] ), .ZN(n6269) );
  AOI22_X1 U4986 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][12] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][12] ), .ZN(n6270) );
  AOI22_X1 U4987 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][12] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][12] ), .ZN(n6271) );
  AOI22_X1 U4989 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][11] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][11] ), .ZN(n6273) );
  AOI22_X1 U4990 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][11] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][11] ), .ZN(n6274) );
  AOI22_X1 U4991 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][11] ), .B1(n6367), 
        .B2(\UUT/regfile/reg_out[24][11] ), .ZN(n6275) );
  AOI22_X1 U4992 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][11] ), .B1(n6370), 
        .B2(\UUT/regfile/reg_out[28][11] ), .ZN(n6276) );
  AOI22_X1 U4993 ( .A1(n6375), .A2(\UUT/regfile/reg_out[5][11] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][11] ), .ZN(n6277) );
  AOI22_X1 U4995 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][10] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][10] ), .ZN(n6279) );
  AOI22_X1 U4996 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][10] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][10] ), .ZN(n6280) );
  AOI22_X1 U4997 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][10] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][10] ), .ZN(n6281) );
  AOI22_X1 U4998 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][10] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][10] ), .ZN(n6282) );
  AOI22_X1 U4999 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][10] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][10] ), .ZN(n6283) );
  INV_X1 U5001 ( .A(\UUT/Mpath/N115 ), .ZN(n6284) );
  NAND3_X1 U5002 ( .A1(n6056), .A2(n6285), .A3(n6286), .ZN(
        \UUT/Mcontrol/d_jump_type[3] ) );
  AOI21_X1 U5003 ( .B1(\UUT/Mcontrol/d_sampled_finstr [19]), .B2(n6062), .A(
        n6045), .ZN(n6286) );
  NAND2_X1 U5004 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1945 ), .A2(n6079), 
        .ZN(n6062) );
  INV_X1 U5005 ( .A(n6054), .ZN(n6056) );
  NAND3_X1 U5006 ( .A1(n6125), .A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
        .A3(n6050), .ZN(n6054) );
  NOR2_X1 U5009 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N25 ), .A2(n6290), .ZN(
        n6291) );
  INV_X1 U5010 ( .A(\UUT/Mcontrol/Nextpc_decoding/N260 ), .ZN(n6290) );
  AOI21_X1 U5012 ( .B1(n6295), .B2(n6294), .A(n6296), .ZN(n6293) );
  INV_X1 U5014 ( .A(\UUT/Mcontrol/Nextpc_decoding/N248 ), .ZN(n6295) );
  INV_X1 U5018 ( .A(\UUT/Mcontrol/Nextpc_decoding/N242 ), .ZN(n6297) );
  AOI22_X1 U5020 ( .A1(n5534), .A2(\UUT/regfile/reg_out[19][31] ), .B1(n5535), 
        .B2(\UUT/regfile/reg_out[18][31] ), .ZN(n6300) );
  AND2_X1 U5025 ( .A1(n6305), .A2(n6306), .ZN(n6301) );
  AOI22_X1 U5026 ( .A1(n5539), .A2(\UUT/regfile/reg_out[21][31] ), .B1(n5540), 
        .B2(\UUT/regfile/reg_out[20][31] ), .ZN(n6307) );
  NAND3_X1 U5029 ( .A1(n6302), .A2(\UUT/rs1_addr [2]), .A3(n6305), .ZN(n5537)
         );
  NAND4_X1 U5030 ( .A1(n6305), .A2(\UUT/rs1_addr [1]), .A3(\UUT/rs1_addr [0]), 
        .A4(\UUT/rs1_addr [2]), .ZN(n5536) );
  NOR2_X1 U5031 ( .A1(n6310), .A2(\UUT/rs1_addr [3]), .ZN(n6305) );
  AOI22_X1 U5032 ( .A1(n5544), .A2(\UUT/regfile/reg_out[25][31] ), .B1(n6368), 
        .B2(\UUT/regfile/reg_out[24][31] ), .ZN(n6311) );
  AND3_X1 U5033 ( .A1(\UUT/rs1_addr [4]), .A2(n6303), .A3(n6312), .ZN(n5545)
         );
  NAND3_X1 U5035 ( .A1(n6302), .A2(\UUT/rs1_addr [4]), .A3(n6314), .ZN(n5542)
         );
  AOI22_X1 U5037 ( .A1(n5549), .A2(\UUT/regfile/reg_out[29][31] ), .B1(n6371), 
        .B2(\UUT/regfile/reg_out[28][31] ), .ZN(n6315) );
  NOR2_X1 U5042 ( .A1(n6310), .A2(n6303), .ZN(n6313) );
  AOI22_X1 U5045 ( .A1(n6376), .A2(\UUT/regfile/reg_out[5][31] ), .B1(n5557), 
        .B2(\UUT/regfile/reg_out[4][31] ), .ZN(n6320) );
  NAND3_X1 U5048 ( .A1(\UUT/rs1_addr [2]), .A2(n6318), .A3(n6319), .ZN(n5554)
         );
  NAND3_X1 U5049 ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/rs1_addr [2]), .A3(n6317), 
        .ZN(n5553) );
  AND2_X1 U5050 ( .A1(n6321), .A2(n6318), .ZN(n6317) );
  NOR2_X1 U5053 ( .A1(n6318), .A2(n6306), .ZN(n6316) );
  NOR2_X1 U5055 ( .A1(n6306), .A2(\UUT/rs1_addr [1]), .ZN(n6309) );
  AND2_X1 U5059 ( .A1(n6302), .A2(n6310), .ZN(n6319) );
  INV_X1 U5061 ( .A(\UUT/rs1_addr [4]), .ZN(n6310) );
  AND2_X1 U5062 ( .A1(n6314), .A2(n6304), .ZN(n6312) );
  INV_X1 U5063 ( .A(\UUT/rs1_addr [1]), .ZN(n6304) );
  NOR2_X1 U5065 ( .A1(n6318), .A2(\UUT/rs1_addr [2]), .ZN(n6314) );
  NAND2_X1 U5066 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1871 ), .A2(n5888), 
        .ZN(\UUT/rs1_addr [2]) );
  INV_X1 U5067 ( .A(\UUT/rs1_addr [3]), .ZN(n6318) );
  NOR2_X1 U5068 ( .A1(n5879), .A2(n6322), .ZN(\UUT/rs1_addr [3]) );
  NOR2_X1 U5069 ( .A1(n6303), .A2(\UUT/rs1_addr [4]), .ZN(n6321) );
  NOR2_X1 U5070 ( .A1(n6322), .A2(n5871), .ZN(\UUT/rs1_addr [4]) );
  INV_X1 U5071 ( .A(\UUT/rs1_addr [0]), .ZN(n6303) );
  NOR2_X1 U5072 ( .A1(n6037), .A2(n6322), .ZN(\UUT/rs1_addr [0]) );
  INV_X1 U5073 ( .A(\UUT/Mcontrol/Operation_decoding32/N1871 ), .ZN(n6322) );
  INV_X1 U5077 ( .A(n6324), .ZN(n6323) );
  NOR3_X1 U5079 ( .A1(\UUT/Mpath/the_shift/N115 ), .A2(
        \UUT/Mpath/the_shift/N118 ), .A3(\UUT/Mpath/the_shift/N111 ), .ZN(
        n6324) );
  INV_X1 U5081 ( .A(\UUT/Mpath/the_shift/N115 ), .ZN(n6325) );
  NOR3_X1 U5082 ( .A1(\UUT/Mpath/the_shift/N115 ), .A2(
        \UUT/Mpath/the_shift/N118 ), .A3(n6326), .ZN(n6201) );
  INV_X1 U5083 ( .A(\UUT/Mpath/the_shift/N111 ), .ZN(n6326) );
  INV_X1 U5084 ( .A(\UUT/Mcontrol/Nextpc_decoding/N254 ), .ZN(n6292) );
  INV_X1 U5085 ( .A(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6287) );
  OAI222_X1 U5086 ( .A1(n6128), .A2(n6027), .B1(n6163), .B2(n5897), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n5881), .ZN(n6327) );
  OAI21_X1 U5088 ( .B1(n6045), .B2(n6066), .A(n6210), .ZN(n6155) );
  NAND2_X1 U5089 ( .A1(n6328), .A2(n6040), .ZN(n6066) );
  INV_X1 U5093 ( .A(\UUT/Mcontrol/Operation_decoding32/N1928 ), .ZN(n6067) );
  NOR2_X1 U5096 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1934 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1940 ), .ZN(n6046) );
  INV_X1 U5097 ( .A(n6053), .ZN(n6285) );
  INV_X1 U5100 ( .A(\UUT/Mcontrol/Operation_decoding32/N1958 ), .ZN(n6040) );
  INV_X1 U5101 ( .A(\UUT/Mcontrol/Operation_decoding32/N1952 ), .ZN(n6328) );
  INV_X1 U5102 ( .A(n6209), .ZN(n6125) );
  NAND2_X1 U5103 ( .A1(n6116), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .ZN(n6209) );
  NOR2_X1 U5104 ( .A1(n6048), .A2(n6170), .ZN(n6172) );
  NOR2_X1 U5105 ( .A1(n6587), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .ZN(n6078) );
  INV_X1 U5106 ( .A(\localbus/N90 ), .ZN(BUS_MW) );
  INV_X1 U5107 ( .A(\localbus/N86 ), .ZN(BUS_MR) );
  NOR2_X1 U5108 ( .A1(n4376), .A2(n6329), .ZN(BUS_DATA_OUTBUS[9]) );
  AOI22_X1 U5109 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[9] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[1]), .ZN(n4376) );
  NOR2_X1 U5110 ( .A1(n4378), .A2(n6329), .ZN(BUS_DATA_OUTBUS[8]) );
  AOI22_X1 U5111 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[8] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[0]), .ZN(n4378) );
  NOR2_X1 U5112 ( .A1(n4380), .A2(n6332), .ZN(BUS_DATA_OUTBUS[7]) );
  NOR2_X1 U5113 ( .A1(n4381), .A2(n6332), .ZN(BUS_DATA_OUTBUS[6]) );
  NOR2_X1 U5114 ( .A1(n4382), .A2(n6332), .ZN(BUS_DATA_OUTBUS[5]) );
  NOR2_X1 U5115 ( .A1(n4383), .A2(n6332), .ZN(BUS_DATA_OUTBUS[4]) );
  NOR2_X1 U5116 ( .A1(n4384), .A2(n6332), .ZN(BUS_DATA_OUTBUS[3]) );
  NOR2_X1 U5117 ( .A1(n4385), .A2(n6329), .ZN(BUS_DATA_OUTBUS[31]) );
  AOI221_X1 U5118 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[7]), .A(n6334), .ZN(n4385) );
  AND2_X1 U5119 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[31] ), .A2(n6335), 
        .ZN(n6334) );
  NOR2_X1 U5120 ( .A1(n4386), .A2(n6329), .ZN(BUS_DATA_OUTBUS[30]) );
  AOI221_X1 U5121 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[6]), .A(n6336), .ZN(n4386) );
  AND2_X1 U5122 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[30] ), .A2(n6335), 
        .ZN(n6336) );
  NOR2_X1 U5123 ( .A1(n4387), .A2(n6332), .ZN(BUS_DATA_OUTBUS[2]) );
  NOR2_X1 U5124 ( .A1(n4388), .A2(n6329), .ZN(BUS_DATA_OUTBUS[29]) );
  AOI221_X1 U5125 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[5]), .A(n6337), .ZN(n4388) );
  AND2_X1 U5126 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[29] ), .A2(n6335), 
        .ZN(n6337) );
  NOR2_X1 U5127 ( .A1(n4389), .A2(n6329), .ZN(BUS_DATA_OUTBUS[28]) );
  AOI221_X1 U5128 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[4]), .A(n6338), .ZN(n4389) );
  AND2_X1 U5129 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[28] ), .A2(n6335), 
        .ZN(n6338) );
  NOR2_X1 U5130 ( .A1(n4390), .A2(n6329), .ZN(BUS_DATA_OUTBUS[27]) );
  AOI221_X1 U5131 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[3]), .A(n6339), .ZN(n4390) );
  AND2_X1 U5132 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[27] ), .A2(n6335), 
        .ZN(n6339) );
  NOR2_X1 U5133 ( .A1(n4391), .A2(n6329), .ZN(BUS_DATA_OUTBUS[26]) );
  AOI221_X1 U5134 ( .B1(n6333), .B2(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
        .C1(n6331), .C2(D_DATA_OUTBUS[2]), .A(n6340), .ZN(n4391) );
  AND2_X1 U5135 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[26] ), .A2(n6335), 
        .ZN(n6340) );
  NOR2_X1 U5136 ( .A1(n4392), .A2(n6329), .ZN(BUS_DATA_OUTBUS[25]) );
  AOI221_X1 U5137 ( .B1(\UUT/Mpath/the_memhandle/smdr_out[9] ), .B2(n6333), 
        .C1(n6331), .C2(D_DATA_OUTBUS[1]), .A(n6341), .ZN(n4392) );
  AND2_X1 U5138 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[25] ), .A2(n6335), 
        .ZN(n6341) );
  NOR2_X1 U5139 ( .A1(n4393), .A2(n6329), .ZN(BUS_DATA_OUTBUS[24]) );
  AOI221_X1 U5140 ( .B1(\UUT/Mpath/the_memhandle/smdr_out[8] ), .B2(n6333), 
        .C1(n6331), .C2(D_DATA_OUTBUS[0]), .A(n6342), .ZN(n4393) );
  AND2_X1 U5141 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[24] ), .A2(n6335), 
        .ZN(n6342) );
  INV_X1 U5142 ( .A(n6343), .ZN(n6333) );
  NOR2_X1 U5143 ( .A1(n4394), .A2(n6329), .ZN(BUS_DATA_OUTBUS[23]) );
  AOI22_X1 U5144 ( .A1(n6344), .A2(D_DATA_OUTBUS[7]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[23] ), .ZN(n4394) );
  NOR2_X1 U5145 ( .A1(n4395), .A2(n6329), .ZN(BUS_DATA_OUTBUS[22]) );
  AOI22_X1 U5146 ( .A1(n6344), .A2(D_DATA_OUTBUS[6]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[22] ), .ZN(n4395) );
  NOR2_X1 U5147 ( .A1(n4396), .A2(n6329), .ZN(BUS_DATA_OUTBUS[21]) );
  AOI22_X1 U5148 ( .A1(n6344), .A2(D_DATA_OUTBUS[5]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[21] ), .ZN(n4396) );
  NOR2_X1 U5149 ( .A1(n4397), .A2(n6329), .ZN(BUS_DATA_OUTBUS[20]) );
  AOI22_X1 U5150 ( .A1(n6344), .A2(D_DATA_OUTBUS[4]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[20] ), .ZN(n4397) );
  NOR2_X1 U5151 ( .A1(n4398), .A2(n6332), .ZN(BUS_DATA_OUTBUS[1]) );
  NOR2_X1 U5152 ( .A1(n4399), .A2(n6329), .ZN(BUS_DATA_OUTBUS[19]) );
  AOI22_X1 U5153 ( .A1(n6344), .A2(D_DATA_OUTBUS[3]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[19] ), .ZN(n4399) );
  NOR2_X1 U5154 ( .A1(n4400), .A2(n6329), .ZN(BUS_DATA_OUTBUS[18]) );
  AOI22_X1 U5155 ( .A1(n6344), .A2(D_DATA_OUTBUS[2]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[18] ), .ZN(n4400) );
  NOR2_X1 U5156 ( .A1(n4401), .A2(n6329), .ZN(BUS_DATA_OUTBUS[17]) );
  AOI22_X1 U5157 ( .A1(n6344), .A2(D_DATA_OUTBUS[1]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[17] ), .ZN(n4401) );
  NOR2_X1 U5158 ( .A1(n4402), .A2(n6329), .ZN(BUS_DATA_OUTBUS[16]) );
  AOI22_X1 U5159 ( .A1(n6344), .A2(D_DATA_OUTBUS[0]), .B1(n6335), .B2(
        \UUT/Mpath/the_memhandle/smdr_out[16] ), .ZN(n4402) );
  AND2_X1 U5160 ( .A1(n6330), .A2(dmem_ishalf), .ZN(n6335) );
  NAND2_X1 U5161 ( .A1(n6345), .A2(n6343), .ZN(n6344) );
  NAND2_X1 U5162 ( .A1(\UUT/Mpath/the_memhandle/N237 ), .A2(n6330), .ZN(n6343)
         );
  NOR2_X1 U5163 ( .A1(n4403), .A2(n6329), .ZN(BUS_DATA_OUTBUS[15]) );
  AOI22_X1 U5164 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[7]), .ZN(n4403) );
  NOR2_X1 U5165 ( .A1(n4404), .A2(n6329), .ZN(BUS_DATA_OUTBUS[14]) );
  AOI22_X1 U5166 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[6]), .ZN(n4404) );
  NOR2_X1 U5167 ( .A1(n4405), .A2(n6329), .ZN(BUS_DATA_OUTBUS[13]) );
  AOI22_X1 U5168 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[5]), .ZN(n4405) );
  NOR2_X1 U5169 ( .A1(n4406), .A2(n6329), .ZN(BUS_DATA_OUTBUS[12]) );
  AOI22_X1 U5170 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[4]), .ZN(n4406) );
  NOR2_X1 U5171 ( .A1(n4407), .A2(n6329), .ZN(BUS_DATA_OUTBUS[11]) );
  AOI22_X1 U5172 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[3]), .ZN(n4407) );
  NOR2_X1 U5173 ( .A1(n4408), .A2(n6329), .ZN(BUS_DATA_OUTBUS[10]) );
  INV_X1 U5174 ( .A(\localbus/N229 ), .ZN(n6329) );
  AOI22_X1 U5175 ( .A1(n6330), .A2(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
        .B1(n6331), .B2(D_DATA_OUTBUS[2]), .ZN(n4408) );
  INV_X1 U5176 ( .A(n6345), .ZN(n6331) );
  NAND2_X1 U5177 ( .A1(\localbus/N51 ), .A2(\UUT/Mpath/the_memhandle/N234 ), 
        .ZN(n6345) );
  AND2_X1 U5178 ( .A1(\localbus/N51 ), .A2(dmem_isbyte), .ZN(n6330) );
  NOR2_X1 U5179 ( .A1(n4409), .A2(n6332), .ZN(BUS_DATA_OUTBUS[0]) );
  NAND2_X1 U5180 ( .A1(\localbus/N229 ), .A2(\localbus/N51 ), .ZN(n6332) );
  NOR2_X1 U5181 ( .A1(n4344), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[9]) );
  NAND2_X1 U5182 ( .A1(n6347), .A2(n6189), .ZN(n4344) );
  NOR2_X1 U5183 ( .A1(n4345), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[8]) );
  NAND2_X1 U5184 ( .A1(n6347), .A2(n6190), .ZN(n4345) );
  NOR2_X1 U5185 ( .A1(n4346), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[7]) );
  NAND2_X1 U5186 ( .A1(n6347), .A2(n6191), .ZN(n4346) );
  NOR2_X1 U5187 ( .A1(n4347), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[6]) );
  NAND2_X1 U5188 ( .A1(n6347), .A2(n6192), .ZN(n4347) );
  NOR2_X1 U5189 ( .A1(n4348), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[5]) );
  NAND2_X1 U5190 ( .A1(n6347), .A2(n6193), .ZN(n4348) );
  NOR2_X1 U5191 ( .A1(n4349), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[4]) );
  NAND2_X1 U5192 ( .A1(n6347), .A2(n6194), .ZN(n4349) );
  NOR2_X1 U5193 ( .A1(n4350), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[3]) );
  NAND2_X1 U5194 ( .A1(n6347), .A2(n6195), .ZN(n4350) );
  NOR2_X1 U5195 ( .A1(n6346), .A2(n4351), .ZN(BUS_ADDR_OUTBUS[31]) );
  NOR2_X1 U5197 ( .A1(n6346), .A2(n4352), .ZN(BUS_ADDR_OUTBUS[30]) );
  NAND2_X1 U5198 ( .A1(n6347), .A2(n6542), .ZN(n4352) );
  NOR2_X1 U5199 ( .A1(n4353), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[2]) );
  NAND2_X1 U5200 ( .A1(n6347), .A2(n6202), .ZN(n4353) );
  NOR2_X1 U5201 ( .A1(n6346), .A2(n4354), .ZN(BUS_ADDR_OUTBUS[29]) );
  NAND2_X1 U5202 ( .A1(n6347), .A2(n5571), .ZN(n4354) );
  NOR2_X1 U5203 ( .A1(n6346), .A2(n4355), .ZN(BUS_ADDR_OUTBUS[28]) );
  NAND2_X1 U5204 ( .A1(n6347), .A2(n6452), .ZN(n4355) );
  NOR2_X1 U5205 ( .A1(n6346), .A2(n4356), .ZN(BUS_ADDR_OUTBUS[27]) );
  NAND2_X1 U5206 ( .A1(n6347), .A2(n5585), .ZN(n4356) );
  NOR2_X1 U5207 ( .A1(n6346), .A2(n4357), .ZN(BUS_ADDR_OUTBUS[26]) );
  NAND2_X1 U5208 ( .A1(n6347), .A2(n5592), .ZN(n4357) );
  NOR2_X1 U5209 ( .A1(n6346), .A2(n4358), .ZN(BUS_ADDR_OUTBUS[25]) );
  NAND2_X1 U5210 ( .A1(n6347), .A2(n5599), .ZN(n4358) );
  NOR2_X1 U5211 ( .A1(n6346), .A2(n4359), .ZN(BUS_ADDR_OUTBUS[24]) );
  NAND2_X1 U5212 ( .A1(n6347), .A2(n5606), .ZN(n4359) );
  NOR2_X1 U5213 ( .A1(n6346), .A2(n4360), .ZN(BUS_ADDR_OUTBUS[23]) );
  NAND2_X1 U5214 ( .A1(n6347), .A2(n6092), .ZN(n4360) );
  NOR2_X1 U5215 ( .A1(n6346), .A2(n4361), .ZN(BUS_ADDR_OUTBUS[22]) );
  NAND2_X1 U5216 ( .A1(n6347), .A2(n6100), .ZN(n4361) );
  NOR2_X1 U5217 ( .A1(n6346), .A2(n4362), .ZN(BUS_ADDR_OUTBUS[21]) );
  NAND2_X1 U5218 ( .A1(n6347), .A2(n6107), .ZN(n4362) );
  NOR2_X1 U5219 ( .A1(n6346), .A2(n4363), .ZN(BUS_ADDR_OUTBUS[20]) );
  NAND2_X1 U5220 ( .A1(n6347), .A2(n6114), .ZN(n4363) );
  NOR2_X1 U5221 ( .A1(n6346), .A2(n4364), .ZN(BUS_ADDR_OUTBUS[1]) );
  NAND2_X1 U5222 ( .A1(D_ADDR_OUTBUS[1]), .A2(\localbus/N50 ), .ZN(n4364) );
  AND2_X1 U5223 ( .A1(\UUT/N3 ), .A2(\UUT/daddr_out [1]), .ZN(D_ADDR_OUTBUS[1]) );
  NOR2_X1 U5224 ( .A1(n6346), .A2(n4365), .ZN(BUS_ADDR_OUTBUS[19]) );
  NAND2_X1 U5225 ( .A1(n6347), .A2(n6124), .ZN(n4365) );
  NOR2_X1 U5226 ( .A1(n6346), .A2(n4366), .ZN(BUS_ADDR_OUTBUS[18]) );
  NAND2_X1 U5227 ( .A1(n6347), .A2(n6134), .ZN(n4366) );
  NOR2_X1 U5228 ( .A1(n6346), .A2(n4367), .ZN(BUS_ADDR_OUTBUS[17]) );
  NAND2_X1 U5229 ( .A1(n6347), .A2(n6152), .ZN(n4367) );
  NOR2_X1 U5230 ( .A1(n6346), .A2(n4368), .ZN(BUS_ADDR_OUTBUS[16]) );
  NAND2_X1 U5231 ( .A1(n6347), .A2(n6161), .ZN(n4368) );
  NOR2_X1 U5232 ( .A1(n6346), .A2(n4369), .ZN(BUS_ADDR_OUTBUS[15]) );
  NAND2_X1 U5233 ( .A1(n6347), .A2(n6169), .ZN(n4369) );
  NOR2_X1 U5234 ( .A1(n6346), .A2(n4370), .ZN(BUS_ADDR_OUTBUS[14]) );
  NAND2_X1 U5235 ( .A1(n6347), .A2(n6180), .ZN(n4370) );
  NOR2_X1 U5236 ( .A1(n6346), .A2(n4371), .ZN(BUS_ADDR_OUTBUS[13]) );
  NAND2_X1 U5237 ( .A1(n6347), .A2(n6187), .ZN(n4371) );
  NOR2_X1 U5238 ( .A1(n4372), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[12]) );
  NAND2_X1 U5239 ( .A1(n6347), .A2(n6203), .ZN(n4372) );
  NOR2_X1 U5240 ( .A1(n4373), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[11]) );
  NAND2_X1 U5241 ( .A1(n6347), .A2(n6204), .ZN(n4373) );
  NOR2_X1 U5242 ( .A1(n4374), .A2(n6346), .ZN(BUS_ADDR_OUTBUS[10]) );
  NAND2_X1 U5243 ( .A1(n6347), .A2(n6205), .ZN(n4374) );
  NAND2_X1 U5244 ( .A1(n6348), .A2(n6350), .ZN(n6349) );
  INV_X1 U5245 ( .A(\UUT/Mpath/the_alu/N492 ), .ZN(n6350) );
  NOR2_X1 U5247 ( .A1(n6346), .A2(n4375), .ZN(BUS_ADDR_OUTBUS[0]) );
  NAND2_X1 U5248 ( .A1(D_ADDR_OUTBUS[0]), .A2(\localbus/N50 ), .ZN(n4375) );
  AND2_X1 U5249 ( .A1(\UUT/N3 ), .A2(\UUT/daddr_out [0]), .ZN(D_ADDR_OUTBUS[0]) );
  OAI21_X1 U5250 ( .B1(\UUT/Mpath/the_alu/N492 ), .B2(n6352), .A(n6353), .ZN(
        n6351) );
  NAND2_X1 U5251 ( .A1(\UUT/Mpath/the_alu/N125 ), .A2(\UUT/Mpath/the_alu/N492 ), .ZN(n6353) );
  AOI22_X1 U5252 ( .A1(n6354), .A2(\UUT/Mpath/the_alu/N485 ), .B1(
        \UUT/Mpath/the_alu/N157 ), .B2(\UUT/Mpath/the_alu/N486 ), .ZN(n6352)
         );
  OAI21_X1 U5253 ( .B1(\UUT/Mpath/the_alu/N480 ), .B2(n6355), .A(n6356), .ZN(
        n6354) );
  NAND2_X1 U5254 ( .A1(\UUT/Mpath/the_alu/N189 ), .A2(\UUT/Mpath/the_alu/N480 ), .ZN(n6356) );
  AOI22_X1 U5255 ( .A1(\UUT/Mpath/the_alu/N221 ), .A2(\UUT/Mpath/the_alu/N474 ), .B1(\UUT/Mpath/the_alu/N473 ), .B2(n6525), .ZN(n6355) );
  BUF_X2 U5257 ( .A(dmem_ishalf), .Z(n6357) );
  BUF_X2 U5258 ( .A(dmem_ishalf), .Z(n6358) );
  BUF_X2 U5259 ( .A(dmem_ishalf), .Z(n6359) );
  BUF_X2 U5260 ( .A(dmem_ishalf), .Z(n6360) );
  BUF_X2 U5261 ( .A(D_ADDR_OUTBUS[1]), .Z(n6361) );
  BUF_X2 U5262 ( .A(dmem_isbyte), .Z(n6362) );
  BUF_X2 U5263 ( .A(dmem_isbyte), .Z(n6363) );
  BUF_X2 U5264 ( .A(dmem_isbyte), .Z(N13) );
  BUF_X2 U5265 ( .A(dmem_isbyte), .Z(N11) );
  BUF_X2 U5266 ( .A(dmem_isbyte), .Z(N9) );
  BUF_X2 U5267 ( .A(dmem_isbyte), .Z(N7) );
  BUF_X2 U5268 ( .A(dmem_ishalf), .Z(N3) );
  BUF_X2 U5269 ( .A(D_ADDR_OUTBUS[1]), .Z(N2) );
  BUF_X2 U5270 ( .A(dmem_ishalf), .Z(N0) );
  INV_X2 U5271 ( .A(n6363), .ZN(N1) );
  INV_X2 U5272 ( .A(n6362), .ZN(N4) );
  INV_X2 U5273 ( .A(n6361), .ZN(N5) );
  INV_X2 U5274 ( .A(n6360), .ZN(N6) );
  INV_X2 U5275 ( .A(n6359), .ZN(N8) );
  INV_X2 U5276 ( .A(n6358), .ZN(N10) );
  INV_X2 U5277 ( .A(n6357), .ZN(N12) );
  up_island_DW01_add_0 \UUT/Mpath/the_mult/accumulate/add_391  ( .A({1'b0, 
        \UUT/Mpath/the_mult/acc_out[63] , \UUT/Mpath/the_mult/acc_out[62] , 
        \UUT/Mpath/the_mult/acc_out[61] , \UUT/Mpath/the_mult/acc_out[60] , 
        \UUT/Mpath/the_mult/acc_out[59] , \UUT/Mpath/the_mult/acc_out[58] , 
        \UUT/Mpath/the_mult/acc_out[57] , \UUT/Mpath/the_mult/acc_out[56] , 
        \UUT/Mpath/the_mult/acc_out[55] , \UUT/Mpath/the_mult/acc_out[54] , 
        \UUT/Mpath/the_mult/acc_out[53] , \UUT/Mpath/the_mult/acc_out[52] , 
        \UUT/Mpath/the_mult/acc_out[51] , \UUT/Mpath/the_mult/acc_out[50] , 
        \UUT/Mpath/the_mult/acc_out[49] , \UUT/Mpath/the_mult/acc_out[48] , 
        \UUT/Mpath/the_mult/acc_out[47] , \UUT/Mpath/the_mult/acc_out[46] , 
        \UUT/Mpath/the_mult/acc_out[45] , \UUT/Mpath/the_mult/acc_out[44] , 
        \UUT/Mpath/the_mult/acc_out[43] , \UUT/Mpath/the_mult/acc_out[42] , 
        \UUT/Mpath/the_mult/acc_out[41] , \UUT/Mpath/the_mult/acc_out[40] , 
        \UUT/Mpath/the_mult/acc_out[39] , \UUT/Mpath/the_mult/acc_out[38] , 
        \UUT/Mpath/the_mult/acc_out[37] , \UUT/Mpath/the_mult/acc_out[36] , 
        \UUT/Mpath/the_mult/acc_out[35] , \UUT/Mpath/the_mult/acc_out[34] , 
        \UUT/Mpath/the_mult/acc_out[33] , \UUT/Mpath/the_mult/acc_out[32] , 
        \UUT/Mpath/the_mult/acc_out[31] , \UUT/Mpath/the_mult/acc_out[30] , 
        \UUT/Mpath/the_mult/acc_out[29] , \UUT/Mpath/the_mult/acc_out[28] , 
        \UUT/Mpath/the_mult/acc_out[27] , \UUT/Mpath/the_mult/acc_out[26] , 
        \UUT/Mpath/the_mult/acc_out[25] , \UUT/Mpath/the_mult/acc_out[24] , 
        \UUT/Mpath/the_mult/acc_out[23] , \UUT/Mpath/the_mult/acc_out[22] , 
        \UUT/Mpath/the_mult/acc_out[21] , \UUT/Mpath/the_mult/acc_out[20] , 
        \UUT/Mpath/the_mult/acc_out[19] , \UUT/Mpath/the_mult/acc_out[18] , 
        \UUT/Mpath/the_mult/acc_out[17] , \UUT/Mpath/the_mult/acc_out[16] , 
        \UUT/Mpath/the_mult/acc_out[15] , \UUT/Mpath/the_mult/acc_out[14] , 
        \UUT/Mpath/the_mult/acc_out[13] , \UUT/Mpath/the_mult/acc_out[12] , 
        \UUT/Mpath/the_mult/acc_out[11] , \UUT/Mpath/the_mult/acc_out[10] , 
        \UUT/Mpath/the_mult/acc_out[9] , \UUT/Mpath/the_mult/acc_out[8] , 
        \UUT/Mpath/the_mult/acc_out[7] , \UUT/Mpath/the_mult/acc_out[6] , 
        \UUT/Mpath/the_mult/acc_out[5] , \UUT/Mpath/the_mult/acc_out[4] , 
        \UUT/Mpath/the_mult/acc_out[3] , \UUT/Mpath/the_mult/acc_out[2] , 
        \UUT/Mpath/the_mult/acc_out[1] , \UUT/Mpath/the_mult/acc_out[0] }), 
        .B({1'b0, \UUT/Mpath/the_mult/Mult_out[63] , 
        \UUT/Mpath/the_mult/Mult_out[62] , \UUT/Mpath/the_mult/Mult_out[61] , 
        \UUT/Mpath/the_mult/Mult_out[60] , \UUT/Mpath/the_mult/Mult_out[59] , 
        \UUT/Mpath/the_mult/Mult_out[58] , \UUT/Mpath/the_mult/Mult_out[57] , 
        \UUT/Mpath/the_mult/Mult_out[56] , \UUT/Mpath/the_mult/Mult_out[55] , 
        \UUT/Mpath/the_mult/Mult_out[54] , \UUT/Mpath/the_mult/Mult_out[53] , 
        \UUT/Mpath/the_mult/Mult_out[52] , \UUT/Mpath/the_mult/Mult_out[51] , 
        \UUT/Mpath/the_mult/Mult_out[50] , \UUT/Mpath/the_mult/Mult_out[49] , 
        \UUT/Mpath/the_mult/Mult_out[48] , \UUT/Mpath/the_mult/Mult_out[47] , 
        \UUT/Mpath/the_mult/Mult_out[46] , \UUT/Mpath/the_mult/Mult_out[45] , 
        \UUT/Mpath/the_mult/Mult_out[44] , \UUT/Mpath/the_mult/Mult_out[43] , 
        \UUT/Mpath/the_mult/Mult_out[42] , \UUT/Mpath/the_mult/Mult_out[41] , 
        \UUT/Mpath/the_mult/Mult_out[40] , \UUT/Mpath/the_mult/Mult_out[39] , 
        \UUT/Mpath/the_mult/Mult_out[38] , \UUT/Mpath/the_mult/Mult_out[37] , 
        \UUT/Mpath/the_mult/Mult_out[36] , \UUT/Mpath/the_mult/Mult_out[35] , 
        \UUT/Mpath/the_mult/Mult_out[34] , \UUT/Mpath/the_mult/Mult_out[33] , 
        \UUT/Mpath/the_mult/Mult_out[32] , \UUT/Mpath/the_mult/Mult_out[31] , 
        \UUT/Mpath/the_mult/Mult_out[30] , \UUT/Mpath/the_mult/Mult_out[29] , 
        \UUT/Mpath/the_mult/Mult_out[28] , \UUT/Mpath/the_mult/Mult_out[27] , 
        \UUT/Mpath/the_mult/Mult_out[26] , \UUT/Mpath/the_mult/Mult_out[25] , 
        \UUT/Mpath/the_mult/Mult_out[24] , \UUT/Mpath/the_mult/Mult_out[23] , 
        \UUT/Mpath/the_mult/Mult_out[22] , \UUT/Mpath/the_mult/Mult_out[21] , 
        \UUT/Mpath/the_mult/Mult_out[20] , \UUT/Mpath/the_mult/Mult_out[19] , 
        \UUT/Mpath/the_mult/Mult_out[18] , \UUT/Mpath/the_mult/Mult_out[17] , 
        \UUT/Mpath/the_mult/Mult_out[16] , \UUT/Mpath/the_mult/Mult_out[15] , 
        \UUT/Mpath/the_mult/Mult_out[14] , \UUT/Mpath/the_mult/Mult_out[13] , 
        \UUT/Mpath/the_mult/Mult_out[12] , \UUT/Mpath/the_mult/Mult_out[11] , 
        \UUT/Mpath/the_mult/Mult_out[10] , \UUT/Mpath/the_mult/Mult_out[9] , 
        \UUT/Mpath/the_mult/Mult_out[8] , \UUT/Mpath/the_mult/Mult_out[7] , 
        \UUT/Mpath/the_mult/Mult_out[6] , \UUT/Mpath/the_mult/Mult_out[5] , 
        \UUT/Mpath/the_mult/Mult_out[4] , \UUT/Mpath/the_mult/Mult_out[3] , 
        \UUT/Mpath/the_mult/Mult_out[2] , \UUT/Mpath/the_mult/Mult_out[1] , 
        \UUT/Mpath/the_mult/Mult_out[0] }), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, \UUT/Mpath/the_mult/Mad_out }) );
  up_island_DW01_add_1 \UUT/Mcontrol/Nextpc_decoding/bta_calc/add_391  ( .A({
        1'b0, \UUT/Mcontrol/f_currpc }), .B({1'b0, \UUT/break_code[23] , 
        \UUT/break_code[22] , \UUT/break_code[21] , \UUT/break_code[20] , 
        \UUT/break_code[19] , \UUT/break_code[18] , \UUT/break_code[17] , 
        \UUT/break_code[16] , \UUT/break_code[15] , \UUT/break_code[14] , 
        \UUT/break_code[13] , \UUT/break_code[12] , \UUT/break_code[11] , 
        \UUT/break_code[10] , \UUT/break_code[9] , \UUT/break_code[8] , 
        \UUT/break_code[7] , \UUT/break_code[6] , \UUT/break_code[5] , 
        \UUT/break_code[4] , \UUT/break_code[3] , \UUT/break_code[2] , 
        \UUT/break_code[1] , \UUT/break_code[0] }), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, \UUT/Mcontrol/Nextpc_decoding/Bta }) );
  up_island_DW01_add_2 \UUT/Mcontrol/Nextpc_decoding/incr/add_391  ( .A({1'b0, 
        \UUT/Mcontrol/f_currpc }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__2, \UUT/jar_in }) );
  up_island_DW01_cmp6_0 r771 ( .A({n6475, \UUT/branch_rega [30:22], n6464, 
        \UUT/branch_rega [20:0]}), .B(\UUT/branch_regb ), .TC(1'b0), .EQ(
        \UUT/Mcontrol/Nextpc_decoding/N22 ), .NE(
        \UUT/Mcontrol/Nextpc_decoding/N25 ) );
  up_island_DW01_sub_0 \UUT/Mpath/the_alu/sub_96  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, 
        \UUT/Mpath/out_regA[0] }), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , 
        \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n6897, n6898, n6899, 
        \UUT/Mpath/out_regB[1] , \UUT/Mpath/out_regB[0] }), .CI(1'b0), .DIFF({
        \UUT/Mpath/the_alu/diff[31] , \UUT/Mpath/the_alu/diff[30] , 
        \UUT/Mpath/the_alu/diff[29] , \UUT/Mpath/the_alu/diff[28] , 
        \UUT/Mpath/the_alu/diff[27] , \UUT/Mpath/the_alu/diff[26] , 
        \UUT/Mpath/the_alu/diff[25] , \UUT/Mpath/the_alu/diff[24] , 
        \UUT/Mpath/the_alu/diff[23] , \UUT/Mpath/the_alu/diff[22] , 
        \UUT/Mpath/the_alu/diff[21] , \UUT/Mpath/the_alu/diff[20] , 
        \UUT/Mpath/the_alu/diff[19] , \UUT/Mpath/the_alu/diff[18] , 
        \UUT/Mpath/the_alu/diff[17] , \UUT/Mpath/the_alu/diff[16] , 
        \UUT/Mpath/the_alu/diff[15] , \UUT/Mpath/the_alu/diff[14] , 
        \UUT/Mpath/the_alu/diff[13] , \UUT/Mpath/the_alu/diff[12] , 
        \UUT/Mpath/the_alu/diff[11] , \UUT/Mpath/the_alu/diff[10] , 
        \UUT/Mpath/the_alu/diff[9] , \UUT/Mpath/the_alu/diff[8] , 
        \UUT/Mpath/the_alu/diff[7] , \UUT/Mpath/the_alu/diff[6] , 
        \UUT/Mpath/the_alu/diff[5] , \UUT/Mpath/the_alu/diff[4] , 
        \UUT/Mpath/the_alu/diff[3] , \UUT/Mpath/the_alu/diff[2] , 
        \UUT/Mpath/the_alu/diff[1] , \UUT/Mpath/the_alu/diff[0] }) );
  up_island_DW01_add_3 \UUT/Mpath/the_alu/add_95  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, 
        \UUT/Mpath/out_regA[0] }), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , 
        \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n6897, n6898, n6899, 
        \UUT/Mpath/out_regB[1] , \UUT/Mpath/out_regB[0] }), .CI(1'b0), .SUM({
        \UUT/Mpath/the_alu/sum[31] , \UUT/Mpath/the_alu/sum[30] , 
        \UUT/Mpath/the_alu/sum[29] , \UUT/Mpath/the_alu/sum[28] , 
        \UUT/Mpath/the_alu/sum[27] , \UUT/Mpath/the_alu/sum[26] , 
        \UUT/Mpath/the_alu/sum[25] , \UUT/Mpath/the_alu/sum[24] , 
        \UUT/Mpath/the_alu/sum[23] , \UUT/Mpath/the_alu/sum[22] , 
        \UUT/Mpath/the_alu/sum[21] , \UUT/Mpath/the_alu/sum[20] , 
        \UUT/Mpath/the_alu/sum[19] , \UUT/Mpath/the_alu/sum[18] , 
        \UUT/Mpath/the_alu/sum[17] , \UUT/Mpath/the_alu/sum[16] , 
        \UUT/Mpath/the_alu/sum[15] , \UUT/Mpath/the_alu/sum[14] , 
        \UUT/Mpath/the_alu/sum[13] , \UUT/Mpath/the_alu/sum[12] , 
        \UUT/Mpath/the_alu/sum[11] , \UUT/Mpath/the_alu/sum[10] , 
        \UUT/Mpath/the_alu/sum[9] , \UUT/Mpath/the_alu/sum[8] , 
        \UUT/Mpath/the_alu/sum[7] , \UUT/Mpath/the_alu/sum[6] , 
        \UUT/Mpath/the_alu/sum[5] , \UUT/Mpath/the_alu/sum[4] , 
        \UUT/Mpath/the_alu/sum[3] , \UUT/Mpath/the_alu/sum[2] , 
        \UUT/Mpath/the_alu/sum[1] , \UUT/Mpath/the_alu/sum[0] }) );
  up_island_DW_mult_tc_1 \UUT/Mpath/the_mult/mult_186  ( .a({
        \UUT/Mpath/the_mult/x_operand1[31] , 
        \UUT/Mpath/the_mult/x_operand1[30] , 
        \UUT/Mpath/the_mult/x_operand1[29] , 
        \UUT/Mpath/the_mult/x_operand1[28] , 
        \UUT/Mpath/the_mult/x_operand1[27] , 
        \UUT/Mpath/the_mult/x_operand1[26] , 
        \UUT/Mpath/the_mult/x_operand1[25] , 
        \UUT/Mpath/the_mult/x_operand1[24] , 
        \UUT/Mpath/the_mult/x_operand1[23] , 
        \UUT/Mpath/the_mult/x_operand1[22] , 
        \UUT/Mpath/the_mult/x_operand1[21] , 
        \UUT/Mpath/the_mult/x_operand1[20] , 
        \UUT/Mpath/the_mult/x_operand1[19] , 
        \UUT/Mpath/the_mult/x_operand1[18] , 
        \UUT/Mpath/the_mult/x_operand1[17] , 
        \UUT/Mpath/the_mult/x_operand1[16] , 
        \UUT/Mpath/the_mult/x_operand1[15] , 
        \UUT/Mpath/the_mult/x_operand1[14] , 
        \UUT/Mpath/the_mult/x_operand1[13] , 
        \UUT/Mpath/the_mult/x_operand1[12] , 
        \UUT/Mpath/the_mult/x_operand1[11] , 
        \UUT/Mpath/the_mult/x_operand1[10] , 
        \UUT/Mpath/the_mult/x_operand1[9] , \UUT/Mpath/the_mult/x_operand1[8] , 
        \UUT/Mpath/the_mult/x_operand1[7] , \UUT/Mpath/the_mult/x_operand1[6] , 
        \UUT/Mpath/the_mult/x_operand1[5] , \UUT/Mpath/the_mult/x_operand1[4] , 
        \UUT/Mpath/the_mult/x_operand1[3] , \UUT/Mpath/the_mult/x_operand1[2] , 
        \UUT/Mpath/the_mult/x_operand1[1] , \UUT/Mpath/the_mult/x_operand1[0] }), .b(\UUT/Mpath/the_mult/x_operand2 ), .product({
        \UUT/Mpath/the_mult/x_mult_out[63] , 
        \UUT/Mpath/the_mult/x_mult_out[62] , 
        \UUT/Mpath/the_mult/x_mult_out[61] , 
        \UUT/Mpath/the_mult/x_mult_out[60] , 
        \UUT/Mpath/the_mult/x_mult_out[59] , 
        \UUT/Mpath/the_mult/x_mult_out[58] , 
        \UUT/Mpath/the_mult/x_mult_out[57] , 
        \UUT/Mpath/the_mult/x_mult_out[56] , 
        \UUT/Mpath/the_mult/x_mult_out[55] , 
        \UUT/Mpath/the_mult/x_mult_out[54] , 
        \UUT/Mpath/the_mult/x_mult_out[53] , 
        \UUT/Mpath/the_mult/x_mult_out[52] , 
        \UUT/Mpath/the_mult/x_mult_out[51] , 
        \UUT/Mpath/the_mult/x_mult_out[50] , 
        \UUT/Mpath/the_mult/x_mult_out[49] , 
        \UUT/Mpath/the_mult/x_mult_out[48] , 
        \UUT/Mpath/the_mult/x_mult_out[47] , 
        \UUT/Mpath/the_mult/x_mult_out[46] , 
        \UUT/Mpath/the_mult/x_mult_out[45] , 
        \UUT/Mpath/the_mult/x_mult_out[44] , 
        \UUT/Mpath/the_mult/x_mult_out[43] , 
        \UUT/Mpath/the_mult/x_mult_out[42] , 
        \UUT/Mpath/the_mult/x_mult_out[41] , 
        \UUT/Mpath/the_mult/x_mult_out[40] , 
        \UUT/Mpath/the_mult/x_mult_out[39] , 
        \UUT/Mpath/the_mult/x_mult_out[38] , 
        \UUT/Mpath/the_mult/x_mult_out[37] , 
        \UUT/Mpath/the_mult/x_mult_out[36] , 
        \UUT/Mpath/the_mult/x_mult_out[35] , 
        \UUT/Mpath/the_mult/x_mult_out[34] , 
        \UUT/Mpath/the_mult/x_mult_out[33] , 
        \UUT/Mpath/the_mult/x_mult_out[32] , 
        \UUT/Mpath/the_mult/x_mult_out[31] , 
        \UUT/Mpath/the_mult/x_mult_out[30] , 
        \UUT/Mpath/the_mult/x_mult_out[29] , 
        \UUT/Mpath/the_mult/x_mult_out[28] , 
        \UUT/Mpath/the_mult/x_mult_out[27] , 
        \UUT/Mpath/the_mult/x_mult_out[26] , 
        \UUT/Mpath/the_mult/x_mult_out[25] , 
        \UUT/Mpath/the_mult/x_mult_out[24] , 
        \UUT/Mpath/the_mult/x_mult_out[23] , 
        \UUT/Mpath/the_mult/x_mult_out[22] , 
        \UUT/Mpath/the_mult/x_mult_out[21] , 
        \UUT/Mpath/the_mult/x_mult_out[20] , 
        \UUT/Mpath/the_mult/x_mult_out[19] , 
        \UUT/Mpath/the_mult/x_mult_out[18] , 
        \UUT/Mpath/the_mult/x_mult_out[17] , 
        \UUT/Mpath/the_mult/x_mult_out[16] , 
        \UUT/Mpath/the_mult/x_mult_out[15] , 
        \UUT/Mpath/the_mult/x_mult_out[14] , 
        \UUT/Mpath/the_mult/x_mult_out[13] , 
        \UUT/Mpath/the_mult/x_mult_out[12] , 
        \UUT/Mpath/the_mult/x_mult_out[11] , 
        \UUT/Mpath/the_mult/x_mult_out[10] , 
        \UUT/Mpath/the_mult/x_mult_out[9] , \UUT/Mpath/the_mult/x_mult_out[8] , 
        \UUT/Mpath/the_mult/x_mult_out[7] , \UUT/Mpath/the_mult/x_mult_out[6] , 
        \UUT/Mpath/the_mult/x_mult_out[5] , \UUT/Mpath/the_mult/x_mult_out[4] , 
        \UUT/Mpath/the_mult/x_mult_out[3] , \UUT/Mpath/the_mult/x_mult_out[2] , 
        \UUT/Mpath/the_mult/x_mult_out[1] , \UUT/Mpath/the_mult/x_mult_out[0] }) );
  up_island_DW_rightsh_1 \UUT/Mpath/the_shift/S_SRL/srl_128  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, n6525}), .SH(
        {n6896, n6898, n6899, n6900, n6675}), .B(\UUT/Mpath/the_shift/sh_srl ), 
        .DATA_TC(1'b0) );
  up_island_DW_sra_1 \UUT/Mpath/the_shift/S_SRA/sra_106  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, n6525}), .SH(
        {n6896, n6898, n6899, \UUT/Mpath/out_regB[1] , n6675}), .B(
        \UUT/Mpath/the_shift/sh_sra ), .SH_TC(1'b0) );
  up_island_DW_rbsh_1 \UUT/Mpath/the_shift/S_ROR/ror_81  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, n6525}), .SH(
        {n6897, n6898, n6899, n6900, n6675}), .B(\UUT/Mpath/the_shift/sh_ror ), 
        .SH_TC(1'b0) );
  up_island_DW01_bsh_1 \UUT/Mpath/the_shift/S_ROL/rol_55  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, n6525}), .SH(
        {n6895, n6898, n6899, \UUT/Mpath/out_regB[1] , n6675}), .B(
        \UUT/Mpath/the_shift/sh_rol ) );
  up_island_DW_leftsh_1 \UUT/Mpath/the_shift/S_SLL/sll_150  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , 
        \UUT/Mpath/out_regA[13] , \UUT/Mpath/out_regA[12] , 
        \UUT/Mpath/out_regA[11] , \UUT/Mpath/out_regA[10] , 
        \UUT/Mpath/out_regA[9] , \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , \UUT/Mpath/out_regA[6] , 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , n6450, n6525}), .SH(
        {n6895, n6898, n6899, n6900, n6675}), .B(\UUT/Mpath/the_shift/sh_sll )
         );
  up_island_DW_cmp_0 \UUT/Mpath/the_alu/lt_114  ( .A({\UUT/Mpath/out_regA[31] , 
        \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[29] , 
        \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[27] , 
        \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[25] , 
        \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[23] , 
        \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[21] , 
        \UUT/Mpath/out_regA[20] , \UUT/Mpath/out_regA[19] , 
        \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[17] , 
        \UUT/Mpath/out_regA[16] , \UUT/Mpath/out_regA[15] , 
        \UUT/Mpath/out_regA[14] , \UUT/Mpath/out_regA[13] , 
        \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[11] , 
        \UUT/Mpath/out_regA[10] , \UUT/Mpath/out_regA[9] , 
        \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[7] , 
        \UUT/Mpath/out_regA[6] , \UUT/Mpath/out_regA[5] , 
        \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[3] , 
        \UUT/Mpath/out_regA[2] , n6450, n6525}), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , 
        \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n6897, n6898, n6899, 
        n6900, n6675}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(\UUT/Mpath/the_alu/N91 ) );
  up_island_DW_cmp_1 \UUT/Mpath/the_alu/lt_120  ( .A({\UUT/Mpath/out_regA[31] , 
        \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[29] , 
        \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[27] , 
        \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[25] , 
        \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[23] , 
        \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[21] , 
        \UUT/Mpath/out_regA[20] , \UUT/Mpath/out_regA[19] , 
        \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[17] , 
        \UUT/Mpath/out_regA[16] , \UUT/Mpath/out_regA[15] , 
        \UUT/Mpath/out_regA[14] , \UUT/Mpath/out_regA[13] , 
        \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[11] , 
        \UUT/Mpath/out_regA[10] , \UUT/Mpath/out_regA[9] , 
        \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[7] , 
        \UUT/Mpath/out_regA[6] , \UUT/Mpath/out_regA[5] , 
        \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[3] , 
        \UUT/Mpath/out_regA[2] , n6450, n6525}), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , 
        \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n6897, n6898, n6899, 
        n6900, n6675}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(\UUT/Mpath/the_alu/N93 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[17]  ( .D(n3169), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[17] ), .QN(
        \UUT/Mpath/the_alu/N49 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[23]  ( .D(n3776), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[23] ), .QN(
        \UUT/Mpath/the_alu/N37 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[20]  ( .D(n3044), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[20] ), .QN(
        \UUT/Mpath/the_alu/N44 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[20]  ( .D(n3049), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[20] ), .QN(
        \UUT/Mpath/the_alu/N43 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[19]  ( .D(n3084), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[19] ), .QN(
        \UUT/Mpath/the_alu/N46 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[19]  ( .D(n3089), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[19] ), .QN(
        \UUT/Mpath/the_alu/N45 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[7]  ( .D(n3501), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[7] ), .QN(
        \UUT/Mpath/the_alu/N69 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[8]  ( .D(n3492), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[8] ), .QN(
        \UUT/Mpath/the_alu/N67 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[14]  ( .D(n3289), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[14] ), .QN(
        \UUT/Mpath/the_alu/N55 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[29]  ( .D(n3943), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[29] ), .QN(
        \UUT/Mpath/the_alu/N25 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[13]  ( .D(n3329), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[13] ), .QN(
        \UUT/Mpath/the_alu/N57 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[25]  ( .D(n2918), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[25] ), .QN(
        \UUT/Mpath/the_alu/N34 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[25]  ( .D(n3811), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[25] ), .QN(
        \UUT/Mpath/the_alu/N33 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[24]  ( .D(n2924), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[24] ), .QN(
        \UUT/Mpath/the_alu/N36 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[24]  ( .D(n2929), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[24] ), .QN(
        \UUT/Mpath/the_alu/N35 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[27]  ( .D(n2906), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[27] ), .QN(
        \UUT/Mpath/the_alu/N30 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[27]  ( .D(n3877), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[27] ), .QN(
        \UUT/Mpath/the_alu/N29 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[6]  ( .D(n3541), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[6] ), .QN(
        \UUT/Mpath/the_alu/N71 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[12]  ( .D(n3369), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[12] ), .QN(
        \UUT/Mpath/the_alu/N59 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[30]  ( .D(n3981), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[30] ), .QN(
        \UUT/Mpath/the_alu/N23 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[18]  ( .D(n3124), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[18] ), .QN(
        \UUT/Mpath/the_alu/N48 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[18]  ( .D(n3129), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[18] ), .QN(
        \UUT/Mpath/the_alu/N47 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[2]  ( .D(n3701), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[2] ), .QN(
        \UUT/Mpath/the_alu/N79 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[5]  ( .D(n3576), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[5] ), .QN(
        \UUT/Mpath/the_alu/N74 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[5]  ( .D(n3581), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[5] ), .QN(
        \UUT/Mpath/the_alu/N73 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[26]  ( .D(n2912), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[26] ), .QN(
        \UUT/Mpath/the_alu/N32 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[26]  ( .D(n3844), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[26] ), .QN(
        \UUT/Mpath/the_alu/N31 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[17]  ( .D(n3164), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[17] ), .QN(
        \UUT/Mpath/the_alu/N50 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[23]  ( .D(n4014), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[23] ), .QN(
        \UUT/Mpath/the_alu/N38 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[28]  ( .D(n2900), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[28] ), .QN(
        \UUT/Mpath/the_alu/N28 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[28]  ( .D(n3910), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[28] ), .QN(
        \UUT/Mpath/the_alu/N27 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[3]  ( .D(n3661), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[3] ), .QN(
        \UUT/Mpath/the_alu/N77 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[10]  ( .D(n3446), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[10] ), .QN(
        \UUT/Mpath/the_alu/N63 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[9]  ( .D(n3454), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[9] ), .QN(
        \UUT/Mpath/the_alu/N65 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[31]  ( .D(n4327), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[31] ), .QN(
        \UUT/Mpath/the_alu/N22 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[31]  ( .D(n4057), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[31] ), .QN(
        \UUT/Mpath/the_alu/N21 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[4]  ( .D(n3621), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[4] ), .QN(
        \UUT/Mpath/the_alu/N75 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[16]  ( .D(n3204), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[16] ), .QN(
        \UUT/Mpath/the_alu/N52 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[16]  ( .D(n3209), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[16] ), .QN(
        \UUT/Mpath/the_alu/N51 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[22]  ( .D(n2964), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[22] ), .QN(
        \UUT/Mpath/the_alu/N40 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[22]  ( .D(n2969), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[22] ), .QN(
        \UUT/Mpath/the_alu/N39 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[11]  ( .D(n3409), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[11] ), .QN(
        \UUT/Mpath/the_alu/N61 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[21]  ( .D(n3009), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[21] ), .QN(
        \UUT/Mpath/the_alu/N41 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[15]  ( .D(n3244), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[15] ), .QN(
        \UUT/Mpath/the_alu/N54 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[15]  ( .D(n3249), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[15] ), .QN(
        \UUT/Mpath/the_alu/N53 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[21]  ( .D(n3004), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[21] ), .QN(
        \UUT/Mpath/the_alu/N42 ) );
  DFFR_X2 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[50]  ( .D(n4307), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[50] ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[14]  ( .D(n3284), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[14] ), .QN(
        \UUT/Mpath/the_alu/N56 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[13]  ( .D(n3324), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[13] ), .QN(
        \UUT/Mpath/the_alu/N58 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[12]  ( .D(n3364), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[12] ), .QN(
        \UUT/Mpath/the_alu/N60 ) );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[11]  ( .D(n3404), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[11] ), .QN(
        \UUT/Mpath/the_alu/N62 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[0]  ( .D(n4256), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[0] ), .QN(
        \UUT/Mpath/the_alu/N83 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[1]  ( .D(n3740), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[1] ), .QN(
        \UUT/Mpath/the_alu/N81 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[5]  ( .D(n3574), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [5]), .QN(
        n2685) );
  DFFS_X2 \UUT/Mcontrol/Program_counter/out_pc_reg[18]  ( .D(n3123), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [18]), .QN(
        n2651) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[31]  ( .D(n4329), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[63] ), .QN(
        n5685) );
  NAND2_X2 syn1555 ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(
        \UUT/Mpath/the_mult/N231 ), .ZN(n6440) );
  INV_X2 syn1525 ( .A(n6445), .ZN(net54953) );
  NAND3_X1 syn1524 ( .A1(n6436), .A2(n6444), .A3(\localbus/N199 ), .ZN(n6445)
         );
  NAND2_X2 syn1522 ( .A1(n6442), .A2(n6441), .ZN(n6444) );
  INV_X2 syn868 ( .A(n6433), .ZN(n139) );
  INV_X2 syn831 ( .A(\UUT/Mpath/the_mult/m_mul_command[3] ), .ZN(n6438) );
  INV_X2 syn768 ( .A(n6443), .ZN(n137) );
  NAND2_X2 syn767 ( .A1(n975), .A2(n6432), .ZN(n6443) );
  INV_X2 syn763 ( .A(\UUT/Mpath/the_mult/N313 ), .ZN(n6427) );
  INV_X2 syn761 ( .A(\localbus/N329 ), .ZN(n6442) );
  INV_X2 syn759 ( .A(\localbus/N331 ), .ZN(n6441) );
  NOR2_X2 syn749 ( .A1(n6426), .A2(n6432), .ZN(n6435) );
  NOR2_X2 syn745 ( .A1(n6429), .A2(net54953), .ZN(n6434) );
  AND2_X2 syn743 ( .A1(n6439), .A2(n6440), .ZN(n6430) );
  NOR2_X2 syn741 ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/m_mul_command[1] ), .ZN(n6439) );
  AND2_X2 syn739 ( .A1(n6437), .A2(n6438), .ZN(n6431) );
  NOR2_X2 syn737 ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(
        \UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(n6437) );
  INV_X2 syn727 ( .A(net87679), .ZN(n6428) );
  NAND3_X1 syn725 ( .A1(n6434), .A2(n6435), .A3(n6427), .ZN(n6433) );
  INV_X2 syn722 ( .A(\UUT/Mpath/the_mult/N285 ), .ZN(n6432) );
  NAND2_X2 syn721 ( .A1(n6430), .A2(n6431), .ZN(n6426) );
  INV_X2 syn720 ( .A(n5413), .ZN(n6429) );
  NAND3_X1 net89067 ( .A1(\UUT/Mpath/the_mult/N285 ), .A2(n6426), .A3(n6427), 
        .ZN(n1183) );
  DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[1]  ( .D(n3735), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [1]), .QN(
        n2698) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[15]  ( .D(n3243), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [15]), .QN(
        n2660) );
  DFFS_X2 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MR]  ( .D(n4060), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/m_mem_command[MR] ), .QN(n5710)
         );
  NOR2_X1 U5278 ( .A1(\localbus/c2_op[MASTER] ), .A2(BUS_NREADY), .ZN(n6436)
         );
  INV_X1 U5279 ( .A(\UUT/branch_rega [4]), .ZN(n6868) );
  INV_X1 U5280 ( .A(\UUT/branch_rega [4]), .ZN(n6874) );
  OR2_X1 U5281 ( .A1(n6794), .A2(\UUT/branch_rega [4]), .ZN(n6787) );
  NOR3_X2 U5282 ( .A1(n933), .A2(n6209), .A3(n2070), .ZN(n2074) );
  NAND2_X2 U5283 ( .A1(n147), .A2(n175), .ZN(n71) );
  OR2_X1 U5284 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N115 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N116 ) );
  OR2_X1 U5285 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N263 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N264 ) );
  OR2_X1 U5286 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N251 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N252 ) );
  OR2_X1 U5287 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N257 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N258 ) );
  OR2_X1 U5288 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N123 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N124 ) );
  INV_X1 U5289 ( .A(\UUT/Mcontrol/d_jump_type[1] ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N224 ) );
  OR2_X1 U5290 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N245 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N246 ) );
  OR2_X1 U5291 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N61 ), .ZN(\UUT/Mcontrol/st_logic/N62 ) );
  OR2_X1 U5292 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N68 ), .ZN(\UUT/Mcontrol/st_logic/N69 ) );
  OR2_X1 U5293 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N106 ), .ZN(\UUT/Mcontrol/st_logic/N107 ) );
  INV_X1 U5294 ( .A(\UUT/Mcontrol/d_jump_type[1] ), .ZN(
        \UUT/Mcontrol/st_logic/N90 ) );
  OR2_X1 U5295 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N86 ), .ZN(\UUT/Mcontrol/st_logic/N87 ) );
  OR2_X1 U5296 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N74 ), .ZN(\UUT/Mcontrol/st_logic/N75 ) );
  OR2_X1 U5297 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N80 ), .ZN(\UUT/Mcontrol/st_logic/N81 ) );
  NOR2_X2 U5298 ( .A1(n5896), .A2(n6322), .ZN(\UUT/rs1_addr [1]) );
  INV_X1 U5299 ( .A(\UUT/branch_rega [5]), .ZN(n6854) );
  INV_X1 U5300 ( .A(\UUT/branch_rega [0]), .ZN(n6832) );
  INV_X1 U5301 ( .A(\UUT/branch_rega [0]), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N191 ) );
  AND2_X1 U5302 ( .A1(\UUT/Mpath/out_regA[18] ), .A2(\UUT/Mpath/out_regB[18] ), 
        .ZN(\UUT/Mpath/the_alu/N107 ) );
  OR2_X1 U5303 ( .A1(\UUT/Mpath/out_regA[18] ), .A2(\UUT/Mpath/out_regB[18] ), 
        .ZN(\UUT/Mpath/the_alu/N139 ) );
  AND2_X2 U5304 ( .A1(\localbus/N50 ), .A2(\UUT/N3 ), .ZN(n6347) );
  INV_X1 U5305 ( .A(\localbus/c1_op[MASTER] ), .ZN(\localbus/N50 ) );
  AND2_X1 U5306 ( .A1(\UUT/Mpath/out_regA[15] ), .A2(\UUT/Mpath/out_regB[15] ), 
        .ZN(\UUT/Mpath/the_alu/N110 ) );
  OR2_X1 U5307 ( .A1(\UUT/Mpath/out_regA[15] ), .A2(\UUT/Mpath/out_regB[15] ), 
        .ZN(\UUT/Mpath/the_alu/N142 ) );
  AND2_X1 U5308 ( .A1(\UUT/Mpath/out_regA[19] ), .A2(\UUT/Mpath/out_regB[19] ), 
        .ZN(\UUT/Mpath/the_alu/N106 ) );
  OR2_X1 U5309 ( .A1(\UUT/Mpath/out_regA[19] ), .A2(\UUT/Mpath/out_regB[19] ), 
        .ZN(\UUT/Mpath/the_alu/N138 ) );
  AND2_X1 U5310 ( .A1(\UUT/Mpath/out_regA[20] ), .A2(\UUT/Mpath/out_regB[20] ), 
        .ZN(\UUT/Mpath/the_alu/N105 ) );
  OR2_X1 U5311 ( .A1(\UUT/Mpath/out_regA[20] ), .A2(\UUT/Mpath/out_regB[20] ), 
        .ZN(\UUT/Mpath/the_alu/N137 ) );
  AND2_X1 U5312 ( .A1(\UUT/Mpath/out_regA[21] ), .A2(\UUT/Mpath/out_regB[21] ), 
        .ZN(\UUT/Mpath/the_alu/N104 ) );
  OR2_X1 U5313 ( .A1(\UUT/Mpath/out_regA[21] ), .A2(\UUT/Mpath/out_regB[21] ), 
        .ZN(\UUT/Mpath/the_alu/N136 ) );
  AND2_X1 U5314 ( .A1(\UUT/Mpath/out_regA[9] ), .A2(\UUT/Mpath/out_regB[9] ), 
        .ZN(\UUT/Mpath/the_alu/N116 ) );
  OR2_X1 U5315 ( .A1(\UUT/Mpath/out_regA[9] ), .A2(\UUT/Mpath/out_regB[9] ), 
        .ZN(\UUT/Mpath/the_alu/N148 ) );
  AND2_X1 U5316 ( .A1(\UUT/Mpath/out_regA[10] ), .A2(\UUT/Mpath/out_regB[10] ), 
        .ZN(\UUT/Mpath/the_alu/N115 ) );
  OR2_X1 U5317 ( .A1(\UUT/Mpath/out_regA[10] ), .A2(\UUT/Mpath/out_regB[10] ), 
        .ZN(\UUT/Mpath/the_alu/N147 ) );
  AND2_X1 U5318 ( .A1(\UUT/Mpath/out_regA[22] ), .A2(\UUT/Mpath/out_regB[22] ), 
        .ZN(\UUT/Mpath/the_alu/N103 ) );
  OR2_X1 U5319 ( .A1(\UUT/Mpath/out_regA[22] ), .A2(\UUT/Mpath/out_regB[22] ), 
        .ZN(\UUT/Mpath/the_alu/N135 ) );
  BUF_X2 U5320 ( .A(n5529), .Z(n6364) );
  OAI21_X1 U5321 ( .B1(\UUT/regfile/N262 ), .B2(n2592), .A(n2593), .ZN(n5529)
         );
  AND3_X2 U5322 ( .A1(n1183), .A2(net54895), .A3(n5413), .ZN(n135) );
  AND2_X1 U5323 ( .A1(\UUT/Mpath/out_regA[23] ), .A2(\UUT/Mpath/out_regB[23] ), 
        .ZN(\UUT/Mpath/the_alu/N102 ) );
  OR2_X1 U5324 ( .A1(\UUT/Mpath/out_regA[23] ), .A2(\UUT/Mpath/out_regB[23] ), 
        .ZN(\UUT/Mpath/the_alu/N134 ) );
  AND2_X2 U5325 ( .A1(\UUT/Mpath/the_alu/N474 ), .A2(n2574), .ZN(n1215) );
  AND2_X2 U5326 ( .A1(n6348), .A2(\UUT/Mpath/the_alu/N492 ), .ZN(n1213) );
  AND2_X1 U5327 ( .A1(\UUT/Mpath/out_regA[8] ), .A2(\UUT/Mpath/out_regB[8] ), 
        .ZN(\UUT/Mpath/the_alu/N117 ) );
  OR2_X1 U5328 ( .A1(\UUT/Mpath/out_regA[8] ), .A2(\UUT/Mpath/out_regB[8] ), 
        .ZN(\UUT/Mpath/the_alu/N149 ) );
  AND2_X1 U5329 ( .A1(\UUT/Mpath/out_regA[16] ), .A2(\UUT/Mpath/out_regB[16] ), 
        .ZN(\UUT/Mpath/the_alu/N109 ) );
  OR2_X1 U5330 ( .A1(\UUT/Mpath/out_regA[16] ), .A2(\UUT/Mpath/out_regB[16] ), 
        .ZN(\UUT/Mpath/the_alu/N141 ) );
  AND2_X1 U5331 ( .A1(\UUT/Mpath/out_regA[17] ), .A2(\UUT/Mpath/out_regB[17] ), 
        .ZN(\UUT/Mpath/the_alu/N108 ) );
  OR2_X1 U5332 ( .A1(\UUT/Mpath/out_regA[17] ), .A2(\UUT/Mpath/out_regB[17] ), 
        .ZN(\UUT/Mpath/the_alu/N140 ) );
  AND2_X1 U5333 ( .A1(\UUT/Mpath/out_regA[28] ), .A2(\UUT/Mpath/out_regB[28] ), 
        .ZN(\UUT/Mpath/the_alu/N97 ) );
  OR2_X1 U5334 ( .A1(\UUT/Mpath/out_regA[28] ), .A2(\UUT/Mpath/out_regB[28] ), 
        .ZN(\UUT/Mpath/the_alu/N129 ) );
  AND2_X1 U5335 ( .A1(\UUT/Mpath/out_regA[27] ), .A2(\UUT/Mpath/out_regB[27] ), 
        .ZN(\UUT/Mpath/the_alu/N98 ) );
  OR2_X1 U5336 ( .A1(\UUT/Mpath/out_regA[27] ), .A2(\UUT/Mpath/out_regB[27] ), 
        .ZN(\UUT/Mpath/the_alu/N130 ) );
  AND2_X1 U5337 ( .A1(\UUT/Mpath/out_regA[25] ), .A2(\UUT/Mpath/out_regB[25] ), 
        .ZN(\UUT/Mpath/the_alu/N100 ) );
  OR2_X1 U5338 ( .A1(\UUT/Mpath/out_regA[25] ), .A2(\UUT/Mpath/out_regB[25] ), 
        .ZN(\UUT/Mpath/the_alu/N132 ) );
  AND2_X1 U5339 ( .A1(\UUT/Mpath/out_regA[30] ), .A2(\UUT/Mpath/out_regB[30] ), 
        .ZN(\UUT/Mpath/the_alu/N95 ) );
  OR2_X1 U5340 ( .A1(\UUT/Mpath/out_regA[30] ), .A2(\UUT/Mpath/out_regB[30] ), 
        .ZN(\UUT/Mpath/the_alu/N127 ) );
  OR2_X2 U5341 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/regfile/N269 ), .ZN(n132) );
  AND3_X2 U5342 ( .A1(n976), .A2(net54895), .A3(n5413), .ZN(n142) );
  AND2_X2 U5343 ( .A1(n6016), .A2(n6025), .ZN(n1291) );
  AND2_X4 U5344 ( .A1(n6312), .A2(n6321), .ZN(n1937) );
  BUF_X2 U5345 ( .A(n1214), .Z(n6365) );
  NOR3_X1 U5346 ( .A1(\UUT/Mpath/the_alu/N486 ), .A2(n6349), .A3(n2577), .ZN(
        n1214) );
  AND2_X1 U5347 ( .A1(\UUT/Mpath/out_regA[7] ), .A2(\UUT/Mpath/out_regB[7] ), 
        .ZN(\UUT/Mpath/the_alu/N118 ) );
  OR2_X1 U5348 ( .A1(\UUT/Mpath/out_regA[7] ), .A2(\UUT/Mpath/out_regB[7] ), 
        .ZN(\UUT/Mpath/the_alu/N150 ) );
  INV_X4 U5349 ( .A(n5553), .ZN(n1938) );
  INV_X2 U5350 ( .A(n5738), .ZN(n1294) );
  AND2_X1 U5351 ( .A1(\UUT/Mpath/out_regA[14] ), .A2(\UUT/Mpath/out_regB[14] ), 
        .ZN(\UUT/Mpath/the_alu/N111 ) );
  OR2_X1 U5352 ( .A1(\UUT/Mpath/out_regA[14] ), .A2(\UUT/Mpath/out_regB[14] ), 
        .ZN(\UUT/Mpath/the_alu/N143 ) );
  OR2_X1 U5353 ( .A1(\UUT/Mpath/out_regA[13] ), .A2(\UUT/Mpath/out_regB[13] ), 
        .ZN(\UUT/Mpath/the_alu/N144 ) );
  AND2_X1 U5354 ( .A1(\UUT/Mpath/out_regA[13] ), .A2(\UUT/Mpath/out_regB[13] ), 
        .ZN(\UUT/Mpath/the_alu/N112 ) );
  AND2_X1 U5355 ( .A1(\UUT/Mpath/out_regA[11] ), .A2(\UUT/Mpath/out_regB[11] ), 
        .ZN(\UUT/Mpath/the_alu/N114 ) );
  OR2_X1 U5356 ( .A1(\UUT/Mpath/out_regA[11] ), .A2(\UUT/Mpath/out_regB[11] ), 
        .ZN(\UUT/Mpath/the_alu/N146 ) );
  AND2_X4 U5357 ( .A1(n6305), .A2(n6308), .ZN(n5540) );
  AND2_X4 U5358 ( .A1(n6301), .A2(n6302), .ZN(n5535) );
  AND2_X2 U5359 ( .A1(n6009), .A2(n6012), .ZN(n5725) );
  AND2_X2 U5360 ( .A1(n6005), .A2(n6006), .ZN(n5720) );
  AND2_X2 U5361 ( .A1(\UUT/Mpath/the_shift/N108 ), .A2(n6324), .ZN(n6199) );
  INV_X1 U5362 ( .A(n5545), .ZN(n6366) );
  INV_X1 U5363 ( .A(n6366), .ZN(n6367) );
  INV_X1 U5364 ( .A(n6366), .ZN(n6368) );
  AND3_X2 U5365 ( .A1(\UUT/rs2_addr [4]), .A2(n6007), .A3(n6016), .ZN(n5730)
         );
  AND3_X4 U5366 ( .A1(n6318), .A2(n6310), .A3(n6308), .ZN(n5557) );
  NAND3_X1 U5367 ( .A1(\UUT/rs1_addr [3]), .A2(\UUT/rs1_addr [4]), .A3(n6308), 
        .ZN(n6369) );
  INV_X1 U5368 ( .A(n6369), .ZN(n6370) );
  INV_X1 U5369 ( .A(n6369), .ZN(n6371) );
  AND3_X2 U5370 ( .A1(n6022), .A2(n6014), .A3(n6012), .ZN(n5742) );
  AND3_X4 U5371 ( .A1(n6308), .A2(n2591), .A3(n6310), .ZN(n1930) );
  AND2_X2 U5372 ( .A1(n6309), .A2(n6303), .ZN(n6308) );
  AND3_X2 U5373 ( .A1(\UUT/rs2_addr [3]), .A2(\UUT/rs2_addr [4]), .A3(n6012), 
        .ZN(n5735) );
  AND2_X1 U5374 ( .A1(\UUT/Mpath/out_regA[12] ), .A2(\UUT/Mpath/out_regB[12] ), 
        .ZN(\UUT/Mpath/the_alu/N113 ) );
  OR2_X1 U5375 ( .A1(\UUT/Mpath/out_regA[12] ), .A2(\UUT/Mpath/out_regB[12] ), 
        .ZN(\UUT/Mpath/the_alu/N145 ) );
  AND3_X2 U5376 ( .A1(n6010), .A2(n6008), .A3(n6021), .ZN(n1282) );
  INV_X2 U5377 ( .A(n5722), .ZN(n1277) );
  NAND2_X2 U5378 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(\UUT/byp_controlB[0] ), 
        .ZN(n5434) );
  NAND3_X2 U5379 ( .A1(\UUT/Mpath/the_mult/N285 ), .A2(n975), .A3(
        \UUT/Mpath/the_mult/N313 ), .ZN(n133) );
  INV_X4 U5380 ( .A(n5537), .ZN(n1926) );
  NAND2_X4 U5381 ( .A1(n6319), .A2(n6316), .ZN(n5558) );
  AND3_X2 U5382 ( .A1(\UUT/Mpath/the_mult/N198 ), .A2(n1194), .A3(
        \UUT/Mpath/the_mult/N216 ), .ZN(n291) );
  AND2_X1 U5383 ( .A1(\UUT/Mpath/out_regA[29] ), .A2(\UUT/Mpath/out_regB[29] ), 
        .ZN(\UUT/Mpath/the_alu/N96 ) );
  OR2_X1 U5384 ( .A1(\UUT/Mpath/out_regA[29] ), .A2(\UUT/Mpath/out_regB[29] ), 
        .ZN(\UUT/Mpath/the_alu/N128 ) );
  NAND2_X2 U5385 ( .A1(n6023), .A2(n6020), .ZN(n5743) );
  OR2_X1 U5386 ( .A1(\UUT/Mpath/out_regA[5] ), .A2(\UUT/Mpath/out_regB[5] ), 
        .ZN(\UUT/Mpath/the_alu/N152 ) );
  AND2_X1 U5387 ( .A1(\UUT/Mpath/out_regA[5] ), .A2(\UUT/Mpath/out_regB[5] ), 
        .ZN(\UUT/Mpath/the_alu/N120 ) );
  AND2_X1 U5388 ( .A1(\UUT/Mpath/out_regA[26] ), .A2(\UUT/Mpath/out_regB[26] ), 
        .ZN(\UUT/Mpath/the_alu/N99 ) );
  OR2_X1 U5389 ( .A1(\UUT/Mpath/out_regA[26] ), .A2(\UUT/Mpath/out_regB[26] ), 
        .ZN(\UUT/Mpath/the_alu/N131 ) );
  AND3_X2 U5390 ( .A1(n6309), .A2(n2591), .A3(n6321), .ZN(n1931) );
  AND3_X2 U5391 ( .A1(n6012), .A2(n1912), .A3(n6014), .ZN(n1284) );
  NAND2_X2 U5392 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/Mcontrol/st_logic/N42 ), .ZN(n129) );
  NAND2_X2 U5393 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(
        \UUT/Mcontrol/st_logic/N42 ), .ZN(n5430) );
  AND4_X2 U5394 ( .A1(net54895), .A2(n971), .A3(n5413), .A4(n972), .ZN(n145)
         );
  OR2_X2 U5395 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(\UUT/regfile/N269 ), .ZN(
        n5432) );
  INV_X1 U5396 ( .A(\UUT/BYP_BRANCH_MUXB/N39 ), .ZN(\UUT/BYP_BRANCH_MUXB/N4 )
         );
  INV_X2 U5397 ( .A(n620), .ZN(n611) );
  INV_X2 U5398 ( .A(n585), .ZN(n576) );
  INV_X2 U5399 ( .A(n560), .ZN(n551) );
  INV_X2 U5400 ( .A(n657), .ZN(n648) );
  INV_X2 U5401 ( .A(n680), .ZN(n671) );
  INV_X2 U5402 ( .A(n534), .ZN(n525) );
  INV_X2 U5403 ( .A(n509), .ZN(n500) );
  INV_X2 U5404 ( .A(n708), .ZN(n699) );
  INV_X2 U5405 ( .A(n731), .ZN(n722) );
  INV_X2 U5406 ( .A(n480), .ZN(n471) );
  INV_X2 U5407 ( .A(n459), .ZN(n447) );
  INV_X2 U5408 ( .A(n754), .ZN(n745) );
  INV_X2 U5409 ( .A(n777), .ZN(n768) );
  INV_X2 U5410 ( .A(n432), .ZN(n423) );
  INV_X2 U5411 ( .A(n410), .ZN(n401) );
  INV_X2 U5412 ( .A(n800), .ZN(n802) );
  INV_X2 U5413 ( .A(n812), .ZN(n814) );
  INV_X2 U5414 ( .A(n388), .ZN(n379) );
  INV_X2 U5415 ( .A(n362), .ZN(n353) );
  INV_X2 U5416 ( .A(n641), .ZN(n958) );
  INV_X2 U5417 ( .A(n605), .ZN(n959) );
  INV_X2 U5418 ( .A(n341), .ZN(n332) );
  INV_X2 U5419 ( .A(n315), .ZN(n303) );
  INV_X2 U5420 ( .A(n1076), .ZN(n960) );
  NAND2_X2 U5421 ( .A1(n6023), .A2(n6018), .ZN(n5745) );
  NAND2_X4 U5422 ( .A1(n6319), .A2(n6314), .ZN(n5560) );
  INV_X4 U5423 ( .A(n5542), .ZN(n1927) );
  INV_X2 U5424 ( .A(n5727), .ZN(n1279) );
  NAND3_X2 U5425 ( .A1(n6007), .A2(n6008), .A3(n6005), .ZN(n5717) );
  NAND3_X4 U5426 ( .A1(n6303), .A2(n6304), .A3(n6301), .ZN(n5532) );
  NAND3_X2 U5427 ( .A1(n6020), .A2(\UUT/rs2_addr [4]), .A3(n6006), .ZN(n5732)
         );
  AND2_X1 U5428 ( .A1(\UUT/Mpath/out_regA[24] ), .A2(\UUT/Mpath/out_regB[24] ), 
        .ZN(\UUT/Mpath/the_alu/N101 ) );
  OR2_X1 U5429 ( .A1(\UUT/Mpath/out_regA[24] ), .A2(\UUT/Mpath/out_regB[24] ), 
        .ZN(\UUT/Mpath/the_alu/N133 ) );
  NAND3_X2 U5430 ( .A1(n6018), .A2(\UUT/rs2_addr [1]), .A3(n6025), .ZN(n5746)
         );
  NAND3_X4 U5431 ( .A1(n6316), .A2(\UUT/rs1_addr [4]), .A3(n6302), .ZN(n5547)
         );
  NOR2_X2 U5432 ( .A1(n6304), .A2(\UUT/rs1_addr [0]), .ZN(n6302) );
  NAND3_X2 U5433 ( .A1(n6314), .A2(\UUT/rs1_addr [1]), .A3(n6321), .ZN(n5561)
         );
  NAND3_X2 U5434 ( .A1(n6313), .A2(n6316), .A3(\UUT/rs1_addr [1]), .ZN(n5546)
         );
  NAND3_X2 U5435 ( .A1(n6017), .A2(n6020), .A3(\UUT/rs2_addr [1]), .ZN(n5731)
         );
  BUF_X1 U5436 ( .A(\UUT/Mcontrol/Nextpc_decoding/N255 ), .Z(n6372) );
  NAND3_X4 U5437 ( .A1(n6303), .A2(n6310), .A3(n6312), .ZN(n1934) );
  OR2_X1 U5438 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N114 ) );
  OR2_X1 U5439 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N262 ) );
  OR2_X1 U5440 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N122 ) );
  OR2_X1 U5441 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N250 ) );
  OR2_X1 U5442 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N256 ) );
  OR2_X1 U5443 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N238 ) );
  OR2_X1 U5444 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N226 ) );
  OR2_X1 U5445 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N232 ) );
  OR2_X1 U5446 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N244 ) );
  OR2_X1 U5447 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N60 ) );
  OR2_X1 U5448 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N67 ) );
  OR2_X1 U5449 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N105 ) );
  OR2_X1 U5450 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N98 ) );
  OR2_X1 U5451 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N92 ) );
  OR2_X1 U5452 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N85 ) );
  OR2_X1 U5453 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N73 ) );
  OR2_X1 U5454 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(n6372), .ZN(
        \UUT/Mcontrol/st_logic/N79 ) );
  AND2_X1 U5455 ( .A1(\UUT/Mpath/out_regA[6] ), .A2(\UUT/Mpath/out_regB[6] ), 
        .ZN(\UUT/Mpath/the_alu/N119 ) );
  OR2_X1 U5456 ( .A1(\UUT/Mpath/out_regA[6] ), .A2(\UUT/Mpath/out_regB[6] ), 
        .ZN(\UUT/Mpath/the_alu/N151 ) );
  NAND3_X2 U5457 ( .A1(n6007), .A2(n6014), .A3(n6016), .ZN(n1287) );
  INV_X2 U5458 ( .A(n5739), .ZN(n1290) );
  INV_X4 U5459 ( .A(\localbus/N226 ), .ZN(n6346) );
  INV_X2 U5460 ( .A(n5721), .ZN(n1275) );
  INV_X4 U5461 ( .A(n5554), .ZN(n1936) );
  NAND2_X2 U5462 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/byp_controlB[0] ), 
        .ZN(n131) );
  INV_X4 U5463 ( .A(n5536), .ZN(n1925) );
  NAND3_X1 U5464 ( .A1(n6306), .A2(n6304), .A3(n6317), .ZN(n6373) );
  INV_X2 U5465 ( .A(\UUT/rs1_addr [2]), .ZN(n6306) );
  NAND3_X2 U5466 ( .A1(n6013), .A2(n1912), .A3(n6025), .ZN(n1288) );
  NAND2_X1 U5467 ( .A1(n6317), .A2(n6309), .ZN(n6374) );
  INV_X1 U5468 ( .A(n6374), .ZN(n6375) );
  INV_X1 U5469 ( .A(n6374), .ZN(n6376) );
  AND2_X2 U5470 ( .A1(n6021), .A2(n6013), .ZN(n5741) );
  AND2_X4 U5471 ( .A1(n6312), .A2(n6313), .ZN(n5544) );
  AND2_X2 U5472 ( .A1(n975), .A2(n973), .ZN(n144) );
  NAND3_X2 U5473 ( .A1(\UUT/rs2_addr [1]), .A2(n6010), .A3(n6021), .ZN(n5737)
         );
  AND2_X2 U5474 ( .A1(n6016), .A2(n6017), .ZN(n5729) );
  NAND3_X2 U5475 ( .A1(\UUT/rs2_addr [1]), .A2(n6020), .A3(n6025), .ZN(n5744)
         );
  NAND3_X2 U5476 ( .A1(\UUT/rs1_addr [1]), .A2(n6306), .A3(n6317), .ZN(n5552)
         );
  AND3_X4 U5477 ( .A1(n6313), .A2(\UUT/rs1_addr [3]), .A3(n6309), .ZN(n5549)
         );
  NAND3_X2 U5478 ( .A1(\UUT/rs1_addr [1]), .A2(n6316), .A3(n6321), .ZN(n5559)
         );
  AND3_X2 U5479 ( .A1(n6013), .A2(\UUT/rs2_addr [0]), .A3(n6009), .ZN(n5724)
         );
  AND3_X2 U5480 ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/rs2_addr [0]), .A3(n6005), 
        .ZN(n5719) );
  AND3_X2 U5481 ( .A1(n6017), .A2(\UUT/rs2_addr [3]), .A3(n6013), .ZN(n5734)
         );
  AND3_X2 U5482 ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/rs1_addr [0]), .A3(n6301), 
        .ZN(n5534) );
  NAND3_X2 U5483 ( .A1(\UUT/rs2_addr [0]), .A2(n6008), .A3(n6005), .ZN(n5716)
         );
  AND3_X4 U5484 ( .A1(n6309), .A2(\UUT/rs1_addr [0]), .A3(n6305), .ZN(n5539)
         );
  NAND3_X2 U5485 ( .A1(\UUT/Mpath/the_mult/N255 ), .A2(n975), .A3(
        \UUT/Mpath/the_mult/N311 ), .ZN(n140) );
  NAND3_X4 U5486 ( .A1(\UUT/rs1_addr [0]), .A2(n6304), .A3(n6301), .ZN(n5531)
         );
  NAND3_X2 U5487 ( .A1(n6010), .A2(n6022), .A3(n6023), .ZN(n5736) );
  NAND3_X4 U5488 ( .A1(n6306), .A2(n6318), .A3(n6319), .ZN(n5551) );
  NAND3_X2 U5489 ( .A1(\UUT/rs1_addr [1]), .A2(n6313), .A3(n6314), .ZN(n5541)
         );
  NAND3_X2 U5490 ( .A1(\UUT/rs2_addr [1]), .A2(n6017), .A3(n6018), .ZN(n5726)
         );
  INV_X2 U5491 ( .A(n831), .ZN(n181) );
  OAI221_X4 U5492 ( .B1(n5873), .B2(n281), .C1(n5710), .C2(n5473), .A(n282), 
        .ZN(n831) );
  INV_X2 U5493 ( .A(n849), .ZN(n130) );
  OAI221_X4 U5494 ( .B1(n5851), .B2(n281), .C1(n5710), .C2(n5464), .A(n282), 
        .ZN(n849) );
  INV_X2 U5495 ( .A(n825), .ZN(n194) );
  OAI221_X4 U5496 ( .B1(n5882), .B2(n281), .C1(n5710), .C2(n5476), .A(n282), 
        .ZN(n825) );
  INV_X2 U5497 ( .A(n843), .ZN(n153) );
  OAI221_X4 U5498 ( .B1(n5857), .B2(n281), .C1(n5710), .C2(n5467), .A(n282), 
        .ZN(n843) );
  INV_X2 U5499 ( .A(n1171), .ZN(n952) );
  OAI221_X4 U5500 ( .B1(n5825), .B2(n281), .C1(n5710), .C2(n5455), .A(n282), 
        .ZN(n1171) );
  INV_X2 U5501 ( .A(n280), .ZN(n209) );
  OAI221_X4 U5502 ( .B1(n5890), .B2(n281), .C1(n5710), .C2(n5479), .A(n282), 
        .ZN(n280) );
  INV_X2 U5503 ( .A(n837), .ZN(n165) );
  OAI221_X4 U5504 ( .B1(n5863), .B2(n281), .C1(n5710), .C2(n5470), .A(n282), 
        .ZN(n837) );
  INV_X2 U5505 ( .A(n869), .ZN(n860) );
  OAI221_X4 U5506 ( .B1(n5832), .B2(n281), .C1(n5710), .C2(n5458), .A(n282), 
        .ZN(n869) );
  INV_X2 U5507 ( .A(n83), .ZN(n82) );
  NOR2_X4 U5508 ( .A1(net54903), .A2(n5530), .ZN(n319) );
  NAND2_X2 U5509 ( .A1(n116), .A2(net54859), .ZN(n83) );
  NOR2_X4 U5510 ( .A1(net54903), .A2(n6364), .ZN(n318) );
  NOR2_X4 U5511 ( .A1(n6409), .A2(n5530), .ZN(n314) );
  NOR2_X4 U5512 ( .A1(n6284), .A2(\UUT/Mpath/N119 ), .ZN(n5612) );
  NOR2_X4 U5513 ( .A1(n6409), .A2(n6364), .ZN(n312) );
  NOR3_X4 U5514 ( .A1(n285), .A2(\UUT/Mpath/N128 ), .A3(n1195), .ZN(n325) );
  OR2_X1 U5515 ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N127 ), .ZN(
        \UUT/Mpath/N128 ) );
  INV_X2 U5516 ( .A(n6674), .ZN(n6675) );
  NOR2_X4 U5517 ( .A1(n2573), .A2(\UUT/Mpath/the_alu/N474 ), .ZN(n1208) );
  NOR2_X4 U5518 ( .A1(n1193), .A2(\UUT/Mpath/the_mult/N216 ), .ZN(n284) );
  OR2_X1 U5519 ( .A1(\UUT/Mpath/the_mult/x_mul_command[0] ), .A2(
        \UUT/Mpath/the_mult/N215 ), .ZN(\UUT/Mpath/the_mult/N216 ) );
  NOR2_X4 U5520 ( .A1(n1211), .A2(n2572), .ZN(n1210) );
  NOR2_X4 U5521 ( .A1(n6325), .A2(\UUT/Mpath/the_shift/N118 ), .ZN(n6198) );
  NOR2_X4 U5522 ( .A1(n6323), .A2(\UUT/Mpath/the_shift/N108 ), .ZN(n6200) );
  NOR2_X4 U5523 ( .A1(n2576), .A2(n6349), .ZN(n1212) );
  NAND2_X4 U5524 ( .A1(\UUT/byp_controlA[2] ), .A2(\UUT/Mcontrol/st_logic/N47 ), .ZN(n5528) );
  NOR2_X4 U5525 ( .A1(n6003), .A2(\localbus/c2_op[MASTER] ), .ZN(n5779) );
  BUF_X2 U5526 ( .A(n5780), .Z(n6377) );
  AND2_X1 U5527 ( .A1(\localbus/N335 ), .A2(\localbus/N337 ), .ZN(
        \localbus/N93 ) );
  NAND2_X4 U5528 ( .A1(\UUT/byp_controlA[2] ), .A2(\UUT/byp_controlA[0] ), 
        .ZN(n5530) );
  BUF_X2 U5529 ( .A(n6201), .Z(n6378) );
  BUF_X2 U5530 ( .A(n290), .Z(n6379) );
  INV_X2 U5531 ( .A(n249), .ZN(n6380) );
  INV_X2 U5532 ( .A(n248), .ZN(n249) );
  NOR2_X4 U5533 ( .A1(\UUT/exe_outsel [0]), .A2(\UUT/Mpath/N121 ), .ZN(n285)
         );
  OR2_X1 U5534 ( .A1(\UUT/Mpath/N116 ), .A2(\UUT/exe_outsel [2]), .ZN(
        \UUT/Mpath/N121 ) );
  INV_X2 U5535 ( .A(n253), .ZN(n6381) );
  INV_X2 U5536 ( .A(n247), .ZN(n6382) );
  INV_X2 U5537 ( .A(n245), .ZN(n6383) );
  INV_X2 U5538 ( .A(n251), .ZN(n6384) );
  INV_X2 U5539 ( .A(n252), .ZN(n253) );
  INV_X2 U5540 ( .A(n246), .ZN(n247) );
  INV_X2 U5541 ( .A(n244), .ZN(n245) );
  INV_X2 U5542 ( .A(n250), .ZN(n251) );
  INV_X2 U5543 ( .A(n243), .ZN(n6385) );
  INV_X2 U5544 ( .A(n257), .ZN(n6386) );
  INV_X2 U5545 ( .A(n255), .ZN(n6387) );
  INV_X2 U5546 ( .A(n241), .ZN(n6388) );
  INV_X2 U5547 ( .A(n242), .ZN(n243) );
  INV_X2 U5548 ( .A(n256), .ZN(n257) );
  INV_X2 U5549 ( .A(n254), .ZN(n255) );
  INV_X2 U5550 ( .A(n240), .ZN(n241) );
  INV_X2 U5551 ( .A(n263), .ZN(n6389) );
  INV_X2 U5552 ( .A(n239), .ZN(n6390) );
  INV_X2 U5553 ( .A(n237), .ZN(n6391) );
  INV_X2 U5554 ( .A(n259), .ZN(n6392) );
  INV_X2 U5555 ( .A(n262), .ZN(n263) );
  INV_X2 U5556 ( .A(n238), .ZN(n239) );
  INV_X2 U5557 ( .A(n236), .ZN(n237) );
  INV_X2 U5558 ( .A(n258), .ZN(n259) );
  INV_X2 U5559 ( .A(n235), .ZN(n6393) );
  INV_X2 U5560 ( .A(n261), .ZN(n6394) );
  INV_X2 U5561 ( .A(n265), .ZN(n6395) );
  INV_X2 U5562 ( .A(n233), .ZN(n6396) );
  INV_X2 U5563 ( .A(n234), .ZN(n235) );
  INV_X2 U5564 ( .A(n260), .ZN(n261) );
  INV_X2 U5565 ( .A(n264), .ZN(n265) );
  INV_X2 U5566 ( .A(n232), .ZN(n233) );
  INV_X2 U5567 ( .A(n271), .ZN(n6397) );
  INV_X2 U5568 ( .A(n231), .ZN(n6398) );
  INV_X2 U5569 ( .A(n227), .ZN(n6399) );
  INV_X2 U5570 ( .A(n267), .ZN(n6400) );
  INV_X2 U5571 ( .A(n270), .ZN(n271) );
  INV_X2 U5572 ( .A(n230), .ZN(n231) );
  INV_X2 U5573 ( .A(n226), .ZN(n227) );
  INV_X2 U5574 ( .A(n266), .ZN(n267) );
  INV_X2 U5575 ( .A(n223), .ZN(n6401) );
  INV_X2 U5576 ( .A(n269), .ZN(n6402) );
  INV_X2 U5577 ( .A(n273), .ZN(n6403) );
  INV_X2 U5578 ( .A(n229), .ZN(n6404) );
  INV_X2 U5579 ( .A(n222), .ZN(n223) );
  INV_X2 U5580 ( .A(n268), .ZN(n269) );
  INV_X2 U5581 ( .A(n272), .ZN(n273) );
  INV_X2 U5582 ( .A(n228), .ZN(n229) );
  INV_X2 U5583 ( .A(n277), .ZN(n6405) );
  INV_X2 U5584 ( .A(n225), .ZN(n6406) );
  INV_X2 U5585 ( .A(n219), .ZN(n6407) );
  INV_X2 U5586 ( .A(n275), .ZN(n6408) );
  INV_X2 U5587 ( .A(n276), .ZN(n277) );
  INV_X2 U5588 ( .A(n224), .ZN(n225) );
  INV_X2 U5589 ( .A(n218), .ZN(n219) );
  INV_X2 U5590 ( .A(n274), .ZN(n275) );
  BUF_X4 U5591 ( .A(n73), .Z(n6409) );
  INV_X2 U5592 ( .A(n221), .ZN(n6410) );
  INV_X2 U5593 ( .A(n279), .ZN(n6411) );
  INV_X2 U5594 ( .A(n6409), .ZN(n147) );
  NOR2_X4 U5595 ( .A1(\UUT/Mpath/N115 ), .A2(\UUT/Mpath/N119 ), .ZN(n5564) );
  INV_X2 U5596 ( .A(n220), .ZN(n221) );
  INV_X2 U5597 ( .A(n278), .ZN(n279) );
  INV_X1 U5598 ( .A(\UUT/jar_in [7]), .ZN(n6650) );
  INV_X1 U5599 ( .A(\UUT/jar_in [3]), .ZN(n6648) );
  INV_X1 U5600 ( .A(\UUT/jar_in [6]), .ZN(n6655) );
  NAND2_X1 U5601 ( .A1(n6466), .A2(n6467), .ZN(n6412) );
  NAND2_X1 U5602 ( .A1(n136), .A2(n6413), .ZN(n2895) );
  INV_X1 U5603 ( .A(n6412), .ZN(n6413) );
  AOI21_X1 U5604 ( .B1(n139), .B2(\UUT/Mpath/the_mult/Mad_out [61]), .A(n6428), 
        .ZN(n136) );
  OR2_X1 U5605 ( .A1(n133), .A2(n134), .ZN(n6466) );
  OR2_X1 U5606 ( .A1(n133), .A2(n154), .ZN(n6414) );
  OR2_X1 U5607 ( .A1(n5689), .A2(n135), .ZN(n6415) );
  NAND3_X1 U5608 ( .A1(n6414), .A2(n6415), .A3(n155), .ZN(n2901) );
  AND2_X1 U5609 ( .A1(n6457), .A2(n6458), .ZN(n155) );
  OR2_X1 U5610 ( .A1(n294), .A2(n466), .ZN(n6416) );
  OR2_X1 U5611 ( .A1(n295), .A2(n2660), .ZN(n6417) );
  NAND3_X1 U5612 ( .A1(n6416), .A2(n6417), .A3(n468), .ZN(n3243) );
  AND3_X1 U5613 ( .A1(n6616), .A2(n6617), .A3(n6618), .ZN(n468) );
  AOI22_X2 U5614 ( .A1(n908), .A2(\UUT/break_code[2] ), .B1(n6449), .B2(
        \UUT/Mcontrol/Nextpc_decoding/Bta [2]), .ZN(n2327) );
  OR2_X1 U5615 ( .A1(n6634), .A2(n6475), .ZN(n6633) );
  OR2_X1 U5616 ( .A1(n787), .A2(n294), .ZN(n6418) );
  OR2_X1 U5617 ( .A1(n295), .A2(n2698), .ZN(n6419) );
  NAND3_X1 U5618 ( .A1(n6418), .A2(n6419), .A3(n790), .ZN(n3735) );
  AND3_X1 U5619 ( .A1(n6536), .A2(n6537), .A3(n6538), .ZN(n790) );
  AND3_X1 U5620 ( .A1(n6703), .A2(n6704), .A3(n2374), .ZN(n571) );
  OR2_X1 U5621 ( .A1(n6716), .A2(n6687), .ZN(n6420) );
  OR2_X1 U5622 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N125 ), .A2(n6688), .ZN(
        n6421) );
  NAND3_X1 U5623 ( .A1(n6420), .A2(n6421), .A3(n2351), .ZN(n6686) );
  INV_X1 U5624 ( .A(\UUT/jar_in [12]), .ZN(n6687) );
  INV_X1 U5625 ( .A(\UUT/branch_rega [12]), .ZN(n6688) );
  NAND2_X1 U5626 ( .A1(n6906), .A2(n6907), .ZN(n6422) );
  NAND3_X1 U5627 ( .A1(n6908), .A2(n6423), .A3(n6905), .ZN(n6909) );
  INV_X1 U5628 ( .A(n6422), .ZN(n6423) );
  NAND2_X1 U5629 ( .A1(\localbus/c1_addr_outbus[30] ), .A2(
        \localbus/c1_addr_outbus[29] ), .ZN(n6424) );
  INV_X1 U5630 ( .A(n6595), .ZN(n6425) );
  AND2_X1 U5631 ( .A1(n6424), .A2(n6425), .ZN(n6903) );
  AND2_X1 U5632 ( .A1(n6347), .A2(n6644), .ZN(n6595) );
  NOR2_X1 U5633 ( .A1(n6480), .A2(n6481), .ZN(n5456) );
  AND2_X1 U5634 ( .A1(n5563), .A2(n5564), .ZN(n6481) );
  BUF_X1 U5635 ( .A(n6128), .Z(n6446) );
  NAND4_X2 U5636 ( .A1(\UUT/Mcontrol/Operation_decoding32/N89 ), .A2(n6285), 
        .A3(n6045), .A4(\UUT/Mcontrol/Operation_decoding32/N1975 ), .ZN(n6128)
         );
  AND4_X1 U5637 ( .A1(n6447), .A2(n4359), .A3(n4357), .A4(n4358), .ZN(n6915)
         );
  NOR4_X1 U5638 ( .A1(\localbus/c1_addr_outbus[28] ), .A2(
        \localbus/c1_addr_outbus[27] ), .A3(n6595), .A4(
        \localbus/c1_addr_outbus[29] ), .ZN(n6447) );
  BUF_X1 U5639 ( .A(n6619), .Z(n6448) );
  NOR2_X1 U5640 ( .A1(n6639), .A2(n6702), .ZN(n6449) );
  NOR2_X1 U5641 ( .A1(n6639), .A2(n6702), .ZN(n6715) );
  BUF_X4 U5642 ( .A(\UUT/Mpath/out_regA[1] ), .Z(n6450) );
  NAND2_X1 U5643 ( .A1(n6468), .A2(n6469), .ZN(n6451) );
  BUF_X1 U5644 ( .A(\UUT/Mpath/out_regB[1] ), .Z(n6900) );
  BUF_X1 U5645 ( .A(n5578), .Z(n6452) );
  BUF_X1 U5646 ( .A(\UUT/Mpath/out_regB[0] ), .Z(n6453) );
  OR2_X1 U5647 ( .A1(n395), .A2(n294), .ZN(n6454) );
  OR2_X1 U5648 ( .A1(n295), .A2(n2651), .ZN(n6455) );
  NAND3_X1 U5649 ( .A1(n6454), .A2(n6455), .A3(n398), .ZN(n3123) );
  BUF_X2 U5650 ( .A(n6488), .Z(n6475) );
  AND2_X1 U5651 ( .A1(n2324), .A2(n295), .ZN(n297) );
  BUF_X1 U5652 ( .A(n2324), .Z(n6646) );
  AND2_X1 U5653 ( .A1(n2324), .A2(n295), .ZN(n6711) );
  BUF_X2 U5654 ( .A(n2324), .Z(n6503) );
  OR2_X1 U5655 ( .A1(n6693), .A2(n6456), .ZN(n6469) );
  NAND2_X1 U5656 ( .A1(n6614), .A2(\UUT/Mcontrol/Nextpc_decoding/Bta [9]), 
        .ZN(n6456) );
  NAND2_X4 U5657 ( .A1(n137), .A2(n156), .ZN(n6457) );
  NAND2_X1 U5658 ( .A1(\UUT/Mpath/the_mult/Mad_out [60]), .A2(n139), .ZN(n6458) );
  NAND2_X1 U5659 ( .A1(n6582), .A2(n6583), .ZN(n6459) );
  NAND2_X1 U5660 ( .A1(n905), .A2(n6460), .ZN(n4041) );
  INV_X1 U5661 ( .A(n6459), .ZN(n6460) );
  NAND2_X1 U5662 ( .A1(\UUT/Mpath/the_mult/Mad_out [63]), .A2(n139), .ZN(n6461) );
  NAND2_X1 U5663 ( .A1(n6461), .A2(net56414), .ZN(n4329) );
  OAI22_X2 U5664 ( .A1(n6633), .A2(n6292), .B1(n6293), .B2(
        \UUT/Mcontrol/Nextpc_decoding/N254 ), .ZN(n6641) );
  NAND2_X1 U5665 ( .A1(n6572), .A2(n6573), .ZN(n6462) );
  AND3_X1 U5666 ( .A1(n6512), .A2(n6513), .A3(n2536), .ZN(n6463) );
  OR2_X1 U5667 ( .A1(n6831), .A2(n6475), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N27 ) );
  AND2_X1 U5668 ( .A1(n6714), .A2(n295), .ZN(n299) );
  AND2_X1 U5669 ( .A1(n6714), .A2(n295), .ZN(n6511) );
  BUF_X1 U5670 ( .A(\UUT/branch_rega [21]), .Z(n6464) );
  AOI22_X1 U5671 ( .A1(n5570), .A2(\UUT/Mpath/N119 ), .B1(n5571), .B2(n5564), 
        .ZN(n5462) );
  OR2_X1 U5672 ( .A1(n6693), .A2(n6465), .ZN(n6573) );
  NAND2_X1 U5673 ( .A1(n6614), .A2(\UUT/Mcontrol/Nextpc_decoding/Bta [10]), 
        .ZN(n6465) );
  OR3_X4 U5674 ( .A1(\localbus/N57 ), .A2(n4340), .A3(n4339), .ZN(n6637) );
  OR2_X1 U5675 ( .A1(n5688), .A2(n135), .ZN(n6467) );
  OAI22_X1 U5676 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N27 ), .A2(n6292), .B1(
        n6293), .B2(\UUT/Mcontrol/Nextpc_decoding/N254 ), .ZN(n6289) );
  OAI222_X1 U5677 ( .A1(n6619), .A2(n5528), .B1(n5414), .B2(n6364), .C1(n5455), 
        .C2(n5530), .ZN(n6488) );
  AND2_X1 U5678 ( .A1(n6845), .A2(n6519), .ZN(n6872) );
  NOR3_X2 U5679 ( .A1(n6676), .A2(n6677), .A3(n6462), .ZN(n979) );
  NAND2_X4 U5680 ( .A1(n137), .A2(n138), .ZN(net87679) );
  NAND2_X1 U5681 ( .A1(n908), .A2(\UUT/break_code[9] ), .ZN(n6468) );
  OAI222_X4 U5682 ( .A1(n5430), .A2(n6448), .B1(n5454), .B2(n5432), .C1(n5455), 
        .C2(n5434), .ZN(\UUT/branch_regb [31]) );
  NAND2_X1 U5683 ( .A1(n1260), .A2(n1259), .ZN(n6470) );
  NAND2_X1 U5684 ( .A1(n1261), .A2(n6471), .ZN(n5563) );
  INV_X1 U5685 ( .A(n6470), .ZN(n6471) );
  AOI21_X1 U5686 ( .B1(n6641), .B2(n6290), .A(n6291), .ZN(n6472) );
  AOI21_X1 U5687 ( .B1(n6641), .B2(n6290), .A(n6291), .ZN(n6645) );
  NAND2_X1 U5688 ( .A1(\UUT/Mpath/the_mult/Mad_out [62]), .A2(n139), .ZN(n6473) );
  NAND2_X1 U5689 ( .A1(n6473), .A2(n6474), .ZN(n3977) );
  AND2_X1 U5690 ( .A1(n6483), .A2(n6694), .ZN(n6474) );
  NAND2_X1 U5691 ( .A1(n6711), .A2(\UUT/jar_in [20]), .ZN(n6476) );
  NAND2_X1 U5692 ( .A1(n298), .A2(\UUT/branch_rega [20]), .ZN(n6477) );
  NAND2_X1 U5693 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [20]), .A2(n299), 
        .ZN(n6478) );
  AND3_X2 U5694 ( .A1(n6476), .A2(n6477), .A3(n6478), .ZN(n350) );
  OAI22_X1 U5695 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6287), .B1(
        n6472), .B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6479) );
  AND2_X1 U5696 ( .A1(n5562), .A2(\UUT/Mpath/N119 ), .ZN(n6480) );
  OAI22_X1 U5697 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6287), .B1(
        n6645), .B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6710) );
  NAND2_X2 U5698 ( .A1(n6843), .A2(n6844), .ZN(n6482) );
  INV_X1 U5699 ( .A(n6482), .ZN(n6483) );
  AOI22_X2 U5700 ( .A1(n6197), .A2(\UUT/Mpath/N119 ), .B1(n6690), .B2(n5564), 
        .ZN(n6619) );
  OR2_X2 U5701 ( .A1(n6770), .A2(n6776), .ZN(n6769) );
  AOI222_X2 U5702 ( .A1(n6107), .A2(n5564), .B1(n346), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[21] ), .C2(n5612), .ZN(n5486) );
  AND2_X2 U5703 ( .A1(n6484), .A2(n6736), .ZN(n6581) );
  INV_X32 U5704 ( .A(n6621), .ZN(n6484) );
  NAND2_X2 U5705 ( .A1(n1255), .A2(n6561), .ZN(n5571) );
  AOI22_X1 U5706 ( .A1(n6197), .A2(\UUT/Mpath/N119 ), .B1(n6690), .B2(n5564), 
        .ZN(n6486) );
  AOI22_X1 U5707 ( .A1(n6197), .A2(\UUT/Mpath/N119 ), .B1(n6690), .B2(n5564), 
        .ZN(n6485) );
  NAND3_X1 U5708 ( .A1(n6703), .A2(n6704), .A3(n2374), .ZN(n6487) );
  OAI222_X1 U5709 ( .A1(n6486), .A2(n5528), .B1(n5414), .B2(n6364), .C1(n5455), 
        .C2(n5530), .ZN(n6489) );
  OAI222_X1 U5710 ( .A1(n6485), .A2(n5528), .B1(n5414), .B2(n6364), .C1(n5455), 
        .C2(n5530), .ZN(\UUT/branch_rega [31]) );
  INV_X1 U5711 ( .A(\UUT/Mcontrol/Operation_decoding32/N1945 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1946 ) );
  OR2_X4 U5712 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1944 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1945 ) );
  INV_X1 U5713 ( .A(n6649), .ZN(n643) );
  OAI221_X1 U5714 ( .B1(n6716), .B2(n6650), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n6733), .A(n2466), .ZN(n6649) );
  NAND2_X1 U5715 ( .A1(\UUT/jar_in [17]), .A2(n297), .ZN(n6490) );
  NAND2_X1 U5716 ( .A1(n298), .A2(\UUT/branch_rega [17]), .ZN(n6491) );
  NAND2_X1 U5717 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [17]), .A2(n299), 
        .ZN(n6492) );
  AND3_X2 U5718 ( .A1(n6490), .A2(n6491), .A3(n6492), .ZN(n420) );
  OAI222_X4 U5719 ( .A1(n5503), .A2(n5530), .B1(n6364), .B2(n2223), .C1(n5528), 
        .C2(n5501), .ZN(\UUT/branch_rega [17]) );
  NAND2_X1 U5720 ( .A1(n908), .A2(\UUT/break_code[4] ), .ZN(n6493) );
  NAND2_X1 U5721 ( .A1(n6715), .A2(\UUT/Mcontrol/Nextpc_decoding/Bta [4]), 
        .ZN(n6494) );
  AND2_X2 U5722 ( .A1(n6493), .A2(n6494), .ZN(n2536) );
  AND3_X1 U5723 ( .A1(n6530), .A2(n6545), .A3(n6544), .ZN(n6640) );
  AOI22_X2 U5724 ( .A1(n6263), .A2(n2328), .B1(n2329), .B2(
        \UUT/Mcontrol/d_sampled_finstr [2]), .ZN(n764) );
  NAND2_X1 U5725 ( .A1(n6630), .A2(n6631), .ZN(n6495) );
  NAND2_X1 U5726 ( .A1(n296), .A2(n6496), .ZN(n2963) );
  INV_X1 U5727 ( .A(n6495), .ZN(n6496) );
  NAND2_X1 U5728 ( .A1(\UUT/jar_in [22]), .A2(n297), .ZN(n6497) );
  NAND2_X1 U5729 ( .A1(n298), .A2(\UUT/branch_rega [22]), .ZN(n6498) );
  NAND2_X1 U5730 ( .A1(n6511), .A2(\UUT/Mcontrol/Nextpc_decoding/Bta [22]), 
        .ZN(n6499) );
  AND3_X2 U5731 ( .A1(n6497), .A2(n6498), .A3(n6499), .ZN(n296) );
  OAI22_X1 U5732 ( .A1(n6297), .A2(n6489), .B1(n6298), .B2(
        \UUT/Mcontrol/Nextpc_decoding/N242 ), .ZN(n6294) );
  BUF_X8 U5733 ( .A(\UUT/Mpath/out_regB[2] ), .Z(n6899) );
  AND2_X1 U5734 ( .A1(\UUT/Mpath/out_regA[4] ), .A2(n6897), .ZN(
        \UUT/Mpath/the_alu/N121 ) );
  OR2_X1 U5735 ( .A1(\UUT/Mpath/out_regA[4] ), .A2(n6897), .ZN(
        \UUT/Mpath/the_alu/N153 ) );
  NAND2_X1 U5736 ( .A1(\UUT/jar_in [16]), .A2(n297), .ZN(n6500) );
  NAND2_X1 U5737 ( .A1(n298), .A2(\UUT/branch_rega [16]), .ZN(n6501) );
  NAND2_X1 U5738 ( .A1(n299), .A2(\UUT/Mcontrol/Nextpc_decoding/Bta [16]), 
        .ZN(n6502) );
  AND3_X2 U5739 ( .A1(n6500), .A2(n6501), .A3(n6502), .ZN(n442) );
  OAI222_X4 U5740 ( .A1(n5506), .A2(n5530), .B1(n6364), .B2(n2243), .C1(n5528), 
        .C2(n5504), .ZN(\UUT/branch_rega [16]) );
  NOR2_X1 U5741 ( .A1(n6725), .A2(n6504), .ZN(n6862) );
  NAND2_X1 U5742 ( .A1(n6505), .A2(n6876), .ZN(n6504) );
  AND2_X2 U5743 ( .A1(n6868), .A2(n6712), .ZN(n6505) );
  OR2_X1 U5744 ( .A1(n6716), .A2(n6849), .ZN(n6506) );
  OR2_X1 U5745 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N125 ), .A2(n6867), .ZN(
        n6507) );
  NAND3_X1 U5746 ( .A1(n6506), .A2(n6507), .A3(n2512), .ZN(n6848) );
  INV_X1 U5747 ( .A(\UUT/jar_in [5]), .ZN(n6849) );
  INV_X1 U5748 ( .A(\UUT/branch_rega [5]), .ZN(n6867) );
  OAI21_X1 U5749 ( .B1(n6710), .B2(n2560), .A(n2561), .ZN(n907) );
  INV_X1 U5750 ( .A(n6654), .ZN(n666) );
  NOR2_X1 U5751 ( .A1(n6615), .A2(n6693), .ZN(n6714) );
  NAND2_X1 U5752 ( .A1(n6596), .A2(n6597), .ZN(n6508) );
  NAND2_X1 U5753 ( .A1(n350), .A2(n6509), .ZN(n3043) );
  INV_X1 U5754 ( .A(n6508), .ZN(n6509) );
  AND2_X1 U5755 ( .A1(n6714), .A2(n295), .ZN(n6510) );
  OR2_X1 U5756 ( .A1(n6716), .A2(n6856), .ZN(n6512) );
  OR2_X1 U5757 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N125 ), .A2(n6857), .ZN(
        n6513) );
  NAND3_X1 U5758 ( .A1(n6512), .A2(n6513), .A3(n2536), .ZN(n6855) );
  INV_X1 U5759 ( .A(\UUT/jar_in [4]), .ZN(n6856) );
  INV_X1 U5760 ( .A(\UUT/branch_rega [4]), .ZN(n6857) );
  NAND2_X1 U5761 ( .A1(n6623), .A2(n6624), .ZN(n6514) );
  NAND2_X1 U5762 ( .A1(n420), .A2(n6515), .ZN(n3163) );
  INV_X1 U5763 ( .A(n6514), .ZN(n6515) );
  OR2_X2 U5764 ( .A1(n6516), .A2(n6576), .ZN(n6690) );
  NAND2_X1 U5765 ( .A1(n6530), .A2(n6696), .ZN(n6516) );
  BUF_X1 U5766 ( .A(\UUT/Mpath/the_mult/Mult_out[1] ), .Z(n6517) );
  BUF_X1 U5767 ( .A(\UUT/Mpath/the_mult/Mult_out[2] ), .Z(n6518) );
  NOR2_X1 U5768 ( .A1(n6522), .A2(n6666), .ZN(n1261) );
  NAND2_X1 U5769 ( .A1(n6523), .A2(n6524), .ZN(n6522) );
  NOR2_X1 U5770 ( .A1(\UUT/branch_rega [26]), .A2(n6745), .ZN(n6519) );
  NAND2_X1 U5771 ( .A1(n1248), .A2(n1247), .ZN(n6520) );
  NAND2_X1 U5772 ( .A1(n1249), .A2(n6521), .ZN(n5578) );
  INV_X1 U5773 ( .A(n6520), .ZN(n6521) );
  NAND2_X1 U5774 ( .A1(\UUT/Mpath/the_alu/diff[30] ), .A2(n1210), .ZN(n6523)
         );
  NAND2_X1 U5775 ( .A1(n1208), .A2(n1262), .ZN(n6524) );
  AND2_X2 U5776 ( .A1(n6503), .A2(\UUT/jar_in [10]), .ZN(n6676) );
  AND2_X2 U5777 ( .A1(n6503), .A2(\UUT/jar_in [9]), .ZN(n6672) );
  BUF_X1 U5778 ( .A(\UUT/Mpath/out_regA[0] ), .Z(n6525) );
  NAND2_X1 U5779 ( .A1(n908), .A2(\UUT/break_code[5] ), .ZN(n6526) );
  NAND2_X1 U5780 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [5]), .A2(n6715), 
        .ZN(n6527) );
  AND2_X2 U5781 ( .A1(n6527), .A2(n6526), .ZN(n2512) );
  INV_X1 U5782 ( .A(n6647), .ZN(n740) );
  NAND2_X1 U5783 ( .A1(n935), .A2(\UUT/Mcontrol/d_instr [6]), .ZN(n6528) );
  NAND2_X1 U5784 ( .A1(n6086), .A2(n6529), .ZN(n2076) );
  INV_X1 U5785 ( .A(n6528), .ZN(n6529) );
  NAND2_X2 U5786 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1945 ), .A2(n6067), 
        .ZN(n6057) );
  INV_X2 U5787 ( .A(n6046), .ZN(n6079) );
  NOR2_X2 U5788 ( .A1(n6079), .A2(n6057), .ZN(n6045) );
  NAND2_X1 U5789 ( .A1(\UUT/Mpath/the_alu/diff[31] ), .A2(n1210), .ZN(n6530)
         );
  OAI22_X2 U5790 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6287), .B1(
        n6288), .B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6693) );
  OAI21_X1 U5791 ( .B1(n6479), .B2(n2560), .A(n2561), .ZN(n6531) );
  NAND3_X2 U5792 ( .A1(n6328), .A2(n6040), .A3(n6210), .ZN(n6053) );
  OR2_X1 U5793 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1889 ) );
  OR2_X1 U5794 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1916 ) );
  OR2_X1 U5795 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1878 ) );
  OR2_X1 U5796 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1923 ) );
  OR2_X1 U5797 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1947 ) );
  OR2_X1 U5798 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1929 ) );
  OR2_X1 U5799 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1935 ) );
  OR2_X1 U5800 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1953 ) );
  OR2_X1 U5801 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1941 ) );
  OR2_X1 U5802 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1965 ) );
  OR2_X1 U5803 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1875 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1959 ) );
  BUF_X2 U5804 ( .A(n6531), .Z(n6716) );
  INV_X1 U5805 ( .A(n6686), .ZN(n545) );
  NOR2_X1 U5806 ( .A1(n6575), .A2(n6532), .ZN(n6819) );
  NAND2_X1 U5807 ( .A1(n6533), .A2(n6820), .ZN(n6532) );
  AND2_X1 U5808 ( .A1(n6549), .A2(n6823), .ZN(n6533) );
  NAND2_X1 U5809 ( .A1(n1242), .A2(n1241), .ZN(n6534) );
  NAND2_X1 U5810 ( .A1(n1243), .A2(n6535), .ZN(n5585) );
  INV_X1 U5811 ( .A(n6534), .ZN(n6535) );
  NAND2_X1 U5812 ( .A1(\UUT/jar_in [1]), .A2(n6711), .ZN(n6536) );
  NAND2_X1 U5813 ( .A1(n298), .A2(\UUT/branch_rega [1]), .ZN(n6537) );
  NAND2_X1 U5814 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [1]), .A2(n299), .ZN(
        n6538) );
  BUF_X1 U5815 ( .A(\UUT/Mcontrol/d_instr [28]), .Z(n6539) );
  BUF_X4 U5816 ( .A(\UUT/Mcontrol/d_instr [28]), .Z(n6541) );
  BUF_X1 U5817 ( .A(\UUT/Mcontrol/d_instr [28]), .Z(n6540) );
  BUF_X1 U5818 ( .A(n5563), .Z(n6542) );
  OR2_X1 U5819 ( .A1(\UUT/Mpath/out_regA[3] ), .A2(n6898), .ZN(
        \UUT/Mpath/the_alu/N154 ) );
  AND2_X1 U5820 ( .A1(\UUT/Mpath/out_regA[3] ), .A2(n6898), .ZN(
        \UUT/Mpath/the_alu/N122 ) );
  OR2_X1 U5821 ( .A1(\localbus/c1_addr_outbus[30] ), .A2(n6910), .ZN(n6543) );
  NAND2_X1 U5822 ( .A1(n6543), .A2(n6909), .ZN(\localbus/N56 ) );
  NAND2_X1 U5823 ( .A1(n1208), .A2(n1209), .ZN(n6544) );
  NAND2_X1 U5824 ( .A1(\UUT/Mpath/the_alu/sum[31] ), .A2(n1211), .ZN(n6545) );
  OR2_X1 U5825 ( .A1(\UUT/branch_rega [28]), .A2(\UUT/branch_rega [29]), .ZN(
        n6875) );
  AND3_X2 U5826 ( .A1(n6546), .A2(n6547), .A3(n6548), .ZN(n1255) );
  INV_X32 U5827 ( .A(n6629), .ZN(n6546) );
  NAND2_X1 U5828 ( .A1(\UUT/Mpath/the_alu/diff[29] ), .A2(n1210), .ZN(n6547)
         );
  NAND2_X1 U5829 ( .A1(\UUT/Mpath/the_alu/sum[29] ), .A2(n1211), .ZN(n6548) );
  OR2_X2 U5830 ( .A1(n5462), .A2(n5528), .ZN(n6608) );
  AND2_X2 U5831 ( .A1(n6825), .A2(n6723), .ZN(n6720) );
  INV_X1 U5832 ( .A(n6752), .ZN(n6753) );
  INV_X1 U5833 ( .A(\UUT/Mcontrol/Nextpc_decoding/N191 ), .ZN(n6808) );
  NOR2_X2 U5834 ( .A1(n6806), .A2(\UUT/branch_rega [29]), .ZN(n6736) );
  AND2_X1 U5835 ( .A1(n6891), .A2(n6574), .ZN(n6549) );
  NOR2_X2 U5836 ( .A1(n6850), .A2(n6550), .ZN(n6838) );
  NAND2_X1 U5837 ( .A1(n6697), .A2(n6885), .ZN(n6550) );
  NAND2_X1 U5838 ( .A1(n1236), .A2(n1235), .ZN(n6551) );
  NAND2_X1 U5839 ( .A1(n1237), .A2(n6552), .ZN(n5592) );
  INV_X1 U5840 ( .A(n6551), .ZN(n6552) );
  NAND2_X1 U5841 ( .A1(n1237), .A2(n6556), .ZN(n6553) );
  NAND2_X1 U5842 ( .A1(n6553), .A2(n6554), .ZN(n5471) );
  OR2_X1 U5843 ( .A1(n6555), .A2(n5564), .ZN(n6554) );
  INV_X1 U5844 ( .A(n6578), .ZN(n6555) );
  AND2_X1 U5845 ( .A1(n6552), .A2(n6578), .ZN(n6556) );
  OAI222_X4 U5846 ( .A1(n5465), .A2(n5528), .B1(n5417), .B2(n6364), .C1(n5467), 
        .C2(n5530), .ZN(\UUT/branch_rega [28]) );
  AOI222_X2 U5847 ( .A1(n1208), .A2(n1250), .B1(\UUT/Mpath/the_alu/diff[28] ), 
        .B2(n1210), .C1(\UUT/Mpath/the_alu/sum[28] ), .C2(n1211), .ZN(n1249)
         );
  AOI22_X2 U5848 ( .A1(n5577), .A2(\UUT/Mpath/N119 ), .B1(n5578), .B2(n5564), 
        .ZN(n5465) );
  INV_X1 U5849 ( .A(n6713), .ZN(n6557) );
  NAND2_X1 U5850 ( .A1(n6558), .A2(n6559), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N222 ) );
  AND2_X2 U5851 ( .A1(n6829), .A2(n6813), .ZN(n6558) );
  NOR2_X2 U5852 ( .A1(n6671), .A2(n6557), .ZN(n6559) );
  NAND2_X1 U5853 ( .A1(n1254), .A2(n1253), .ZN(n6560) );
  INV_X1 U5854 ( .A(n6560), .ZN(n6561) );
  NAND2_X1 U5855 ( .A1(\UUT/jar_in [18]), .A2(n6711), .ZN(n6562) );
  NAND2_X1 U5856 ( .A1(n298), .A2(\UUT/branch_rega [18]), .ZN(n6563) );
  NAND2_X1 U5857 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [18]), .A2(n6511), 
        .ZN(n6564) );
  AND3_X2 U5858 ( .A1(n6562), .A2(n6563), .A3(n6564), .ZN(n398) );
  OAI222_X4 U5859 ( .A1(n5462), .A2(n5430), .B1(n5463), .B2(n5432), .C1(n5464), 
        .C2(n5434), .ZN(\UUT/branch_regb [29]) );
  NAND2_X1 U5860 ( .A1(n6609), .A2(n6610), .ZN(n6565) );
  NAND2_X2 U5861 ( .A1(n6608), .A2(n6566), .ZN(\UUT/branch_rega [29]) );
  INV_X1 U5862 ( .A(n6565), .ZN(n6566) );
  OR2_X1 U5863 ( .A1(n369), .A2(n294), .ZN(n6567) );
  OR2_X1 U5864 ( .A1(n295), .A2(n2648), .ZN(n6568) );
  NAND3_X1 U5865 ( .A1(n6567), .A2(n6568), .A3(n372), .ZN(n3083) );
  NAND2_X1 U5866 ( .A1(\UUT/jar_in [19]), .A2(n6711), .ZN(n6569) );
  NAND2_X1 U5867 ( .A1(n298), .A2(\UUT/branch_rega [19]), .ZN(n6570) );
  NAND2_X1 U5868 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [19]), .A2(n6511), 
        .ZN(n6571) );
  AND3_X2 U5869 ( .A1(n6569), .A2(n6570), .A3(n6571), .ZN(n372) );
  OR2_X1 U5870 ( .A1(n5464), .A2(n5530), .ZN(n6610) );
  NAND2_X1 U5871 ( .A1(n908), .A2(\UUT/break_code[10] ), .ZN(n6572) );
  OR2_X2 U5872 ( .A1(n5456), .A2(n5528), .ZN(n6663) );
  AND2_X1 U5873 ( .A1(\UUT/Mpath/out_regA[2] ), .A2(n6899), .ZN(
        \UUT/Mpath/the_alu/N123 ) );
  OR2_X1 U5874 ( .A1(\UUT/Mpath/out_regA[2] ), .A2(n6899), .ZN(
        \UUT/Mpath/the_alu/N155 ) );
  INV_X1 U5875 ( .A(n6828), .ZN(n6574) );
  NAND2_X1 U5876 ( .A1(n6838), .A2(n6836), .ZN(n6575) );
  AND2_X1 U5877 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N159 ), .A2(n6870), .ZN(
        n6829) );
  AND2_X2 U5878 ( .A1(n6819), .A2(n6814), .ZN(n6813) );
  OAI22_X4 U5879 ( .A1(\UUT/Mpath/the_alu/N520 ), .A2(n2575), .B1(
        \UUT/Mpath/the_alu/N526 ), .B2(\UUT/Mpath/the_alu/N468 ), .ZN(n1211)
         );
  OR2_X2 U5880 ( .A1(n6755), .A2(\UUT/branch_rega [6]), .ZN(n6754) );
  INV_X8 U5881 ( .A(n6720), .ZN(n6721) );
  INV_X1 U5882 ( .A(\UUT/branch_rega [6]), .ZN(n6724) );
  OAI222_X4 U5883 ( .A1(n5443), .A2(n5530), .B1(n6364), .B2(n2491), .C1(n5528), 
        .C2(n5441), .ZN(\UUT/branch_rega [6]) );
  NAND2_X1 U5884 ( .A1(n6545), .A2(n6577), .ZN(n6576) );
  INV_X32 U5885 ( .A(n6632), .ZN(n6577) );
  OR2_X2 U5886 ( .A1(\UUT/branch_rega [26]), .A2(\UUT/branch_rega [25]), .ZN(
        n6858) );
  AND2_X2 U5887 ( .A1(\UUT/Mpath/the_alu/sum[27] ), .A2(n1211), .ZN(n6591) );
  INV_X32 U5888 ( .A(n6700), .ZN(n6578) );
  NOR2_X2 U5889 ( .A1(n6742), .A2(n6579), .ZN(n6789) );
  NAND2_X1 U5890 ( .A1(n6580), .A2(n6783), .ZN(n6579) );
  AND2_X2 U5891 ( .A1(n6811), .A2(n6719), .ZN(n6580) );
  NAND2_X1 U5892 ( .A1(n6663), .A2(n6581), .ZN(n6689) );
  OR2_X1 U5893 ( .A1(n117), .A2(n294), .ZN(n6582) );
  OR2_X1 U5894 ( .A1(n295), .A2(n2727), .ZN(n6583) );
  NAND2_X1 U5895 ( .A1(\UUT/jar_in [23]), .A2(n297), .ZN(n6584) );
  NAND2_X1 U5896 ( .A1(n298), .A2(\UUT/branch_rega [23]), .ZN(n6585) );
  NAND2_X1 U5897 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [23]), .A2(n6510), 
        .ZN(n6586) );
  AND3_X2 U5898 ( .A1(n6586), .A2(n6585), .A3(n6584), .ZN(n905) );
  OAI222_X1 U5899 ( .A1(n6446), .A2(n6026), .B1(n6163), .B2(n5881), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n6035), .ZN(n6272) );
  NAND3_X2 U5900 ( .A1(n6028), .A2(\UUT/Mcontrol/Operation_decoding32/N2036 ), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N2030 ), .ZN(n6587) );
  INV_X4 U5901 ( .A(n6587), .ZN(n931) );
  INV_X1 U5902 ( .A(\UUT/Mcontrol/Operation_decoding32/N2036 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2037 ) );
  OR2_X1 U5903 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2035 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2036 ) );
  BUF_X1 U5904 ( .A(\UUT/break_code[0] ), .Z(n6588) );
  OAI222_X4 U5905 ( .A1(n5485), .A2(n5530), .B1(n6364), .B2(n2098), .C1(n5528), 
        .C2(n5483), .ZN(\UUT/branch_rega [22]) );
  OR2_X1 U5906 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2086 ) );
  OR2_X1 U5907 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2080 ) );
  OR2_X1 U5908 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2074 ) );
  OR2_X1 U5909 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2068 ) );
  OR2_X1 U5910 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2062 ) );
  OR2_X1 U5911 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2056 ) );
  OR2_X1 U5912 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2050 ) );
  OR2_X1 U5913 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2020 ) );
  OR2_X1 U5914 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2014 ) );
  OR2_X1 U5915 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2008 ) );
  OR2_X1 U5916 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2002 ) );
  OR2_X1 U5917 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1996 ) );
  OR2_X1 U5918 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1990 ) );
  OR2_X1 U5919 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1983 ) );
  OR2_X1 U5920 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1971 ) );
  OR2_X1 U5921 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2026 ) );
  OR2_X1 U5922 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2032 ) );
  OR2_X1 U5923 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2038 ) );
  OR2_X1 U5924 ( .A1(\UUT/Mcontrol/d_instr [30]), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2044 ) );
  OR2_X1 U5925 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1876 ), .A2(
        \UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1977 ) );
  AND2_X2 U5926 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1969 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1963 ), .ZN(n6210) );
  INV_X1 U5927 ( .A(\UUT/Mcontrol/Operation_decoding32/N1969 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1970 ) );
  INV_X1 U5928 ( .A(\UUT/Mcontrol/Operation_decoding32/N1963 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1964 ) );
  OAI222_X4 U5929 ( .A1(n6029), .A2(n6446), .B1(n6163), .B2(n6035), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n6032), .ZN(n6181) );
  OAI222_X4 U5930 ( .A1(n6031), .A2(n6446), .B1(n6163), .B2(n6036), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n6033), .ZN(n6188) );
  OAI222_X4 U5931 ( .A1(n6034), .A2(n6128), .B1(n6163), .B2(n5889), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1975 ), .C2(n6036), .ZN(n6278) );
  AND2_X1 U5932 ( .A1(n1208), .A2(n1244), .ZN(n6589) );
  AND2_X1 U5933 ( .A1(\UUT/Mpath/the_alu/diff[27] ), .A2(n1210), .ZN(n6590) );
  NOR3_X2 U5934 ( .A1(n6589), .A2(n6590), .A3(n6591), .ZN(n1243) );
  OR2_X2 U5935 ( .A1(n5468), .A2(n5528), .ZN(n6592) );
  OR2_X1 U5936 ( .A1(n5418), .A2(n6364), .ZN(n6593) );
  OR2_X2 U5937 ( .A1(n5470), .A2(n5530), .ZN(n6594) );
  NAND3_X2 U5938 ( .A1(n6592), .A2(n6593), .A3(n6594), .ZN(
        \UUT/branch_rega [27]) );
  AND2_X2 U5939 ( .A1(n6827), .A2(n6851), .ZN(n6826) );
  INV_X4 U5940 ( .A(\UUT/branch_rega [16]), .ZN(n6851) );
  INV_X4 U5941 ( .A(\UUT/branch_rega [16]), .ZN(n6853) );
  NAND2_X1 U5942 ( .A1(n6803), .A2(n6884), .ZN(n6788) );
  NOR2_X1 U5943 ( .A1(n6743), .A2(n6751), .ZN(n6735) );
  INV_X1 U5944 ( .A(n6802), .ZN(n6803) );
  NAND2_X4 U5945 ( .A1(n6155), .A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n6163) );
  INV_X4 U5946 ( .A(n6595), .ZN(n4351) );
  OR2_X1 U5947 ( .A1(n348), .A2(n294), .ZN(n6596) );
  OR2_X1 U5948 ( .A1(n295), .A2(n2645), .ZN(n6597) );
  OR2_X4 U5949 ( .A1(\localbus/N57 ), .A2(\localbus/N62 ), .ZN(n4337) );
  NAND2_X4 U5950 ( .A1(n4337), .A2(\localbus/N338 ), .ZN(\localbus/N227 ) );
  INV_X4 U5951 ( .A(n6071), .ZN(\UUT/Mcontrol/d_instr [29]) );
  AOI22_X2 U5952 ( .A1(n935), .A2(n6085), .B1(n6030), .B2(n2077), .ZN(n2061)
         );
  INV_X4 U5953 ( .A(n6070), .ZN(\UUT/Mcontrol/d_instr [30]) );
  OR2_X1 U5954 ( .A1(n327), .A2(n294), .ZN(n6598) );
  OR2_X1 U5955 ( .A1(n295), .A2(n2642), .ZN(n6599) );
  NAND3_X1 U5956 ( .A1(n6598), .A2(n6599), .A3(n329), .ZN(n3003) );
  NAND2_X1 U5957 ( .A1(\UUT/jar_in [21]), .A2(n297), .ZN(n6600) );
  NAND2_X1 U5958 ( .A1(n298), .A2(n6464), .ZN(n6601) );
  NAND2_X1 U5959 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [21]), .A2(n6510), 
        .ZN(n6602) );
  AND3_X2 U5960 ( .A1(n6600), .A2(n6601), .A3(n6602), .ZN(n329) );
  OR2_X1 U5961 ( .A1(n6658), .A2(n6603), .ZN(n6604) );
  INV_X1 U5962 ( .A(n6790), .ZN(n6603) );
  AND2_X1 U5963 ( .A1(n6605), .A2(n6789), .ZN(n6660) );
  INV_X32 U5964 ( .A(n6604), .ZN(n6605) );
  OR2_X1 U5965 ( .A1(n495), .A2(n294), .ZN(n6606) );
  OR2_X1 U5966 ( .A1(n295), .A2(n2663), .ZN(n6607) );
  NAND3_X1 U5967 ( .A1(n6606), .A2(n6607), .A3(n497), .ZN(n3283) );
  OR2_X1 U5968 ( .A1(n5416), .A2(n6364), .ZN(n6609) );
  NAND2_X1 U5969 ( .A1(\UUT/jar_in [14]), .A2(n297), .ZN(n6611) );
  NAND2_X1 U5970 ( .A1(n298), .A2(\UUT/branch_rega [14]), .ZN(n6612) );
  NAND2_X1 U5971 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [14]), .A2(n6511), 
        .ZN(n6613) );
  AND3_X2 U5972 ( .A1(n6611), .A2(n6612), .A3(n6613), .ZN(n497) );
  OAI222_X4 U5973 ( .A1(n5512), .A2(n5530), .B1(n6364), .B2(n2283), .C1(n5528), 
        .C2(n5510), .ZN(\UUT/branch_rega [14]) );
  OAI222_X4 U5974 ( .A1(n5468), .A2(n5430), .B1(n5469), .B2(n5432), .C1(n5470), 
        .C2(n5434), .ZN(\UUT/branch_regb [27]) );
  INV_X1 U5975 ( .A(\UUT/branch_rega [27]), .ZN(n6744) );
  INV_X1 U5976 ( .A(\UUT/branch_rega [27]), .ZN(n6841) );
  NOR2_X1 U5977 ( .A1(n2559), .A2(n2560), .ZN(n6614) );
  INV_X1 U5978 ( .A(n6614), .ZN(n6615) );
  NAND2_X1 U5979 ( .A1(\UUT/jar_in [15]), .A2(n6711), .ZN(n6616) );
  NAND2_X1 U5980 ( .A1(n298), .A2(\UUT/branch_rega [15]), .ZN(n6617) );
  NAND2_X1 U5981 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [15]), .A2(n6510), 
        .ZN(n6618) );
  OAI222_X4 U5982 ( .A1(n5509), .A2(n5530), .B1(n6364), .B2(n2263), .C1(n5528), 
        .C2(n5507), .ZN(\UUT/branch_rega [15]) );
  INV_X4 U5983 ( .A(n6069), .ZN(\UUT/Mcontrol/d_instr [31]) );
  INV_X1 U5984 ( .A(\UUT/Mcontrol/Operation_decoding32/N1920 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N89 ) );
  NAND2_X1 U5985 ( .A1(n6664), .A2(n6665), .ZN(n6621) );
  NAND2_X2 U5986 ( .A1(n6663), .A2(n6622), .ZN(\UUT/branch_rega [30]) );
  INV_X1 U5987 ( .A(n6621), .ZN(n6622) );
  OR2_X1 U5988 ( .A1(n417), .A2(n294), .ZN(n6623) );
  OR2_X1 U5989 ( .A1(n295), .A2(n2654), .ZN(n6624) );
  OR2_X1 U5990 ( .A1(n5458), .A2(n5530), .ZN(n6665) );
  BUF_X4 U5991 ( .A(\UUT/Mpath/out_regB[4] ), .Z(n6897) );
  BUF_X1 U5992 ( .A(n5456), .Z(n6625) );
  AOI22_X2 U5993 ( .A1(n5584), .A2(\UUT/Mpath/N119 ), .B1(n5585), .B2(n5564), 
        .ZN(n5468) );
  NOR2_X1 U5994 ( .A1(n6785), .A2(n6658), .ZN(n6626) );
  AND2_X1 U5995 ( .A1(n6626), .A2(n6627), .ZN(n6831) );
  AND2_X1 U5996 ( .A1(n6628), .A2(n6659), .ZN(n6627) );
  INV_X1 U5997 ( .A(n6657), .ZN(n6628) );
  AND2_X1 U5998 ( .A1(n1208), .A2(n1256), .ZN(n6629) );
  OR2_X1 U5999 ( .A1(n292), .A2(n294), .ZN(n6630) );
  OR2_X1 U6000 ( .A1(n295), .A2(n2639), .ZN(n6631) );
  AND2_X1 U6001 ( .A1(n1208), .A2(n1209), .ZN(n6632) );
  NOR2_X1 U6002 ( .A1(n6777), .A2(n6657), .ZN(n6634) );
  AND2_X1 U6003 ( .A1(n6635), .A2(n6636), .ZN(n6681) );
  NOR2_X1 U6004 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N160 ), .A2(
        \UUT/branch_rega [29]), .ZN(n6635) );
  NOR2_X1 U6005 ( .A1(n6683), .A2(\UUT/branch_rega [28]), .ZN(n6636) );
  INV_X4 U6006 ( .A(n6637), .ZN(\localbus/c1_op[SLAVE][0] ) );
  BUF_X1 U6007 ( .A(n6531), .Z(n6638) );
  NOR3_X2 U6008 ( .A1(n6672), .A2(n6451), .A3(n6673), .ZN(n909) );
  OAI22_X1 U6009 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6287), .B1(
        n6288), .B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6639) );
  NOR3_X1 U6010 ( .A1(n6672), .A2(n6673), .A3(n6451), .ZN(n6642) );
  NOR3_X1 U6011 ( .A1(n6676), .A2(n6677), .A3(n6462), .ZN(n6643) );
  NAND2_X1 U6012 ( .A1(n6640), .A2(n6696), .ZN(n6644) );
  AOI21_X1 U6013 ( .B1(n6289), .B2(n6290), .A(n6291), .ZN(n6288) );
  OAI221_X1 U6014 ( .B1(n6716), .B2(n6648), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n6876), .A(n2558), .ZN(n6647) );
  INV_X4 U6015 ( .A(\UUT/branch_rega [3]), .ZN(n6876) );
  OAI222_X4 U6016 ( .A1(n5440), .A2(n5530), .B1(n6364), .B2(n2468), .C1(n5528), 
        .C2(n5438), .ZN(\UUT/branch_rega [7]) );
  INV_X1 U6017 ( .A(n6453), .ZN(n6674) );
  AND2_X1 U6018 ( .A1(n6489), .A2(\UUT/Mcontrol/Nextpc_decoding/N236 ), .ZN(
        n6651) );
  NOR2_X1 U6019 ( .A1(n6299), .A2(n6651), .ZN(n6298) );
  NAND2_X1 U6020 ( .A1(n6646), .A2(\UUT/jar_in [8]), .ZN(n6652) );
  NAND2_X1 U6021 ( .A1(n2325), .A2(\UUT/branch_rega [8]), .ZN(n6653) );
  AND3_X2 U6022 ( .A1(n6652), .A2(n6653), .A3(n2443), .ZN(n631) );
  INV_X1 U6023 ( .A(\UUT/Mcontrol/Nextpc_decoding/N235 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N236 ) );
  OAI222_X4 U6024 ( .A1(n5437), .A2(n5530), .B1(n5529), .B2(n2445), .C1(n5528), 
        .C2(n5435), .ZN(\UUT/branch_rega [8]) );
  OAI221_X1 U6025 ( .B1(n6638), .B2(n6655), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n6656), .A(n2489), .ZN(n6654) );
  INV_X32 U6026 ( .A(\UUT/branch_rega [6]), .ZN(n6656) );
  NAND2_X1 U6027 ( .A1(n6779), .A2(n6832), .ZN(n6657) );
  INV_X1 U6028 ( .A(n6847), .ZN(n6658) );
  NAND2_X1 U6029 ( .A1(n6660), .A2(n6659), .ZN(n6777) );
  INV_X32 U6030 ( .A(n6784), .ZN(n6659) );
  OR2_X1 U6031 ( .A1(n520), .A2(n294), .ZN(n6661) );
  OR2_X1 U6032 ( .A1(n295), .A2(n2666), .ZN(n6662) );
  NAND3_X1 U6033 ( .A1(n6661), .A2(n6662), .A3(n522), .ZN(n3323) );
  OR2_X1 U6034 ( .A1(n5415), .A2(n6364), .ZN(n6664) );
  AND2_X1 U6035 ( .A1(\UUT/Mpath/the_alu/sum[30] ), .A2(n1211), .ZN(n6666) );
  NAND2_X1 U6036 ( .A1(\UUT/jar_in [13]), .A2(n297), .ZN(n6667) );
  NAND2_X1 U6037 ( .A1(n298), .A2(\UUT/branch_rega [13]), .ZN(n6668) );
  NAND2_X1 U6038 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [13]), .A2(n6510), 
        .ZN(n6669) );
  AND3_X2 U6039 ( .A1(n6667), .A2(n6668), .A3(n6669), .ZN(n522) );
  OAI222_X4 U6040 ( .A1(n5515), .A2(n5530), .B1(n6364), .B2(n2303), .C1(n5528), 
        .C2(n5513), .ZN(\UUT/branch_rega [13]) );
  INV_X1 U6041 ( .A(n6705), .ZN(n6670) );
  NAND2_X1 U6042 ( .A1(n6886), .A2(n6670), .ZN(n6671) );
  AND2_X1 U6043 ( .A1(n2325), .A2(\UUT/branch_rega [9]), .ZN(n6673) );
  OR2_X2 U6044 ( .A1(\UUT/branch_rega [13]), .A2(\UUT/branch_rega [12]), .ZN(
        n6865) );
  INV_X1 U6045 ( .A(\UUT/branch_rega [12]), .ZN(n6807) );
  INV_X1 U6046 ( .A(\UUT/branch_rega [12]), .ZN(n6886) );
  OAI222_X4 U6047 ( .A1(n5518), .A2(n5530), .B1(n6364), .B2(n2353), .C1(n5528), 
        .C2(n5516), .ZN(\UUT/branch_rega [12]) );
  INV_X1 U6048 ( .A(n6858), .ZN(n6859) );
  AND2_X1 U6049 ( .A1(n2325), .A2(\UUT/branch_rega [10]), .ZN(n6677) );
  OAI222_X4 U6050 ( .A1(n5524), .A2(n5530), .B1(n6364), .B2(n2399), .C1(n5528), 
        .C2(n5522), .ZN(\UUT/branch_rega [10]) );
  NOR2_X1 U6051 ( .A1(n2559), .A2(n2560), .ZN(n6678) );
  NOR2_X1 U6052 ( .A1(\UUT/Mcontrol/Nextpc_decoding/condition ), .A2(n6679), 
        .ZN(n906) );
  INV_X1 U6053 ( .A(n6678), .ZN(n6679) );
  OR2_X1 U6054 ( .A1(n6489), .A2(\UUT/branch_rega [30]), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N160 ) );
  INV_X1 U6055 ( .A(n6809), .ZN(n6680) );
  NAND2_X1 U6056 ( .A1(n6681), .A2(n6682), .ZN(n6725) );
  NOR2_X1 U6057 ( .A1(\UUT/branch_rega [26]), .A2(n6680), .ZN(n6682) );
  INV_X1 U6058 ( .A(n6841), .ZN(n6683) );
  NAND2_X1 U6059 ( .A1(n6646), .A2(\UUT/jar_in [2]), .ZN(n6684) );
  NAND2_X1 U6060 ( .A1(n2325), .A2(\UUT/branch_rega [2]), .ZN(n6685) );
  AND3_X2 U6061 ( .A1(n6684), .A2(n6685), .A3(n2327), .ZN(n763) );
  OAI222_X4 U6062 ( .A1(n5461), .A2(n5530), .B1(n5529), .B2(n2330), .C1(n5528), 
        .C2(n5459), .ZN(\UUT/branch_rega [2]) );
  NOR2_X1 U6063 ( .A1(n6689), .A2(n6488), .ZN(n6845) );
  OR2_X1 U6064 ( .A1(n439), .A2(n294), .ZN(n6691) );
  OR2_X1 U6065 ( .A1(n295), .A2(n2657), .ZN(n6692) );
  NAND3_X1 U6066 ( .A1(n6691), .A2(n6692), .A3(n442), .ZN(n3203) );
  NAND2_X2 U6067 ( .A1(n137), .A2(n863), .ZN(n6694) );
  NAND2_X1 U6068 ( .A1(n1205), .A2(n1206), .ZN(n6695) );
  INV_X1 U6069 ( .A(n6695), .ZN(n6696) );
  OR2_X2 U6070 ( .A1(n6799), .A2(\UUT/branch_rega [3]), .ZN(n6794) );
  OAI222_X4 U6071 ( .A1(n5452), .A2(n5530), .B1(n5529), .B2(n2565), .C1(n5528), 
        .C2(n5450), .ZN(\UUT/branch_rega [3]) );
  OR2_X1 U6072 ( .A1(n6525), .A2(n6675), .ZN(\UUT/Mpath/the_alu/N157 ) );
  AND2_X1 U6073 ( .A1(n6525), .A2(n6675), .ZN(\UUT/Mpath/the_alu/N125 ) );
  NOR2_X1 U6074 ( .A1(n6840), .A2(\UUT/branch_rega [22]), .ZN(n6697) );
  AND2_X1 U6075 ( .A1(n6877), .A2(n6698), .ZN(n6699) );
  INV_X1 U6076 ( .A(\UUT/branch_rega [27]), .ZN(n6698) );
  AND2_X1 U6077 ( .A1(n5591), .A2(\UUT/Mpath/N119 ), .ZN(n6700) );
  NOR2_X1 U6078 ( .A1(n2559), .A2(n2560), .ZN(n6701) );
  INV_X1 U6079 ( .A(n6701), .ZN(n6702) );
  NAND2_X1 U6080 ( .A1(n6646), .A2(\UUT/jar_in [11]), .ZN(n6703) );
  NAND2_X1 U6081 ( .A1(n2325), .A2(\UUT/branch_rega [11]), .ZN(n6704) );
  OR2_X1 U6082 ( .A1(\UUT/branch_rega [14]), .A2(n6706), .ZN(n6705) );
  INV_X1 U6083 ( .A(n6878), .ZN(n6706) );
  AND2_X1 U6084 ( .A1(n1208), .A2(n1238), .ZN(n6707) );
  AND2_X1 U6085 ( .A1(\UUT/Mpath/the_alu/diff[26] ), .A2(n1210), .ZN(n6708) );
  AND2_X1 U6086 ( .A1(\UUT/Mpath/the_alu/sum[26] ), .A2(n1211), .ZN(n6709) );
  NOR3_X2 U6087 ( .A1(n6707), .A2(n6708), .A3(n6709), .ZN(n1237) );
  OAI222_X4 U6088 ( .A1(n5521), .A2(n5530), .B1(n6364), .B2(n2376), .C1(n5528), 
        .C2(n5519), .ZN(\UUT/branch_rega [11]) );
  INV_X1 U6089 ( .A(n6848), .ZN(n694) );
  OAI222_X4 U6090 ( .A1(n5471), .A2(n5430), .B1(n5472), .B2(n5432), .C1(n5473), 
        .C2(n5434), .ZN(\UUT/branch_regb [26]) );
  OAI22_X1 U6091 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6287), .B1(
        n6472), .B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/condition ) );
  NAND2_X4 U6092 ( .A1(net54875), .A2(n978), .ZN(n546) );
  INV_X8 U6093 ( .A(n546), .ZN(n295) );
  INV_X1 U6094 ( .A(n6718), .ZN(n6712) );
  INV_X32 U6095 ( .A(n6721), .ZN(n6713) );
  AND2_X1 U6096 ( .A1(n6882), .A2(n6883), .ZN(net56414) );
  INV_X1 U6097 ( .A(n6726), .ZN(n6717) );
  NAND2_X1 U6098 ( .A1(n6867), .A2(n6717), .ZN(n6718) );
  AND2_X2 U6099 ( .A1(n6740), .A2(n6733), .ZN(n6732) );
  OR2_X2 U6100 ( .A1(n6793), .A2(\UUT/branch_rega [21]), .ZN(n6792) );
  INV_X1 U6101 ( .A(\UUT/branch_rega [18]), .ZN(n6834) );
  OAI222_X4 U6102 ( .A1(n5500), .A2(n5530), .B1(n5529), .B2(n2203), .C1(n5528), 
        .C2(n5498), .ZN(\UUT/branch_rega [18]) );
  AOI222_X2 U6103 ( .A1(n6134), .A2(n5564), .B1(n415), .B2(\UUT/Mpath/N119 ), 
        .C1(\UUT/Mpath/out_jar[18] ), .C2(n5612), .ZN(n5498) );
  INV_X1 U6104 ( .A(n6727), .ZN(n6719) );
  INV_X1 U6105 ( .A(n6753), .ZN(n6722) );
  NOR2_X2 U6106 ( .A1(n6730), .A2(n6722), .ZN(n6723) );
  INV_X4 U6107 ( .A(n6764), .ZN(n6766) );
  NAND2_X1 U6108 ( .A1(n6732), .A2(n6724), .ZN(n6726) );
  NAND2_X1 U6109 ( .A1(n6728), .A2(n6805), .ZN(n6727) );
  AND2_X2 U6110 ( .A1(n6818), .A2(n6729), .ZN(n6728) );
  INV_X1 U6111 ( .A(n6734), .ZN(n6729) );
  NAND2_X1 U6112 ( .A1(n6757), .A2(n6731), .ZN(n6730) );
  INV_X32 U6113 ( .A(n6737), .ZN(n6731) );
  INV_X1 U6114 ( .A(\UUT/branch_rega [7]), .ZN(n6733) );
  NAND2_X1 U6115 ( .A1(n6735), .A2(n6812), .ZN(n6734) );
  OR2_X1 U6116 ( .A1(n6738), .A2(\UUT/branch_rega [9]), .ZN(n6737) );
  INV_X1 U6117 ( .A(n6739), .ZN(n6738) );
  INV_X32 U6118 ( .A(\UUT/branch_rega [8]), .ZN(n6739) );
  AND2_X1 U6119 ( .A1(n6746), .A2(n6741), .ZN(n6740) );
  INV_X1 U6120 ( .A(\UUT/branch_rega [8]), .ZN(n6741) );
  NAND2_X1 U6121 ( .A1(n6822), .A2(n6821), .ZN(n6742) );
  INV_X1 U6122 ( .A(n6807), .ZN(n6743) );
  NAND2_X1 U6123 ( .A1(n6744), .A2(n6852), .ZN(n6745) );
  INV_X1 U6124 ( .A(\UUT/branch_rega [23]), .ZN(n6885) );
  OAI222_X4 U6125 ( .A1(n5482), .A2(n5530), .B1(n6364), .B2(n2078), .C1(n5528), 
        .C2(n5480), .ZN(\UUT/branch_rega [23]) );
  AND2_X1 U6126 ( .A1(n6756), .A2(n6747), .ZN(n6746) );
  INV_X1 U6127 ( .A(\UUT/branch_rega [9]), .ZN(n6747) );
  INV_X1 U6128 ( .A(n6759), .ZN(n6748) );
  NAND2_X1 U6129 ( .A1(n6880), .A2(n6748), .ZN(n6749) );
  INV_X1 U6130 ( .A(n6749), .ZN(n6750) );
  NAND2_X1 U6131 ( .A1(n6830), .A2(n6750), .ZN(n6751) );
  OR2_X1 U6132 ( .A1(\UUT/branch_rega [7]), .A2(n6754), .ZN(n6752) );
  INV_X1 U6133 ( .A(n6766), .ZN(n6755) );
  AND2_X1 U6134 ( .A1(n6761), .A2(n6757), .ZN(n6756) );
  INV_X1 U6135 ( .A(\UUT/branch_rega [10]), .ZN(n6757) );
  INV_X1 U6136 ( .A(n6782), .ZN(n6758) );
  NAND2_X1 U6137 ( .A1(n6763), .A2(n6758), .ZN(n6759) );
  INV_X1 U6138 ( .A(n6824), .ZN(n6760) );
  NOR2_X2 U6139 ( .A1(n6767), .A2(n6760), .ZN(n6761) );
  INV_X1 U6140 ( .A(n6873), .ZN(n6762) );
  NOR2_X2 U6141 ( .A1(n6769), .A2(n6762), .ZN(n6763) );
  INV_X1 U6142 ( .A(\UUT/branch_rega [19]), .ZN(n6833) );
  INV_X1 U6143 ( .A(\UUT/branch_rega [19]), .ZN(n6891) );
  INV_X1 U6144 ( .A(n6796), .ZN(n6798) );
  INV_X1 U6145 ( .A(\UUT/branch_rega [19]), .ZN(n6879) );
  OR2_X1 U6146 ( .A1(\UUT/branch_rega [5]), .A2(n6765), .ZN(n6764) );
  INV_X1 U6147 ( .A(n6774), .ZN(n6765) );
  OR2_X1 U6148 ( .A1(n6771), .A2(n6768), .ZN(n6767) );
  INV_X4 U6149 ( .A(n6817), .ZN(n6768) );
  INV_X1 U6150 ( .A(n6853), .ZN(n6770) );
  NAND2_X1 U6151 ( .A1(n6772), .A2(n6826), .ZN(n6771) );
  NOR2_X1 U6152 ( .A1(n6786), .A2(n6778), .ZN(n6772) );
  INV_X1 U6153 ( .A(n6808), .ZN(n6773) );
  NOR2_X2 U6154 ( .A1(n6787), .A2(n6773), .ZN(n6774) );
  INV_X1 U6155 ( .A(\UUT/branch_rega [17]), .ZN(n6775) );
  NAND2_X1 U6156 ( .A1(n6781), .A2(n6775), .ZN(n6776) );
  INV_X1 U6157 ( .A(n6842), .ZN(n6778) );
  INV_X32 U6158 ( .A(\UUT/branch_rega [2]), .ZN(n6779) );
  INV_X1 U6159 ( .A(\UUT/branch_rega [24]), .ZN(n6877) );
  OAI222_X4 U6160 ( .A1(n5477), .A2(n5528), .B1(n5421), .B2(n6364), .C1(n5479), 
        .C2(n5530), .ZN(\UUT/branch_rega [24]) );
  INV_X1 U6161 ( .A(n6879), .ZN(n6780) );
  NOR2_X1 U6162 ( .A1(n6788), .A2(n6780), .ZN(n6781) );
  INV_X32 U6163 ( .A(n6846), .ZN(n6782) );
  INV_X32 U6164 ( .A(\UUT/branch_rega [6]), .ZN(n6783) );
  INV_X32 U6165 ( .A(n6835), .ZN(n6784) );
  NAND2_X1 U6166 ( .A1(n6789), .A2(n6790), .ZN(n6785) );
  OR2_X1 U6167 ( .A1(\UUT/branch_rega [22]), .A2(n6792), .ZN(n6786) );
  AND2_X1 U6168 ( .A1(n6791), .A2(n6854), .ZN(n6790) );
  INV_X1 U6169 ( .A(n6795), .ZN(n6791) );
  INV_X1 U6170 ( .A(n6798), .ZN(n6793) );
  INV_X32 U6171 ( .A(n6874), .ZN(n6795) );
  OR2_X1 U6172 ( .A1(\UUT/branch_rega [20]), .A2(n6797), .ZN(n6796) );
  INV_X1 U6173 ( .A(n6801), .ZN(n6797) );
  OR2_X1 U6174 ( .A1(n6800), .A2(\UUT/branch_rega [2]), .ZN(n6799) );
  INV_X1 U6175 ( .A(n6847), .ZN(n6800) );
  AND2_X1 U6176 ( .A1(n6834), .A2(n6833), .ZN(n6801) );
  INV_X4 U6177 ( .A(\UUT/branch_rega [1]), .ZN(n6847) );
  OR2_X1 U6178 ( .A1(\UUT/branch_rega [21]), .A2(\UUT/branch_rega [20]), .ZN(
        n6802) );
  OR2_X1 U6179 ( .A1(\UUT/branch_rega [9]), .A2(\UUT/branch_rega [8]), .ZN(
        n6804) );
  INV_X32 U6180 ( .A(n6804), .ZN(n6805) );
  INV_X1 U6181 ( .A(n6837), .ZN(n6806) );
  AND2_X1 U6182 ( .A1(n6810), .A2(n6816), .ZN(n6809) );
  INV_X1 U6183 ( .A(\UUT/branch_rega [23]), .ZN(n6810) );
  INV_X1 U6184 ( .A(n6815), .ZN(n6816) );
  INV_X1 U6185 ( .A(\UUT/branch_rega [28]), .ZN(n6837) );
  INV_X32 U6186 ( .A(\UUT/branch_rega [7]), .ZN(n6811) );
  INV_X32 U6187 ( .A(\UUT/branch_rega [11]), .ZN(n6812) );
  INV_X1 U6188 ( .A(\UUT/branch_rega [15]), .ZN(n6814) );
  OR2_X1 U6189 ( .A1(\UUT/branch_rega [25]), .A2(\UUT/branch_rega [24]), .ZN(
        n6815) );
  INV_X32 U6190 ( .A(\UUT/branch_rega [14]), .ZN(n6817) );
  INV_X32 U6191 ( .A(\UUT/branch_rega [10]), .ZN(n6818) );
  INV_X1 U6192 ( .A(\UUT/branch_rega [16]), .ZN(n6820) );
  INV_X32 U6193 ( .A(\UUT/branch_rega [23]), .ZN(n6821) );
  AND2_X2 U6194 ( .A1(n6871), .A2(n6872), .ZN(n6822) );
  INV_X1 U6195 ( .A(\UUT/branch_rega [17]), .ZN(n6823) );
  AND2_X1 U6196 ( .A1(n6825), .A2(n6866), .ZN(n6824) );
  INV_X1 U6197 ( .A(\UUT/branch_rega [11]), .ZN(n6825) );
  INV_X1 U6198 ( .A(\UUT/branch_rega [15]), .ZN(n6827) );
  INV_X1 U6199 ( .A(n6892), .ZN(n6828) );
  INV_X32 U6200 ( .A(\UUT/branch_rega [22]), .ZN(n6830) );
  INV_X32 U6201 ( .A(\UUT/branch_rega [3]), .ZN(n6835) );
  INV_X1 U6202 ( .A(\UUT/branch_rega [20]), .ZN(n6836) );
  INV_X4 U6203 ( .A(n6464), .ZN(n6839) );
  INV_X32 U6204 ( .A(n6839), .ZN(n6840) );
  INV_X32 U6205 ( .A(\UUT/branch_rega [17]), .ZN(n6842) );
  OR2_X1 U6206 ( .A1(n133), .A2(n861), .ZN(n6843) );
  OR2_X1 U6207 ( .A1(n5686), .A2(n135), .ZN(n6844) );
  OAI222_X4 U6208 ( .A1(n5471), .A2(n5528), .B1(n5419), .B2(n6364), .C1(n5473), 
        .C2(n5530), .ZN(\UUT/branch_rega [26]) );
  OAI222_X4 U6209 ( .A1(n5474), .A2(n5528), .B1(n5420), .B2(n6364), .C1(n5476), 
        .C2(n5530), .ZN(\UUT/branch_rega [25]) );
  INV_X32 U6210 ( .A(\UUT/branch_rega [14]), .ZN(n6846) );
  INV_X1 U6211 ( .A(n907), .ZN(n2324) );
  OR2_X1 U6212 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N124 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N125 ) );
  NAND2_X1 U6213 ( .A1(n6699), .A2(n6859), .ZN(n6850) );
  INV_X32 U6214 ( .A(\UUT/branch_rega [25]), .ZN(n6852) );
  INV_X1 U6215 ( .A(n6475), .ZN(n6861) );
  INV_X1 U6216 ( .A(n6489), .ZN(n6860) );
  NAND2_X1 U6217 ( .A1(n6862), .A2(n6863), .ZN(n6887) );
  AND2_X1 U6218 ( .A1(n6864), .A2(n6890), .ZN(n6863) );
  INV_X1 U6219 ( .A(n6889), .ZN(n6864) );
  INV_X32 U6220 ( .A(n6865), .ZN(n6866) );
  BUF_X1 U6221 ( .A(\UUT/Mpath/the_mult/Mult_out[0] ), .Z(n6869) );
  NOR2_X1 U6222 ( .A1(\UUT/branch_rega [30]), .A2(n6875), .ZN(n6870) );
  INV_X32 U6223 ( .A(\UUT/branch_rega [24]), .ZN(n6871) );
  INV_X32 U6224 ( .A(\UUT/branch_rega [15]), .ZN(n6873) );
  INV_X32 U6225 ( .A(\UUT/branch_rega [13]), .ZN(n6878) );
  INV_X32 U6226 ( .A(\UUT/branch_rega [13]), .ZN(n6880) );
  NAND2_X1 U6227 ( .A1(n6893), .A2(n6894), .ZN(n6881) );
  INV_X1 U6228 ( .A(n6881), .ZN(n6882) );
  NAND2_X2 U6229 ( .A1(n137), .A2(n948), .ZN(n6883) );
  INV_X32 U6230 ( .A(\UUT/branch_rega [18]), .ZN(n6884) );
  NAND2_X1 U6231 ( .A1(n6887), .A2(n6888), .ZN(n6296) );
  OR2_X1 U6232 ( .A1(n6295), .A2(n6861), .ZN(n6888) );
  OR2_X1 U6233 ( .A1(\UUT/branch_rega [0]), .A2(n6295), .ZN(n6889) );
  NOR2_X1 U6234 ( .A1(\UUT/branch_rega [2]), .A2(\UUT/branch_rega [1]), .ZN(
        n6890) );
  AOI21_X2 U6235 ( .B1(\UUT/Mcontrol/Nextpc_decoding/N32 ), .B2(
        \UUT/Mcontrol/Nextpc_decoding/N230 ), .A(
        \UUT/Mcontrol/Nextpc_decoding/N236 ), .ZN(n6299) );
  INV_X32 U6236 ( .A(\UUT/branch_rega [18]), .ZN(n6892) );
  INV_X1 U6237 ( .A(\UUT/branch_rega [31]), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N159 ) );
  OR2_X1 U6238 ( .A1(n133), .A2(n1142), .ZN(n6893) );
  OR2_X1 U6239 ( .A1(n5685), .A2(n135), .ZN(n6894) );
  BUF_X1 U6240 ( .A(\UUT/Mpath/out_regB[4] ), .Z(n6895) );
  BUF_X1 U6241 ( .A(\UUT/Mpath/out_regB[4] ), .Z(n6896) );
  BUF_X4 U6242 ( .A(\UUT/Mpath/out_regB[3] ), .Z(n6898) );
  INV_X1 U6243 ( .A(net54903), .ZN(net54843) );
  INV_X1 U6244 ( .A(net54903), .ZN(net54845) );
  INV_X1 U6245 ( .A(net54903), .ZN(net54847) );
  INV_X1 U6246 ( .A(net54903), .ZN(net54849) );
  INV_X1 U6247 ( .A(net54903), .ZN(net54851) );
  INV_X1 U6248 ( .A(net54953), .ZN(net54853) );
  INV_X1 U6249 ( .A(net54953), .ZN(net54855) );
  INV_X1 U6250 ( .A(net54953), .ZN(net54857) );
  INV_X1 U6251 ( .A(net54953), .ZN(net54859) );
  INV_X1 U6252 ( .A(net54953), .ZN(net54861) );
  INV_X1 U6253 ( .A(net54953), .ZN(net54863) );
  INV_X1 U6254 ( .A(net54953), .ZN(net54865) );
  INV_X1 U6255 ( .A(net54953), .ZN(net54867) );
  INV_X1 U6256 ( .A(net54953), .ZN(net54869) );
  INV_X1 U6257 ( .A(net54953), .ZN(net54871) );
  INV_X1 U6258 ( .A(net54953), .ZN(net54873) );
  INV_X1 U6259 ( .A(net54953), .ZN(net54875) );
  INV_X1 U6260 ( .A(net54953), .ZN(net54877) );
  INV_X1 U6261 ( .A(net54953), .ZN(net54879) );
  INV_X1 U6262 ( .A(net54953), .ZN(net54881) );
  INV_X1 U6263 ( .A(net54953), .ZN(net54883) );
  INV_X1 U6264 ( .A(net54953), .ZN(net54885) );
  INV_X1 U6265 ( .A(net54953), .ZN(net54887) );
  INV_X1 U6266 ( .A(net54953), .ZN(net54889) );
  INV_X1 U6267 ( .A(net54953), .ZN(net54891) );
  INV_X1 U6268 ( .A(net54953), .ZN(net54893) );
  INV_X1 U6269 ( .A(net54953), .ZN(net54895) );
  BUF_X4 U6270 ( .A(net54949), .Z(net54903) );
  BUF_X4 U6271 ( .A(net54949), .Z(net54905) );
  BUF_X4 U6272 ( .A(net54949), .Z(net54907) );
  BUF_X4 U6273 ( .A(net54947), .Z(net54909) );
  BUF_X4 U6274 ( .A(net54947), .Z(net54911) );
  BUF_X4 U6275 ( .A(net54947), .Z(net54913) );
  BUF_X4 U6276 ( .A(net54945), .Z(net54915) );
  BUF_X4 U6277 ( .A(net54945), .Z(net54917) );
  BUF_X4 U6278 ( .A(net54945), .Z(net54919) );
  BUF_X4 U6279 ( .A(net54943), .Z(net54921) );
  BUF_X4 U6280 ( .A(net54943), .Z(net54923) );
  BUF_X4 U6281 ( .A(net54943), .Z(net54925) );
  BUF_X4 U6282 ( .A(net54941), .Z(net54927) );
  BUF_X4 U6283 ( .A(net54941), .Z(net54929) );
  BUF_X4 U6284 ( .A(net54941), .Z(net54931) );
  BUF_X4 U6285 ( .A(net54939), .Z(net54933) );
  BUF_X4 U6286 ( .A(net54939), .Z(net54935) );
  BUF_X4 U6287 ( .A(net54939), .Z(net54937) );
  BUF_X4 U6288 ( .A(net54953), .Z(net54939) );
  BUF_X4 U6289 ( .A(net54953), .Z(net54941) );
  BUF_X4 U6290 ( .A(net54953), .Z(net54943) );
  BUF_X4 U6291 ( .A(net54953), .Z(net54945) );
  BUF_X4 U6292 ( .A(net54953), .Z(net54947) );
  BUF_X4 U6293 ( .A(net54953), .Z(net54949) );
  NAND4_X1 U6294 ( .A1(n6595), .A2(\localbus/c1_addr_outbus[30] ), .A3(
        \localbus/c1_addr_outbus[29] ), .A4(\localbus/c1_addr_outbus[28] ), 
        .ZN(\localbus/N61 ) );
  OAI21_X1 U6295 ( .B1(\localbus/c1_addr_outbus[29] ), .B2(
        \localbus/c1_addr_outbus[28] ), .A(\localbus/c1_addr_outbus[30] ), 
        .ZN(n6902) );
  INV_X1 U6296 ( .A(n6595), .ZN(n6901) );
  NAND2_X1 U6297 ( .A1(n6902), .A2(n6901), .ZN(\localbus/N60 ) );
  INV_X1 U6298 ( .A(n6903), .ZN(n6910) );
  OR2_X1 U6299 ( .A1(\localbus/c1_addr_outbus[14] ), .A2(
        \localbus/c1_addr_outbus[13] ), .ZN(n6904) );
  AOI221_X1 U6300 ( .B1(\localbus/c1_addr_outbus[16] ), .B2(
        \localbus/c1_addr_outbus[15] ), .C1(\localbus/c1_addr_outbus[16] ), 
        .C2(n6904), .A(n6910), .ZN(n6908) );
  NOR4_X1 U6301 ( .A1(\localbus/c1_addr_outbus[20] ), .A2(
        \localbus/c1_addr_outbus[19] ), .A3(\localbus/c1_addr_outbus[18] ), 
        .A4(\localbus/c1_addr_outbus[17] ), .ZN(n6907) );
  NOR4_X1 U6302 ( .A1(\localbus/c1_addr_outbus[24] ), .A2(
        \localbus/c1_addr_outbus[23] ), .A3(\localbus/c1_addr_outbus[22] ), 
        .A4(\localbus/c1_addr_outbus[21] ), .ZN(n6906) );
  NOR4_X1 U6303 ( .A1(\localbus/c1_addr_outbus[28] ), .A2(
        \localbus/c1_addr_outbus[27] ), .A3(\localbus/c1_addr_outbus[26] ), 
        .A4(\localbus/c1_addr_outbus[25] ), .ZN(n6905) );
  NOR2_X1 U6304 ( .A1(n6595), .A2(\localbus/c1_addr_outbus[30] ), .ZN(n6914)
         );
  NOR4_X1 U6305 ( .A1(\localbus/c1_addr_outbus[19] ), .A2(
        \localbus/c1_addr_outbus[18] ), .A3(\localbus/c1_addr_outbus[17] ), 
        .A4(\localbus/c1_addr_outbus[16] ), .ZN(n6912) );
  NOR4_X1 U6306 ( .A1(\localbus/c1_addr_outbus[23] ), .A2(
        \localbus/c1_addr_outbus[22] ), .A3(\localbus/c1_addr_outbus[21] ), 
        .A4(\localbus/c1_addr_outbus[20] ), .ZN(n6911) );
  AND2_X1 U6307 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  OAI22_X1 U6308 ( .A1(n6915), .A2(n6914), .B1(n6913), .B2(n6914), .ZN(
        \localbus/N55 ) );
  XNOR2_X1 U6309 ( .A(\UUT/Mcontrol/x_rd[0] ), .B(\UUT/rs2_addr [0]), .ZN(
        n6918) );
  XNOR2_X1 U6310 ( .A(\UUT/Mcontrol/x_rd[2] ), .B(\UUT/rs2_addr [2]), .ZN(
        n6917) );
  XNOR2_X1 U6311 ( .A(\UUT/Mcontrol/x_rd[1] ), .B(\UUT/rs2_addr [1]), .ZN(
        n6916) );
  NAND3_X1 U6312 ( .A1(n6918), .A2(n6917), .A3(n6916), .ZN(n6921) );
  XOR2_X1 U6313 ( .A(\UUT/Mcontrol/x_rd[3] ), .B(\UUT/rs2_addr [3]), .Z(n6920)
         );
  XOR2_X1 U6314 ( .A(\UUT/Mcontrol/x_rd[4] ), .B(\UUT/rs2_addr [4]), .Z(n6919)
         );
  NOR3_X1 U6315 ( .A1(n6921), .A2(n6920), .A3(n6919), .ZN(
        \UUT/Mcontrol/bp_logicB/N2 ) );
  XNOR2_X1 U6316 ( .A(\UUT/Mcontrol/m_sampled_xrd[0] ), .B(\UUT/rs2_addr [0]), 
        .ZN(n6924) );
  XNOR2_X1 U6317 ( .A(\UUT/Mcontrol/m_sampled_xrd[2] ), .B(\UUT/rs2_addr [2]), 
        .ZN(n6923) );
  XNOR2_X1 U6318 ( .A(\UUT/Mcontrol/m_sampled_xrd[1] ), .B(\UUT/rs2_addr [1]), 
        .ZN(n6922) );
  NAND3_X1 U6319 ( .A1(n6924), .A2(n6923), .A3(n6922), .ZN(n6927) );
  XOR2_X1 U6320 ( .A(\UUT/Mcontrol/m_sampled_xrd[3] ), .B(\UUT/rs2_addr [3]), 
        .Z(n6926) );
  XOR2_X1 U6321 ( .A(\UUT/Mcontrol/m_sampled_xrd[4] ), .B(\UUT/rs2_addr [4]), 
        .Z(n6925) );
  NOR3_X1 U6322 ( .A1(n6927), .A2(n6926), .A3(n6925), .ZN(
        \UUT/Mcontrol/bp_logicB/N3 ) );
  XNOR2_X1 U6323 ( .A(\UUT/Mcontrol/x_rd[0] ), .B(\UUT/rs1_addr [0]), .ZN(
        n6930) );
  XNOR2_X1 U6324 ( .A(\UUT/Mcontrol/x_rd[2] ), .B(\UUT/rs1_addr [2]), .ZN(
        n6929) );
  XNOR2_X1 U6325 ( .A(\UUT/Mcontrol/x_rd[1] ), .B(\UUT/rs1_addr [1]), .ZN(
        n6928) );
  NAND3_X1 U6326 ( .A1(n6930), .A2(n6929), .A3(n6928), .ZN(n6933) );
  XOR2_X1 U6327 ( .A(\UUT/Mcontrol/x_rd[3] ), .B(\UUT/rs1_addr [3]), .Z(n6932)
         );
  XOR2_X1 U6328 ( .A(\UUT/Mcontrol/x_rd[4] ), .B(\UUT/rs1_addr [4]), .Z(n6931)
         );
  NOR3_X1 U6329 ( .A1(n6933), .A2(n6932), .A3(n6931), .ZN(
        \UUT/Mcontrol/bp_logicA/N2 ) );
  XNOR2_X1 U6330 ( .A(\UUT/Mcontrol/m_sampled_xrd[0] ), .B(\UUT/rs1_addr [0]), 
        .ZN(n6936) );
  XNOR2_X1 U6331 ( .A(\UUT/Mcontrol/m_sampled_xrd[2] ), .B(\UUT/rs1_addr [2]), 
        .ZN(n6935) );
  XNOR2_X1 U6332 ( .A(\UUT/Mcontrol/m_sampled_xrd[1] ), .B(\UUT/rs1_addr [1]), 
        .ZN(n6934) );
  NAND3_X1 U6333 ( .A1(n6936), .A2(n6935), .A3(n6934), .ZN(n6939) );
  XOR2_X1 U6334 ( .A(\UUT/Mcontrol/m_sampled_xrd[3] ), .B(\UUT/rs1_addr [3]), 
        .Z(n6938) );
  XOR2_X1 U6335 ( .A(\UUT/Mcontrol/m_sampled_xrd[4] ), .B(\UUT/rs1_addr [4]), 
        .Z(n6937) );
  NOR3_X1 U6336 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(
        \UUT/Mcontrol/bp_logicA/N3 ) );
endmodule

