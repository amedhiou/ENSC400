---------------------------------------------------------------------------
--                      XI_memhandle.vhd                                 --
--                                                                       --
-- Created 2000 by F.M.Campi , fcampi@deis.unibo.it                      --
-- DEIS, Department of Electronics Informatics and Systems,              --
-- University of Bologna, BOLOGNA , ITALY                                -- 
---------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- "The contents of this file are subject to the Source Code Public License 
-- Version 1.0 (the "License"); you may not use this file except in compliance 
-- with the License. 
-- You may obtain a copy of the License at http://xirisc.deis.unibo.it/license.txt
--
-- Software distributed under the License is distributed on an "AS IS" basis, 
-- WITHOUT WARRANTY OF ANY KIND, either express or implied. 
-- See the License for the specific language governing rights and limitations
-- under the License.
--
-- This code was initially developed at "Department of electronics, computer 
-- science and Systems", (D.E.I.S.), University of Bologna, Bologna, Italy.
--
-- This license is a modification of the Cadence Design Systems Source Code Public 
-- License Version 1.0 which is similar to the Netscape public license.  
-- We believe this license conforms to requirements adopted by OpenSource.org.  
--
-- Please direct any comments regarding this license to xirisc@deis.unibo.it
-------------------------------------------------------------------------------

-- This vhdl block represents all the functionalities to master the XiRisc processor's
-- DATA memory bus cycle.
-- 


library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_arith.all;
  use work.menu.all;
  use work.basic.all;
  use work.components.all;


entity mem_handle is
  generic ( Word_Width      : positive := 32 );
  port ( clk,reset     : in  Std_logic;
         smdr_enable   : in  Std_logic;
         mem_baddr : in std_logic_vector(1 downto 0);
         -- The data to be stored => datapath in_regB signal
         stored_data   : in  std_logic_vector(word_width-1 downto 0);
         -- The data read from memory
         read_data     : out std_logic_vector(word_width-1 downto 0);
         -- Memory access control signals
         x_mem_command,m_mem_command   : in  mem_control;
         -- ddata_in bus
         data_in       : in  std_logic_vector(word_width-1 downto 0);
         -- ddata_out bus 
         data_out      : out std_logic_vector(word_width-1 downto 0)  );   
end mem_handle;


architecture STRUCTURAL of mem_handle is

  signal smdr_out : std_logic_vector(word_width-1 downto 0);
  
begin  -- STRUCTURAL


----------------------------------------------------------------------------
-- DATA HANDLE    logic                                                   --
----------------------------------------------------------------------------
    
  -- MEMORY STORE :In case a store operation is being executed,the value
  -- that is to be tranferred into dmemory is copied on the output data_bus port.
  --  
  -- Store_in_Memory_Data_Register: 
  -- This register is used to hold the data to be sent to external memory
  -- in case of STORE operations, that is specified by the rb source field
  -- of the instruction, bypassing the alu that is contemporaneusly used for
  -- the destination address calculation.

  SMDR: Data_Reg
     generic map ( init_value => 0, reg_width => word_width )
     port map ( clk,reset,smdr_enable,stored_data,smdr_out );
  
  store_output_reordering:process(smdr_out,x_mem_command)
  begin
    if x_mem_command.mb='0' then
      data_out <= smdr_out(7 downto 0) & smdr_out(7 downto 0) & smdr_out(7 downto 0) & smdr_out(7 downto 0);
    elsif x_mem_command.mh='0' then
      data_out <= smdr_out(15 downto 0) & smdr_out(15 downto 0);
    else
      data_out <= smdr_out;
    end if;
  end process;

  
  -- MEMORY LOAD:In case a load operation is being executed,the value that
  -- is being read is copied from the bidirectional data_bus.
  -- If this value is not 32-bits wide it is extended according to 
  -- the input signals control_logic generated by the control_logic.
  -- Note: Very recent Addition, fcampi@sfu.ca Jan 2013
  -- Based on the address, I am also choosing the approprite byte
  -- Before now, I assumed that was done on the outside!
  load_input_reorder_extension:
    process( data_in,mem_baddr,m_mem_command )
    begin
        if m_mem_command.sign = '0' and m_mem_command.mb = '0' then
          case mem_baddr is
            when "00" => read_data <= SXT(data_in(31 downto 24),word_width);
            when "01" => read_data <= SXT(data_in(23 downto 16),word_width);
            when "10" => read_data <= SXT(data_in(15 downto  8),word_width);
            when "11" => read_data <= SXT(data_in( 7 downto  0),word_width); 
            when others => read_data <= SXT(data_in(7 downto 0),word_width);
          end case;
        elsif m_mem_command.sign = '1' and m_mem_command.mb = '0' then
          case mem_baddr is
            when "00" => read_data <= EXT(data_in(31 downto 24),word_width);
            when "01" => read_data <= EXT(data_in(23 downto 16),word_width);
            when "10" => read_data <= EXT(data_in(15 downto  8),word_width);
            when "11" => read_data <= EXT(data_in( 7 downto  0),word_width); 
            when others => read_data <= EXT(data_in(7 downto 0),word_width);
          end case;
        elsif m_mem_command.sign = '0' and m_mem_command.mh = '0' then
          case mem_baddr(1) is
             when '0' => read_data <= SXT(data_in(31 downto 16),word_width);
             when '1' => read_data <= SXT(data_in(15 downto 0),word_width);
             when others => read_data <= SXT(data_in(15 downto 0),word_width);
          end case;
        elsif m_mem_command.sign = '1' and m_mem_command.mh = '0' then
          case mem_baddr(1) is
             when '0' => read_data <= EXT(data_in(31 downto 16),word_width);
             when '1' => read_data <= EXT(data_in(15 downto 0),word_width);
             when others => read_data <= ( others => '0');
          end case;
        else
              read_data <= data_in;         
        end if;
     end process;  

end STRUCTURAL;
