
module up_island_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96;

  XNOR2_X2 U41 ( .A(n82), .B(A[14]), .ZN(n39) );
  XNOR2_X1 U102 ( .A(n92), .B(A[4]), .ZN(n57) );
  INV_X1 U103 ( .A(B[30]), .ZN(n66) );
  INV_X1 U104 ( .A(B[31]), .ZN(n65) );
  NOR2_X1 U105 ( .A1(n11), .A2(n10), .ZN(n9) );
  BUF_X2 U106 ( .A(n1), .Z(NE) );
  INV_X1 U107 ( .A(B[2]), .ZN(n94) );
  INV_X1 U108 ( .A(B[8]), .ZN(n88) );
  XNOR2_X1 U109 ( .A(n88), .B(A[8]), .ZN(n49) );
  NOR2_X1 U110 ( .A1(n49), .A2(n48), .ZN(n47) );
  INV_X1 U111 ( .A(B[0]), .ZN(n96) );
  XNOR2_X1 U112 ( .A(n96), .B(A[0]), .ZN(n64) );
  NOR2_X1 U113 ( .A1(n64), .A2(n63), .ZN(n62) );
  XNOR2_X1 U114 ( .A(n78), .B(A[18]), .ZN(n31) );
  INV_X1 U115 ( .A(B[18]), .ZN(n78) );
  NOR2_X2 U116 ( .A1(n28), .A2(n21), .ZN(n3) );
  NOR2_X1 U117 ( .A1(n24), .A2(n23), .ZN(n22) );
  XNOR2_X1 U118 ( .A(n74), .B(A[22]), .ZN(n24) );
  INV_X1 U119 ( .A(B[22]), .ZN(n74) );
  INV_X1 U120 ( .A(B[5]), .ZN(n91) );
  XNOR2_X1 U121 ( .A(n70), .B(A[26]), .ZN(n17) );
  INV_X2 U122 ( .A(B[26]), .ZN(n70) );
  INV_X1 U123 ( .A(B[12]), .ZN(n84) );
  XNOR2_X1 U124 ( .A(n84), .B(A[12]), .ZN(n42) );
  NOR2_X1 U125 ( .A1(n42), .A2(n41), .ZN(n40) );
  XNOR2_X1 U126 ( .A(n72), .B(A[24]), .ZN(n20) );
  INV_X1 U127 ( .A(B[24]), .ZN(n72) );
  INV_X1 U128 ( .A(B[11]), .ZN(n85) );
  XNOR2_X1 U129 ( .A(n83), .B(A[13]), .ZN(n41) );
  INV_X1 U130 ( .A(B[13]), .ZN(n83) );
  NOR2_X1 U131 ( .A1(n58), .A2(n51), .ZN(n50) );
  NOR2_X1 U132 ( .A1(n54), .A2(n53), .ZN(n52) );
  XNOR2_X1 U133 ( .A(n89), .B(A[7]), .ZN(n53) );
  INV_X1 U134 ( .A(B[7]), .ZN(n89) );
  NAND2_X1 U135 ( .A1(n62), .A2(n59), .ZN(n58) );
  NOR2_X1 U136 ( .A1(n61), .A2(n60), .ZN(n59) );
  INV_X1 U137 ( .A(B[3]), .ZN(n93) );
  XNOR2_X1 U138 ( .A(n90), .B(A[6]), .ZN(n54) );
  INV_X1 U139 ( .A(B[6]), .ZN(n90) );
  CLKBUF_X1 U140 ( .A(n5), .Z(EQ) );
  NAND2_X1 U141 ( .A1(n3), .A2(n7), .ZN(n6) );
  XNOR2_X1 U142 ( .A(n75), .B(A[21]), .ZN(n26) );
  INV_X1 U143 ( .A(B[21]), .ZN(n75) );
  INV_X1 U144 ( .A(B[20]), .ZN(n76) );
  NAND2_X1 U145 ( .A1(n50), .A2(n35), .ZN(n2) );
  XNOR2_X1 U146 ( .A(n95), .B(A[1]), .ZN(n63) );
  INV_X1 U147 ( .A(B[1]), .ZN(n95) );
  NOR2_X1 U148 ( .A1(n34), .A2(n33), .ZN(n32) );
  INV_X1 U149 ( .A(B[16]), .ZN(n80) );
  NOR2_X2 U150 ( .A1(n4), .A2(n8), .ZN(n7) );
  NOR2_X1 U151 ( .A1(n17), .A2(n16), .ZN(n15) );
  XNOR2_X1 U152 ( .A(n69), .B(A[27]), .ZN(n16) );
  INV_X1 U153 ( .A(B[27]), .ZN(n69) );
  NOR2_X2 U154 ( .A1(n43), .A2(n36), .ZN(n35) );
  INV_X1 U155 ( .A(B[9]), .ZN(n87) );
  INV_X1 U156 ( .A(B[17]), .ZN(n79) );
  NOR2_X1 U157 ( .A1(n39), .A2(n38), .ZN(n37) );
  NAND2_X1 U158 ( .A1(n40), .A2(n37), .ZN(n36) );
  INV_X1 U159 ( .A(B[14]), .ZN(n82) );
  XNOR2_X1 U160 ( .A(n68), .B(A[28]), .ZN(n14) );
  NAND2_X1 U161 ( .A1(n25), .A2(n22), .ZN(n21) );
  NOR2_X2 U162 ( .A1(n27), .A2(n26), .ZN(n25) );
  XNOR2_X1 U163 ( .A(n76), .B(A[20]), .ZN(n27) );
  NOR2_X1 U164 ( .A1(n14), .A2(n13), .ZN(n12) );
  NAND2_X1 U165 ( .A1(n12), .A2(n9), .ZN(n8) );
  INV_X1 U166 ( .A(B[28]), .ZN(n68) );
  INV_X1 U167 ( .A(n5), .ZN(n1) );
  NOR2_X2 U168 ( .A1(n2), .A2(n6), .ZN(n5) );
  INV_X1 U169 ( .A(B[23]), .ZN(n73) );
  NAND2_X1 U170 ( .A1(n55), .A2(n52), .ZN(n51) );
  NOR2_X1 U171 ( .A1(n57), .A2(n56), .ZN(n55) );
  INV_X1 U172 ( .A(B[4]), .ZN(n92) );
  NAND2_X1 U173 ( .A1(n18), .A2(n15), .ZN(n4) );
  NOR2_X1 U174 ( .A1(n20), .A2(n19), .ZN(n18) );
  INV_X1 U175 ( .A(B[25]), .ZN(n71) );
  NAND2_X1 U176 ( .A1(n32), .A2(n29), .ZN(n28) );
  NOR2_X1 U177 ( .A1(n31), .A2(n30), .ZN(n29) );
  INV_X1 U178 ( .A(B[19]), .ZN(n77) );
  INV_X1 U179 ( .A(B[15]), .ZN(n81) );
  INV_X1 U180 ( .A(B[29]), .ZN(n67) );
  NAND2_X1 U181 ( .A1(n47), .A2(n44), .ZN(n43) );
  NOR2_X1 U182 ( .A1(n46), .A2(n45), .ZN(n44) );
  XNOR2_X1 U183 ( .A(n86), .B(A[10]), .ZN(n46) );
  INV_X1 U184 ( .A(B[10]), .ZN(n86) );
  XNOR2_X1 U185 ( .A(n94), .B(A[2]), .ZN(n61) );
  XNOR2_X1 U186 ( .A(n87), .B(A[9]), .ZN(n48) );
  XNOR2_X1 U187 ( .A(n71), .B(A[25]), .ZN(n19) );
  XNOR2_X1 U188 ( .A(n73), .B(A[23]), .ZN(n23) );
  XNOR2_X1 U189 ( .A(n81), .B(A[15]), .ZN(n38) );
  XNOR2_X1 U190 ( .A(n80), .B(A[16]), .ZN(n34) );
  XNOR2_X1 U191 ( .A(n91), .B(A[5]), .ZN(n56) );
  XNOR2_X1 U192 ( .A(n79), .B(A[17]), .ZN(n33) );
  XNOR2_X1 U193 ( .A(n77), .B(A[19]), .ZN(n30) );
  XNOR2_X1 U194 ( .A(n67), .B(A[29]), .ZN(n13) );
  XNOR2_X1 U195 ( .A(n66), .B(A[30]), .ZN(n11) );
  XNOR2_X1 U196 ( .A(n85), .B(A[11]), .ZN(n45) );
  XNOR2_X1 U197 ( .A(n93), .B(A[3]), .ZN(n60) );
  XNOR2_X1 U198 ( .A(n65), .B(A[31]), .ZN(n10) );
endmodule


module up_island_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  OAI21_X4 U1 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  AOI21_X4 U3 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  AOI21_X4 U7 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  OAI21_X4 U9 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U14 ( .A1(n22), .A2(n20), .ZN(n18) );
  OAI21_X4 U15 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  AOI21_X4 U21 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  NOR2_X4 U22 ( .A1(n28), .A2(n26), .ZN(n24) );
  OAI21_X4 U23 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U28 ( .A1(n34), .A2(n32), .ZN(n30) );
  OAI21_X4 U29 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NAND2_X4 U33 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  OAI21_X4 U35 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  NOR2_X4 U108 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  NAND2_X4 U109 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  NOR2_X4 U118 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X4 U119 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NAND2_X4 U120 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  NOR2_X1 U157 ( .A1(n151), .A2(B[31]), .ZN(n14) );
  NAND2_X1 U158 ( .A1(n151), .A2(B[31]), .ZN(n15) );
  INV_X1 U159 ( .A(A[29]), .ZN(n149) );
  INV_X4 U160 ( .A(A[0]), .ZN(n120) );
  INV_X4 U161 ( .A(A[2]), .ZN(n122) );
  INV_X1 U162 ( .A(A[14]), .ZN(n134) );
  INV_X1 U163 ( .A(A[13]), .ZN(n133) );
  INV_X1 U164 ( .A(A[15]), .ZN(n135) );
  OAI21_X1 U165 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X1 U166 ( .A1(n56), .A2(n54), .ZN(n52) );
  AOI21_X1 U167 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NAND2_X1 U168 ( .A1(n58), .A2(n52), .ZN(n50) );
  INV_X1 U169 ( .A(A[12]), .ZN(n132) );
  INV_X2 U170 ( .A(A[16]), .ZN(n136) );
  INV_X1 U171 ( .A(A[7]), .ZN(n127) );
  INV_X1 U172 ( .A(A[6]), .ZN(n126) );
  INV_X1 U173 ( .A(A[10]), .ZN(n130) );
  INV_X2 U174 ( .A(A[8]), .ZN(n128) );
  NAND2_X1 U175 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X1 U176 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  INV_X2 U177 ( .A(A[20]), .ZN(n140) );
  INV_X2 U178 ( .A(A[17]), .ZN(n137) );
  INV_X1 U179 ( .A(A[5]), .ZN(n125) );
  INV_X4 U180 ( .A(A[30]), .ZN(n150) );
  NAND2_X1 U181 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X1 U182 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  INV_X4 U183 ( .A(A[1]), .ZN(n121) );
  INV_X1 U184 ( .A(A[9]), .ZN(n129) );
  NAND2_X1 U185 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X1 U186 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  NAND2_X1 U187 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X1 U188 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  NAND2_X1 U189 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X1 U190 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NAND2_X1 U191 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X1 U192 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X1 U193 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X1 U194 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NOR2_X1 U195 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X1 U196 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  NAND2_X1 U197 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X1 U198 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  INV_X4 U199 ( .A(A[28]), .ZN(n148) );
  NAND2_X1 U200 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X1 U201 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NAND2_X1 U202 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  NOR2_X1 U203 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  INV_X4 U204 ( .A(A[3]), .ZN(n123) );
  INV_X4 U205 ( .A(A[4]), .ZN(n124) );
  INV_X4 U206 ( .A(A[26]), .ZN(n146) );
  INV_X4 U207 ( .A(A[27]), .ZN(n147) );
  NAND2_X1 U208 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X1 U209 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NAND2_X1 U210 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  NOR2_X1 U211 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X1 U212 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X1 U213 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NOR2_X1 U214 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X1 U215 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  NOR2_X1 U216 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X1 U217 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  INV_X4 U218 ( .A(A[23]), .ZN(n143) );
  INV_X4 U219 ( .A(A[22]), .ZN(n142) );
  INV_X4 U220 ( .A(A[24]), .ZN(n144) );
  INV_X4 U221 ( .A(A[25]), .ZN(n145) );
  INV_X4 U222 ( .A(A[31]), .ZN(n151) );
  INV_X4 U223 ( .A(A[19]), .ZN(n139) );
  INV_X4 U224 ( .A(A[21]), .ZN(n141) );
  INV_X2 U225 ( .A(A[18]), .ZN(n138) );
  INV_X4 U226 ( .A(A[11]), .ZN(n131) );
endmodule


module up_island_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  OAI21_X4 U1 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  AOI21_X4 U3 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  AOI21_X4 U7 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  OAI21_X4 U9 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U14 ( .A1(n22), .A2(n20), .ZN(n18) );
  OAI21_X4 U15 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  AOI21_X4 U21 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  NOR2_X4 U22 ( .A1(n28), .A2(n26), .ZN(n24) );
  OAI21_X4 U23 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U28 ( .A1(n34), .A2(n32), .ZN(n30) );
  OAI21_X4 U29 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NAND2_X4 U33 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  OAI21_X4 U35 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  NOR2_X4 U108 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  NAND2_X4 U109 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  NOR2_X4 U118 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X4 U119 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NAND2_X4 U120 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  INV_X1 U157 ( .A(B[31]), .ZN(n151) );
  INV_X1 U158 ( .A(A[29]), .ZN(n149) );
  INV_X4 U159 ( .A(A[0]), .ZN(n120) );
  INV_X4 U160 ( .A(A[2]), .ZN(n122) );
  INV_X1 U161 ( .A(A[14]), .ZN(n134) );
  INV_X1 U162 ( .A(A[13]), .ZN(n133) );
  INV_X1 U163 ( .A(A[15]), .ZN(n135) );
  OAI21_X1 U164 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X1 U165 ( .A1(n56), .A2(n54), .ZN(n52) );
  AOI21_X1 U166 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NAND2_X1 U167 ( .A1(n58), .A2(n52), .ZN(n50) );
  INV_X1 U168 ( .A(A[12]), .ZN(n132) );
  INV_X2 U169 ( .A(A[16]), .ZN(n136) );
  INV_X1 U170 ( .A(A[7]), .ZN(n127) );
  INV_X1 U171 ( .A(A[6]), .ZN(n126) );
  INV_X1 U172 ( .A(A[10]), .ZN(n130) );
  INV_X2 U173 ( .A(A[8]), .ZN(n128) );
  NAND2_X1 U174 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X1 U175 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  INV_X2 U176 ( .A(A[20]), .ZN(n140) );
  INV_X2 U177 ( .A(A[17]), .ZN(n137) );
  INV_X1 U178 ( .A(A[5]), .ZN(n125) );
  INV_X4 U179 ( .A(A[30]), .ZN(n150) );
  NAND2_X1 U180 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X1 U181 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  INV_X4 U182 ( .A(A[1]), .ZN(n121) );
  INV_X1 U183 ( .A(A[9]), .ZN(n129) );
  NAND2_X1 U184 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X1 U185 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  NAND2_X1 U186 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X1 U187 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  NAND2_X1 U188 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X1 U189 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NAND2_X1 U190 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X1 U191 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X1 U192 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X1 U193 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NOR2_X1 U194 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X1 U195 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  NAND2_X1 U196 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X1 U197 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  INV_X4 U198 ( .A(A[28]), .ZN(n148) );
  NAND2_X1 U199 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X1 U200 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NAND2_X1 U201 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  NOR2_X1 U202 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  INV_X4 U203 ( .A(A[3]), .ZN(n123) );
  INV_X4 U204 ( .A(A[4]), .ZN(n124) );
  INV_X4 U205 ( .A(A[26]), .ZN(n146) );
  INV_X4 U206 ( .A(A[27]), .ZN(n147) );
  NAND2_X1 U207 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X1 U208 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NAND2_X1 U209 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  NOR2_X1 U210 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X1 U211 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X1 U212 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NOR2_X1 U213 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X1 U214 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  NOR2_X1 U215 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X1 U216 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  INV_X4 U217 ( .A(A[23]), .ZN(n143) );
  INV_X4 U218 ( .A(A[22]), .ZN(n142) );
  INV_X4 U219 ( .A(A[24]), .ZN(n144) );
  INV_X4 U220 ( .A(A[25]), .ZN(n145) );
  NAND2_X1 U221 ( .A1(n151), .A2(A[31]), .ZN(n15) );
  NOR2_X1 U222 ( .A1(n151), .A2(A[31]), .ZN(n14) );
  INV_X4 U223 ( .A(A[19]), .ZN(n139) );
  INV_X4 U224 ( .A(A[21]), .ZN(n141) );
  INV_X2 U225 ( .A(A[18]), .ZN(n138) );
  INV_X4 U226 ( .A(A[11]), .ZN(n131) );
endmodule


module up_island_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636;

  NAND2_X1 U107 ( .A1(n1220), .A2(n1221), .ZN(B[8]) );
  NAND2_X1 U108 ( .A1(n1227), .A2(n1228), .ZN(B[7]) );
  NAND2_X1 U109 ( .A1(n1440), .A2(n1441), .ZN(B[22]) );
  NAND2_X1 U110 ( .A1(n1457), .A2(n1458), .ZN(B[21]) );
  NAND2_X1 U111 ( .A1(A[0]), .A2(n1178), .ZN(n1636) );
  NAND2_X1 U112 ( .A1(n1423), .A2(n1424), .ZN(B[23]) );
  NAND2_X1 U113 ( .A1(A[2]), .A2(n1175), .ZN(n1520) );
  INV_X1 U114 ( .A(A[2]), .ZN(n1634) );
  INV_X4 U115 ( .A(SH[2]), .ZN(n1183) );
  NAND2_X1 U116 ( .A1(A[1]), .A2(n1175), .ZN(n1534) );
  INV_X1 U117 ( .A(A[1]), .ZN(n1620) );
  NAND2_X1 U118 ( .A1(n1279), .A2(n1280), .ZN(B[31]) );
  NAND2_X1 U119 ( .A1(A[3]), .A2(n1176), .ZN(n1613) );
  INV_X1 U120 ( .A(A[3]), .ZN(n1605) );
  NAND2_X1 U121 ( .A1(A[4]), .A2(n1177), .ZN(n1626) );
  INV_X1 U122 ( .A(A[4]), .ZN(n1594) );
  INV_X1 U123 ( .A(A[26]), .ZN(n1387) );
  INV_X1 U124 ( .A(A[0]), .ZN(n1628) );
  INV_X1 U125 ( .A(A[27]), .ZN(n1370) );
  INV_X1 U126 ( .A(A[23]), .ZN(n1438) );
  INV_X1 U127 ( .A(A[22]), .ZN(n1455) );
  INV_X1 U128 ( .A(A[24]), .ZN(n1421) );
  INV_X1 U129 ( .A(A[25]), .ZN(n1404) );
  INV_X1 U130 ( .A(A[19]), .ZN(n1371) );
  INV_X1 U131 ( .A(A[21]), .ZN(n1472) );
  INV_X1 U132 ( .A(A[15]), .ZN(n1439) );
  INV_X1 U133 ( .A(A[18]), .ZN(n1388) );
  INV_X1 U134 ( .A(A[17]), .ZN(n1405) );
  INV_X1 U135 ( .A(A[13]), .ZN(n1473) );
  NAND2_X1 U136 ( .A1(A[7]), .A2(n1176), .ZN(n1614) );
  INV_X1 U137 ( .A(A[7]), .ZN(n1559) );
  INV_X1 U138 ( .A(A[11]), .ZN(n1504) );
  INV_X1 U139 ( .A(A[20]), .ZN(n1489) );
  INV_X1 U140 ( .A(A[16]), .ZN(n1422) );
  INV_X1 U141 ( .A(A[9]), .ZN(n1531) );
  INV_X1 U142 ( .A(A[12]), .ZN(n1490) );
  NAND2_X1 U143 ( .A1(A[6]), .A2(n1178), .ZN(n1632) );
  INV_X1 U144 ( .A(A[6]), .ZN(n1571) );
  INV_X1 U145 ( .A(A[14]), .ZN(n1456) );
  INV_X1 U146 ( .A(A[8]), .ZN(n1545) );
  INV_X1 U147 ( .A(A[10]), .ZN(n1517) );
  NAND2_X1 U148 ( .A1(A[5]), .A2(n1177), .ZN(n1618) );
  INV_X1 U149 ( .A(A[5]), .ZN(n1583) );
  INV_X1 U150 ( .A(n1172), .ZN(n1162) );
  INV_X1 U151 ( .A(n1172), .ZN(n1163) );
  INV_X1 U152 ( .A(n1172), .ZN(n1164) );
  INV_X1 U153 ( .A(n1172), .ZN(n1165) );
  INV_X1 U154 ( .A(n1171), .ZN(n1166) );
  CLKBUF_X3 U155 ( .A(SH[4]), .Z(n1167) );
  CLKBUF_X3 U156 ( .A(SH[4]), .Z(n1168) );
  CLKBUF_X3 U157 ( .A(SH[4]), .Z(n1169) );
  CLKBUF_X3 U158 ( .A(SH[4]), .Z(n1170) );
  CLKBUF_X3 U159 ( .A(SH[4]), .Z(n1171) );
  CLKBUF_X3 U160 ( .A(SH[4]), .Z(n1172) );
  INV_X1 U161 ( .A(n1179), .ZN(n1173) );
  INV_X1 U162 ( .A(n1179), .ZN(n1174) );
  INV_X1 U163 ( .A(SH[3]), .ZN(n1175) );
  INV_X1 U164 ( .A(SH[3]), .ZN(n1176) );
  INV_X1 U165 ( .A(SH[3]), .ZN(n1177) );
  INV_X1 U166 ( .A(SH[3]), .ZN(n1178) );
  INV_X1 U167 ( .A(SH[3]), .ZN(n1179) );
  INV_X1 U168 ( .A(n1183), .ZN(n1180) );
  INV_X1 U169 ( .A(n1183), .ZN(n1181) );
  INV_X1 U170 ( .A(n1183), .ZN(n1182) );
  INV_X1 U171 ( .A(n1189), .ZN(n1184) );
  INV_X1 U172 ( .A(n1188), .ZN(n1185) );
  INV_X1 U173 ( .A(n1189), .ZN(n1186) );
  INV_X1 U174 ( .A(n1188), .ZN(n1187) );
  INV_X2 U175 ( .A(SH[1]), .ZN(n1188) );
  INV_X2 U176 ( .A(SH[1]), .ZN(n1189) );
  INV_X1 U177 ( .A(n1196), .ZN(n1190) );
  INV_X1 U178 ( .A(n1199), .ZN(n1191) );
  INV_X1 U179 ( .A(n1200), .ZN(n1192) );
  INV_X1 U180 ( .A(n1201), .ZN(n1193) );
  INV_X1 U181 ( .A(n1202), .ZN(n1194) );
  CLKBUF_X3 U182 ( .A(SH[0]), .Z(n1195) );
  CLKBUF_X3 U183 ( .A(SH[0]), .Z(n1196) );
  CLKBUF_X3 U184 ( .A(SH[0]), .Z(n1197) );
  CLKBUF_X3 U185 ( .A(SH[0]), .Z(n1198) );
  CLKBUF_X3 U186 ( .A(SH[0]), .Z(n1199) );
  CLKBUF_X3 U187 ( .A(SH[0]), .Z(n1200) );
  CLKBUF_X3 U188 ( .A(SH[0]), .Z(n1201) );
  CLKBUF_X3 U189 ( .A(SH[0]), .Z(n1202) );
  CLKBUF_X3 U190 ( .A(SH[0]), .Z(n1203) );
  CLKBUF_X3 U191 ( .A(SH[0]), .Z(n1204) );
  CLKBUF_X3 U192 ( .A(SH[0]), .Z(n1205) );
  CLKBUF_X3 U193 ( .A(SH[0]), .Z(n1206) );
  CLKBUF_X3 U194 ( .A(SH[0]), .Z(n1207) );
  CLKBUF_X3 U195 ( .A(SH[0]), .Z(n1208) );
  CLKBUF_X3 U196 ( .A(SH[0]), .Z(n1209) );
  NAND2_X2 U197 ( .A1(n1210), .A2(n1211), .ZN(B[9]) );
  MUX2_X1 U198 ( .A(n1212), .B(n1213), .S(n1184), .Z(n1211) );
  NAND2_X2 U199 ( .A1(n1208), .A2(n1214), .ZN(n1213) );
  NAND2_X2 U200 ( .A1(n1209), .A2(n1215), .ZN(n1212) );
  MUX2_X1 U201 ( .A(n1216), .B(n1217), .S(n1187), .Z(n1210) );
  NAND2_X2 U202 ( .A1(n1218), .A2(n1192), .ZN(n1217) );
  NAND2_X2 U203 ( .A1(n1219), .A2(n1190), .ZN(n1216) );
  MUX2_X1 U204 ( .A(n1222), .B(n1223), .S(n1187), .Z(n1221) );
  NAND2_X2 U205 ( .A1(n1209), .A2(n1224), .ZN(n1223) );
  NAND2_X2 U206 ( .A1(n1208), .A2(n1218), .ZN(n1222) );
  MUX2_X1 U207 ( .A(n1225), .B(n1226), .S(n1187), .Z(n1220) );
  NAND2_X2 U208 ( .A1(n1214), .A2(n1190), .ZN(n1226) );
  NAND2_X2 U209 ( .A1(n1215), .A2(n1190), .ZN(n1225) );
  MUX2_X1 U210 ( .A(n1229), .B(n1230), .S(n1187), .Z(n1228) );
  NAND2_X2 U211 ( .A1(n1208), .A2(n1231), .ZN(n1230) );
  NAND2_X2 U212 ( .A1(n1207), .A2(n1214), .ZN(n1229) );
  MUX2_X1 U213 ( .A(n1232), .B(n1233), .S(n1187), .Z(n1227) );
  NAND2_X2 U214 ( .A1(n1224), .A2(n1190), .ZN(n1233) );
  NAND2_X2 U215 ( .A1(n1218), .A2(n1190), .ZN(n1232) );
  NAND2_X2 U216 ( .A1(n1234), .A2(n1235), .ZN(B[6]) );
  MUX2_X1 U217 ( .A(n1236), .B(n1237), .S(n1186), .Z(n1235) );
  NAND2_X2 U218 ( .A1(n1238), .A2(n1195), .ZN(n1237) );
  NAND2_X2 U219 ( .A1(n1208), .A2(n1224), .ZN(n1236) );
  MUX2_X1 U220 ( .A(n1239), .B(n1240), .S(n1186), .Z(n1234) );
  NAND2_X2 U221 ( .A1(n1231), .A2(n1190), .ZN(n1240) );
  NAND2_X2 U222 ( .A1(n1214), .A2(n1190), .ZN(n1239) );
  INV_X2 U223 ( .A(n1241), .ZN(n1214) );
  MUX2_X1 U224 ( .A(n1242), .B(n1243), .S(n1180), .Z(n1241) );
  NAND2_X2 U225 ( .A1(n1244), .A2(n1164), .ZN(n1243) );
  NAND2_X2 U226 ( .A1(n1245), .A2(n1162), .ZN(n1242) );
  NAND2_X2 U227 ( .A1(n1246), .A2(n1247), .ZN(B[5]) );
  MUX2_X1 U228 ( .A(n1248), .B(n1249), .S(n1186), .Z(n1247) );
  NAND2_X2 U229 ( .A1(n1250), .A2(n1195), .ZN(n1249) );
  NAND2_X2 U230 ( .A1(n1207), .A2(n1231), .ZN(n1248) );
  MUX2_X1 U231 ( .A(n1251), .B(n1252), .S(n1186), .Z(n1246) );
  NAND2_X2 U232 ( .A1(n1238), .A2(n1190), .ZN(n1252) );
  NAND2_X2 U233 ( .A1(n1224), .A2(n1190), .ZN(n1251) );
  INV_X2 U234 ( .A(n1253), .ZN(n1224) );
  MUX2_X1 U235 ( .A(n1254), .B(n1255), .S(n1182), .Z(n1253) );
  NAND2_X2 U236 ( .A1(n1256), .A2(n1162), .ZN(n1255) );
  NAND2_X2 U237 ( .A1(n1257), .A2(n1162), .ZN(n1254) );
  NAND2_X2 U238 ( .A1(n1258), .A2(n1259), .ZN(B[4]) );
  MUX2_X1 U239 ( .A(n1260), .B(n1261), .S(n1186), .Z(n1259) );
  NAND2_X2 U240 ( .A1(n1262), .A2(n1195), .ZN(n1261) );
  NAND2_X2 U241 ( .A1(n1238), .A2(n1196), .ZN(n1260) );
  MUX2_X1 U242 ( .A(n1263), .B(n1264), .S(n1186), .Z(n1258) );
  NAND2_X2 U243 ( .A1(n1250), .A2(n1190), .ZN(n1264) );
  NAND2_X2 U244 ( .A1(n1231), .A2(n1190), .ZN(n1263) );
  INV_X2 U245 ( .A(n1265), .ZN(n1231) );
  MUX2_X1 U246 ( .A(n1266), .B(n1267), .S(n1182), .Z(n1265) );
  NAND2_X2 U247 ( .A1(n1268), .A2(n1162), .ZN(n1267) );
  NAND2_X2 U248 ( .A1(n1269), .A2(n1162), .ZN(n1266) );
  NAND2_X2 U249 ( .A1(n1270), .A2(n1271), .ZN(B[3]) );
  MUX2_X1 U250 ( .A(n1272), .B(n1273), .S(n1186), .Z(n1271) );
  NAND2_X2 U251 ( .A1(n1274), .A2(n1196), .ZN(n1273) );
  NAND2_X2 U252 ( .A1(n1250), .A2(n1195), .ZN(n1272) );
  MUX2_X1 U253 ( .A(n1275), .B(n1276), .S(n1186), .Z(n1270) );
  NAND2_X2 U254 ( .A1(n1262), .A2(n1190), .ZN(n1276) );
  NAND2_X2 U255 ( .A1(n1238), .A2(n1191), .ZN(n1275) );
  INV_X2 U256 ( .A(n1277), .ZN(n1238) );
  NAND3_X1 U257 ( .A1(n1183), .A2(n1166), .A3(n1278), .ZN(n1277) );
  MUX2_X1 U258 ( .A(n1281), .B(n1282), .S(n1186), .Z(n1280) );
  NAND2_X2 U259 ( .A1(n1207), .A2(n1283), .ZN(n1282) );
  NAND2_X2 U260 ( .A1(n1207), .A2(n1284), .ZN(n1281) );
  MUX2_X1 U261 ( .A(n1285), .B(n1286), .S(n1186), .Z(n1279) );
  NAND2_X2 U262 ( .A1(n1287), .A2(n1191), .ZN(n1286) );
  OAI21_X2 U263 ( .B1(n1288), .B2(n1289), .A(n1194), .ZN(n1285) );
  MUX2_X1 U264 ( .A(n1290), .B(n1291), .S(n1182), .Z(n1289) );
  AND2_X2 U265 ( .A1(n1292), .A2(n1165), .ZN(n1291) );
  AND2_X2 U266 ( .A1(n1293), .A2(n1165), .ZN(n1290) );
  MUX2_X1 U267 ( .A(A[31]), .B(A[23]), .S(n1173), .Z(n1293) );
  MUX2_X1 U268 ( .A(n1294), .B(n1295), .S(n1182), .Z(n1288) );
  AND2_X2 U269 ( .A1(n1172), .A2(n1296), .ZN(n1295) );
  AND2_X2 U270 ( .A1(n1172), .A2(n1297), .ZN(n1294) );
  NAND2_X2 U271 ( .A1(n1298), .A2(n1299), .ZN(B[30]) );
  MUX2_X1 U272 ( .A(n1300), .B(n1301), .S(n1186), .Z(n1299) );
  NAND2_X2 U273 ( .A1(n1206), .A2(n1302), .ZN(n1301) );
  NAND2_X2 U274 ( .A1(n1206), .A2(n1287), .ZN(n1300) );
  MUX2_X1 U275 ( .A(n1303), .B(n1304), .S(n1186), .Z(n1298) );
  NAND2_X2 U276 ( .A1(n1283), .A2(n1191), .ZN(n1304) );
  NAND2_X2 U277 ( .A1(n1284), .A2(n1191), .ZN(n1303) );
  NAND2_X2 U278 ( .A1(n1305), .A2(n1306), .ZN(n1284) );
  MUX2_X1 U279 ( .A(n1307), .B(n1308), .S(n1182), .Z(n1306) );
  NAND2_X2 U280 ( .A1(n1171), .A2(n1309), .ZN(n1308) );
  NAND2_X2 U281 ( .A1(n1171), .A2(n1310), .ZN(n1307) );
  MUX2_X1 U282 ( .A(n1311), .B(n1312), .S(n1182), .Z(n1305) );
  NAND2_X2 U283 ( .A1(n1313), .A2(n1162), .ZN(n1312) );
  NAND2_X2 U284 ( .A1(n1314), .A2(n1162), .ZN(n1311) );
  MUX2_X1 U285 ( .A(A[30]), .B(A[22]), .S(n1173), .Z(n1314) );
  NAND2_X2 U286 ( .A1(n1315), .A2(n1316), .ZN(B[2]) );
  NAND3_X1 U287 ( .A1(n1194), .A2(n1189), .A3(n1250), .ZN(n1316) );
  INV_X2 U288 ( .A(n1317), .ZN(n1250) );
  NAND3_X1 U289 ( .A1(n1183), .A2(n1166), .A3(n1244), .ZN(n1317) );
  MUX2_X1 U290 ( .A(n1318), .B(n1319), .S(n1197), .Z(n1315) );
  NAND2_X2 U291 ( .A1(n1262), .A2(n1188), .ZN(n1319) );
  NAND2_X2 U292 ( .A1(n1274), .A2(n1184), .ZN(n1318) );
  NAND2_X2 U293 ( .A1(n1320), .A2(n1321), .ZN(B[29]) );
  MUX2_X1 U294 ( .A(n1322), .B(n1323), .S(n1186), .Z(n1321) );
  NAND2_X2 U295 ( .A1(n1206), .A2(n1324), .ZN(n1323) );
  NAND2_X2 U296 ( .A1(n1206), .A2(n1283), .ZN(n1322) );
  MUX2_X1 U297 ( .A(n1325), .B(n1326), .S(n1186), .Z(n1320) );
  NAND2_X2 U298 ( .A1(n1302), .A2(n1191), .ZN(n1326) );
  NAND2_X2 U299 ( .A1(n1287), .A2(n1191), .ZN(n1325) );
  NAND2_X2 U300 ( .A1(n1327), .A2(n1328), .ZN(n1287) );
  MUX2_X1 U301 ( .A(n1329), .B(n1330), .S(n1182), .Z(n1328) );
  NAND2_X2 U302 ( .A1(n1170), .A2(n1331), .ZN(n1330) );
  NAND2_X2 U303 ( .A1(n1170), .A2(n1332), .ZN(n1329) );
  MUX2_X1 U304 ( .A(n1333), .B(n1334), .S(n1182), .Z(n1327) );
  NAND2_X2 U305 ( .A1(n1335), .A2(n1162), .ZN(n1334) );
  NAND2_X2 U306 ( .A1(n1336), .A2(n1162), .ZN(n1333) );
  MUX2_X1 U307 ( .A(A[29]), .B(A[21]), .S(n1173), .Z(n1336) );
  NAND2_X2 U308 ( .A1(n1337), .A2(n1338), .ZN(B[28]) );
  MUX2_X1 U309 ( .A(n1339), .B(n1340), .S(n1186), .Z(n1338) );
  NAND2_X2 U310 ( .A1(n1205), .A2(n1341), .ZN(n1340) );
  NAND2_X2 U311 ( .A1(n1205), .A2(n1302), .ZN(n1339) );
  MUX2_X1 U312 ( .A(n1342), .B(n1343), .S(n1186), .Z(n1337) );
  NAND2_X2 U313 ( .A1(n1324), .A2(n1191), .ZN(n1343) );
  NAND2_X2 U314 ( .A1(n1283), .A2(n1191), .ZN(n1342) );
  NAND2_X2 U315 ( .A1(n1344), .A2(n1345), .ZN(n1283) );
  MUX2_X1 U316 ( .A(n1346), .B(n1347), .S(n1181), .Z(n1345) );
  NAND2_X2 U317 ( .A1(n1170), .A2(n1348), .ZN(n1347) );
  NAND2_X2 U318 ( .A1(n1170), .A2(n1349), .ZN(n1346) );
  MUX2_X1 U319 ( .A(n1350), .B(n1351), .S(n1181), .Z(n1344) );
  NAND2_X2 U320 ( .A1(n1352), .A2(n1162), .ZN(n1351) );
  NAND2_X2 U321 ( .A1(n1353), .A2(n1162), .ZN(n1350) );
  MUX2_X1 U322 ( .A(A[28]), .B(A[20]), .S(n1173), .Z(n1353) );
  NAND2_X2 U323 ( .A1(n1354), .A2(n1355), .ZN(B[27]) );
  MUX2_X1 U324 ( .A(n1356), .B(n1357), .S(n1186), .Z(n1355) );
  NAND2_X2 U325 ( .A1(n1205), .A2(n1358), .ZN(n1357) );
  NAND2_X2 U326 ( .A1(n1205), .A2(n1324), .ZN(n1356) );
  MUX2_X1 U327 ( .A(n1359), .B(n1360), .S(n1186), .Z(n1354) );
  NAND2_X2 U328 ( .A1(n1341), .A2(n1191), .ZN(n1360) );
  NAND2_X2 U329 ( .A1(n1302), .A2(n1191), .ZN(n1359) );
  NAND2_X2 U330 ( .A1(n1361), .A2(n1362), .ZN(n1302) );
  MUX2_X1 U331 ( .A(n1363), .B(n1364), .S(n1181), .Z(n1362) );
  NAND2_X2 U332 ( .A1(n1170), .A2(n1365), .ZN(n1364) );
  NAND2_X2 U333 ( .A1(n1169), .A2(n1296), .ZN(n1363) );
  MUX2_X1 U334 ( .A(n1366), .B(n1367), .S(n1181), .Z(n1361) );
  NAND2_X2 U335 ( .A1(n1368), .A2(n1162), .ZN(n1367) );
  NAND2_X2 U336 ( .A1(n1292), .A2(n1163), .ZN(n1366) );
  INV_X2 U337 ( .A(n1369), .ZN(n1292) );
  MUX2_X1 U338 ( .A(n1370), .B(n1371), .S(n1173), .Z(n1369) );
  NAND2_X2 U339 ( .A1(n1372), .A2(n1373), .ZN(B[26]) );
  MUX2_X1 U340 ( .A(n1374), .B(n1375), .S(n1185), .Z(n1373) );
  NAND2_X2 U341 ( .A1(n1204), .A2(n1376), .ZN(n1375) );
  NAND2_X2 U342 ( .A1(n1204), .A2(n1341), .ZN(n1374) );
  MUX2_X1 U343 ( .A(n1377), .B(n1378), .S(n1185), .Z(n1372) );
  NAND2_X2 U344 ( .A1(n1358), .A2(n1191), .ZN(n1378) );
  NAND2_X2 U345 ( .A1(n1324), .A2(n1191), .ZN(n1377) );
  NAND2_X2 U346 ( .A1(n1379), .A2(n1380), .ZN(n1324) );
  MUX2_X1 U347 ( .A(n1381), .B(n1382), .S(n1181), .Z(n1380) );
  NAND2_X2 U348 ( .A1(n1169), .A2(n1245), .ZN(n1382) );
  NAND2_X2 U349 ( .A1(n1169), .A2(n1309), .ZN(n1381) );
  MUX2_X1 U350 ( .A(n1383), .B(n1384), .S(n1181), .Z(n1379) );
  NAND2_X2 U351 ( .A1(n1385), .A2(n1163), .ZN(n1384) );
  NAND2_X2 U352 ( .A1(n1313), .A2(n1163), .ZN(n1383) );
  INV_X2 U353 ( .A(n1386), .ZN(n1313) );
  MUX2_X1 U354 ( .A(n1387), .B(n1388), .S(n1173), .Z(n1386) );
  NAND2_X2 U355 ( .A1(n1389), .A2(n1390), .ZN(B[25]) );
  MUX2_X1 U356 ( .A(n1391), .B(n1392), .S(n1185), .Z(n1390) );
  NAND2_X2 U357 ( .A1(n1204), .A2(n1393), .ZN(n1392) );
  NAND2_X2 U358 ( .A1(n1204), .A2(n1358), .ZN(n1391) );
  MUX2_X1 U359 ( .A(n1394), .B(n1395), .S(n1185), .Z(n1389) );
  NAND2_X2 U360 ( .A1(n1376), .A2(n1192), .ZN(n1395) );
  NAND2_X2 U361 ( .A1(n1341), .A2(n1192), .ZN(n1394) );
  NAND2_X2 U362 ( .A1(n1396), .A2(n1397), .ZN(n1341) );
  MUX2_X1 U363 ( .A(n1398), .B(n1399), .S(n1181), .Z(n1397) );
  NAND2_X2 U364 ( .A1(n1169), .A2(n1257), .ZN(n1399) );
  NAND2_X2 U365 ( .A1(n1169), .A2(n1331), .ZN(n1398) );
  MUX2_X1 U366 ( .A(n1400), .B(n1401), .S(n1181), .Z(n1396) );
  NAND2_X2 U367 ( .A1(n1402), .A2(n1163), .ZN(n1401) );
  NAND2_X2 U368 ( .A1(n1335), .A2(n1163), .ZN(n1400) );
  INV_X2 U369 ( .A(n1403), .ZN(n1335) );
  MUX2_X1 U370 ( .A(n1404), .B(n1405), .S(n1173), .Z(n1403) );
  NAND2_X2 U371 ( .A1(n1406), .A2(n1407), .ZN(B[24]) );
  MUX2_X1 U372 ( .A(n1408), .B(n1409), .S(n1185), .Z(n1407) );
  NAND2_X2 U373 ( .A1(n1203), .A2(n1410), .ZN(n1409) );
  NAND2_X2 U374 ( .A1(n1203), .A2(n1376), .ZN(n1408) );
  MUX2_X1 U375 ( .A(n1411), .B(n1412), .S(n1185), .Z(n1406) );
  NAND2_X2 U376 ( .A1(n1393), .A2(n1192), .ZN(n1412) );
  NAND2_X2 U377 ( .A1(n1358), .A2(n1192), .ZN(n1411) );
  NAND2_X2 U378 ( .A1(n1413), .A2(n1414), .ZN(n1358) );
  MUX2_X1 U379 ( .A(n1415), .B(n1416), .S(n1181), .Z(n1414) );
  NAND2_X2 U380 ( .A1(n1168), .A2(n1269), .ZN(n1416) );
  NAND2_X2 U381 ( .A1(n1168), .A2(n1348), .ZN(n1415) );
  MUX2_X1 U382 ( .A(n1417), .B(n1418), .S(n1181), .Z(n1413) );
  NAND2_X2 U383 ( .A1(n1419), .A2(n1163), .ZN(n1418) );
  NAND2_X2 U384 ( .A1(n1352), .A2(n1163), .ZN(n1417) );
  INV_X2 U385 ( .A(n1420), .ZN(n1352) );
  MUX2_X1 U386 ( .A(n1421), .B(n1422), .S(n1173), .Z(n1420) );
  MUX2_X1 U387 ( .A(n1425), .B(n1426), .S(n1185), .Z(n1424) );
  NAND2_X2 U388 ( .A1(n1203), .A2(n1427), .ZN(n1426) );
  NAND2_X2 U389 ( .A1(n1202), .A2(n1393), .ZN(n1425) );
  MUX2_X1 U390 ( .A(n1428), .B(n1429), .S(n1185), .Z(n1423) );
  NAND2_X2 U391 ( .A1(n1410), .A2(n1192), .ZN(n1429) );
  NAND2_X2 U392 ( .A1(n1376), .A2(n1192), .ZN(n1428) );
  NAND2_X2 U393 ( .A1(n1430), .A2(n1431), .ZN(n1376) );
  MUX2_X1 U394 ( .A(n1432), .B(n1433), .S(n1181), .Z(n1431) );
  NAND2_X2 U395 ( .A1(n1168), .A2(n1278), .ZN(n1433) );
  NAND2_X2 U396 ( .A1(n1168), .A2(n1365), .ZN(n1432) );
  MUX2_X1 U397 ( .A(n1434), .B(n1435), .S(n1181), .Z(n1430) );
  NAND2_X2 U398 ( .A1(n1436), .A2(n1163), .ZN(n1435) );
  NAND2_X2 U399 ( .A1(n1368), .A2(n1163), .ZN(n1434) );
  INV_X2 U400 ( .A(n1437), .ZN(n1368) );
  MUX2_X1 U401 ( .A(n1438), .B(n1439), .S(n1173), .Z(n1437) );
  MUX2_X1 U402 ( .A(n1442), .B(n1443), .S(n1185), .Z(n1441) );
  NAND2_X2 U403 ( .A1(n1202), .A2(n1444), .ZN(n1443) );
  NAND2_X2 U404 ( .A1(n1202), .A2(n1410), .ZN(n1442) );
  MUX2_X1 U405 ( .A(n1445), .B(n1446), .S(n1185), .Z(n1440) );
  NAND2_X2 U406 ( .A1(n1427), .A2(n1192), .ZN(n1446) );
  NAND2_X2 U407 ( .A1(n1393), .A2(n1192), .ZN(n1445) );
  NAND2_X2 U408 ( .A1(n1447), .A2(n1448), .ZN(n1393) );
  MUX2_X1 U409 ( .A(n1449), .B(n1450), .S(n1181), .Z(n1448) );
  NAND2_X2 U410 ( .A1(n1168), .A2(n1244), .ZN(n1450) );
  NAND2_X2 U411 ( .A1(n1167), .A2(n1245), .ZN(n1449) );
  MUX2_X1 U412 ( .A(n1451), .B(n1452), .S(n1181), .Z(n1447) );
  NAND2_X2 U413 ( .A1(n1453), .A2(n1163), .ZN(n1452) );
  NAND2_X2 U414 ( .A1(n1385), .A2(n1163), .ZN(n1451) );
  INV_X2 U415 ( .A(n1454), .ZN(n1385) );
  MUX2_X1 U416 ( .A(n1455), .B(n1456), .S(n1173), .Z(n1454) );
  MUX2_X1 U417 ( .A(n1459), .B(n1460), .S(n1185), .Z(n1458) );
  NAND2_X2 U418 ( .A1(n1202), .A2(n1461), .ZN(n1460) );
  NAND2_X2 U419 ( .A1(n1201), .A2(n1427), .ZN(n1459) );
  MUX2_X1 U420 ( .A(n1462), .B(n1463), .S(n1185), .Z(n1457) );
  NAND2_X2 U421 ( .A1(n1444), .A2(n1192), .ZN(n1463) );
  NAND2_X2 U422 ( .A1(n1410), .A2(n1192), .ZN(n1462) );
  NAND2_X2 U423 ( .A1(n1464), .A2(n1465), .ZN(n1410) );
  MUX2_X1 U424 ( .A(n1466), .B(n1467), .S(n1181), .Z(n1465) );
  NAND2_X2 U425 ( .A1(n1167), .A2(n1256), .ZN(n1467) );
  NAND2_X2 U426 ( .A1(n1167), .A2(n1257), .ZN(n1466) );
  MUX2_X1 U427 ( .A(n1468), .B(n1469), .S(n1181), .Z(n1464) );
  NAND2_X2 U428 ( .A1(n1470), .A2(n1163), .ZN(n1469) );
  NAND2_X2 U429 ( .A1(n1402), .A2(n1164), .ZN(n1468) );
  INV_X2 U430 ( .A(n1471), .ZN(n1402) );
  MUX2_X1 U431 ( .A(n1472), .B(n1473), .S(n1173), .Z(n1471) );
  NAND2_X2 U432 ( .A1(n1474), .A2(n1475), .ZN(B[20]) );
  MUX2_X1 U433 ( .A(n1476), .B(n1477), .S(n1185), .Z(n1475) );
  NAND2_X2 U434 ( .A1(n1201), .A2(n1478), .ZN(n1477) );
  NAND2_X2 U435 ( .A1(n1201), .A2(n1444), .ZN(n1476) );
  MUX2_X1 U436 ( .A(n1479), .B(n1480), .S(n1185), .Z(n1474) );
  NAND2_X2 U437 ( .A1(n1461), .A2(n1192), .ZN(n1480) );
  NAND2_X2 U438 ( .A1(n1427), .A2(n1193), .ZN(n1479) );
  NAND2_X2 U439 ( .A1(n1481), .A2(n1482), .ZN(n1427) );
  MUX2_X1 U440 ( .A(n1483), .B(n1484), .S(n1180), .Z(n1482) );
  NAND2_X2 U441 ( .A1(n1167), .A2(n1268), .ZN(n1484) );
  NAND2_X2 U442 ( .A1(n1167), .A2(n1269), .ZN(n1483) );
  MUX2_X1 U443 ( .A(n1485), .B(n1486), .S(n1180), .Z(n1481) );
  NAND2_X2 U444 ( .A1(n1487), .A2(n1164), .ZN(n1486) );
  NAND2_X2 U445 ( .A1(n1419), .A2(n1164), .ZN(n1485) );
  INV_X2 U446 ( .A(n1488), .ZN(n1419) );
  MUX2_X1 U447 ( .A(n1489), .B(n1490), .S(n1173), .Z(n1488) );
  MUX2_X1 U448 ( .A(n1491), .B(n1492), .S(n1198), .Z(B[1]) );
  AND2_X2 U449 ( .A1(n1274), .A2(n1188), .ZN(n1492) );
  AND2_X2 U450 ( .A1(n1262), .A2(n1188), .ZN(n1491) );
  INV_X2 U451 ( .A(n1493), .ZN(n1262) );
  NAND3_X1 U452 ( .A1(n1183), .A2(n1165), .A3(n1256), .ZN(n1493) );
  NAND2_X2 U453 ( .A1(n1494), .A2(n1495), .ZN(B[19]) );
  MUX2_X1 U454 ( .A(n1496), .B(n1497), .S(n1185), .Z(n1495) );
  NAND2_X2 U455 ( .A1(n1201), .A2(n1498), .ZN(n1497) );
  NAND2_X2 U456 ( .A1(n1200), .A2(n1461), .ZN(n1496) );
  MUX2_X1 U457 ( .A(n1499), .B(n1500), .S(n1185), .Z(n1494) );
  NAND2_X2 U458 ( .A1(n1478), .A2(n1193), .ZN(n1500) );
  NAND2_X2 U459 ( .A1(n1444), .A2(n1193), .ZN(n1499) );
  NAND2_X2 U460 ( .A1(n1501), .A2(n1502), .ZN(n1444) );
  NAND3_X1 U461 ( .A1(n1183), .A2(n1166), .A3(n1436), .ZN(n1502) );
  INV_X2 U462 ( .A(n1503), .ZN(n1436) );
  MUX2_X1 U463 ( .A(n1371), .B(n1504), .S(n1174), .Z(n1503) );
  MUX2_X1 U464 ( .A(n1505), .B(n1506), .S(n1171), .Z(n1501) );
  NAND2_X2 U465 ( .A1(n1278), .A2(n1183), .ZN(n1506) );
  NAND2_X2 U466 ( .A1(n1180), .A2(n1297), .ZN(n1505) );
  NAND2_X2 U467 ( .A1(n1507), .A2(n1508), .ZN(B[18]) );
  MUX2_X1 U468 ( .A(n1509), .B(n1510), .S(n1185), .Z(n1508) );
  NAND2_X2 U469 ( .A1(n1200), .A2(n1511), .ZN(n1510) );
  NAND2_X2 U470 ( .A1(n1200), .A2(n1478), .ZN(n1509) );
  MUX2_X1 U471 ( .A(n1512), .B(n1513), .S(n1184), .Z(n1507) );
  NAND2_X2 U472 ( .A1(n1498), .A2(n1193), .ZN(n1513) );
  NAND2_X2 U473 ( .A1(n1461), .A2(n1193), .ZN(n1512) );
  NAND2_X2 U474 ( .A1(n1514), .A2(n1515), .ZN(n1461) );
  NAND3_X1 U475 ( .A1(n1183), .A2(n1166), .A3(n1453), .ZN(n1515) );
  INV_X2 U476 ( .A(n1516), .ZN(n1453) );
  MUX2_X1 U477 ( .A(n1388), .B(n1517), .S(n1174), .Z(n1516) );
  MUX2_X1 U478 ( .A(n1518), .B(n1519), .S(n1171), .Z(n1514) );
  NAND2_X2 U479 ( .A1(n1244), .A2(n1183), .ZN(n1519) );
  INV_X2 U480 ( .A(n1520), .ZN(n1244) );
  NAND2_X2 U481 ( .A1(n1180), .A2(n1310), .ZN(n1518) );
  NAND2_X2 U482 ( .A1(n1521), .A2(n1522), .ZN(B[17]) );
  MUX2_X1 U483 ( .A(n1523), .B(n1524), .S(n1184), .Z(n1522) );
  NAND2_X2 U484 ( .A1(n1200), .A2(n1525), .ZN(n1524) );
  NAND2_X2 U485 ( .A1(n1199), .A2(n1498), .ZN(n1523) );
  MUX2_X1 U486 ( .A(n1526), .B(n1527), .S(n1184), .Z(n1521) );
  NAND2_X2 U487 ( .A1(n1511), .A2(n1193), .ZN(n1527) );
  NAND2_X2 U488 ( .A1(n1478), .A2(n1193), .ZN(n1526) );
  NAND2_X2 U489 ( .A1(n1528), .A2(n1529), .ZN(n1478) );
  NAND3_X1 U490 ( .A1(n1183), .A2(n1166), .A3(n1470), .ZN(n1529) );
  INV_X2 U491 ( .A(n1530), .ZN(n1470) );
  MUX2_X1 U492 ( .A(n1405), .B(n1531), .S(n1174), .Z(n1530) );
  MUX2_X1 U493 ( .A(n1532), .B(n1533), .S(n1171), .Z(n1528) );
  NAND2_X2 U494 ( .A1(n1256), .A2(n1183), .ZN(n1533) );
  INV_X2 U495 ( .A(n1534), .ZN(n1256) );
  NAND2_X2 U496 ( .A1(n1180), .A2(n1332), .ZN(n1532) );
  NAND2_X2 U497 ( .A1(n1535), .A2(n1536), .ZN(B[16]) );
  MUX2_X1 U498 ( .A(n1537), .B(n1538), .S(n1184), .Z(n1536) );
  NAND2_X2 U499 ( .A1(n1198), .A2(n1539), .ZN(n1538) );
  NAND2_X2 U500 ( .A1(n1198), .A2(n1511), .ZN(n1537) );
  MUX2_X1 U501 ( .A(n1540), .B(n1541), .S(n1184), .Z(n1535) );
  NAND2_X2 U502 ( .A1(n1525), .A2(n1193), .ZN(n1541) );
  NAND2_X2 U503 ( .A1(n1498), .A2(n1193), .ZN(n1540) );
  NAND2_X2 U504 ( .A1(n1542), .A2(n1543), .ZN(n1498) );
  NAND3_X1 U505 ( .A1(n1183), .A2(n1166), .A3(n1487), .ZN(n1543) );
  INV_X2 U506 ( .A(n1544), .ZN(n1487) );
  MUX2_X1 U507 ( .A(n1422), .B(n1545), .S(n1174), .Z(n1544) );
  MUX2_X1 U508 ( .A(n1546), .B(n1547), .S(n1171), .Z(n1542) );
  NAND2_X2 U509 ( .A1(n1268), .A2(n1183), .ZN(n1547) );
  NAND2_X2 U510 ( .A1(n1180), .A2(n1349), .ZN(n1546) );
  NAND2_X2 U511 ( .A1(n1548), .A2(n1549), .ZN(B[15]) );
  MUX2_X1 U512 ( .A(n1550), .B(n1551), .S(n1184), .Z(n1549) );
  NAND2_X2 U513 ( .A1(n1197), .A2(n1552), .ZN(n1551) );
  NAND2_X2 U514 ( .A1(n1199), .A2(n1525), .ZN(n1550) );
  MUX2_X1 U515 ( .A(n1553), .B(n1554), .S(n1184), .Z(n1548) );
  NAND2_X2 U516 ( .A1(n1539), .A2(n1193), .ZN(n1554) );
  NAND2_X2 U517 ( .A1(n1511), .A2(n1193), .ZN(n1553) );
  INV_X2 U518 ( .A(n1555), .ZN(n1511) );
  MUX2_X1 U519 ( .A(n1556), .B(n1557), .S(n1180), .Z(n1555) );
  NAND2_X2 U520 ( .A1(n1296), .A2(n1164), .ZN(n1557) );
  NAND2_X2 U521 ( .A1(n1297), .A2(n1164), .ZN(n1556) );
  INV_X2 U522 ( .A(n1558), .ZN(n1297) );
  MUX2_X1 U523 ( .A(n1439), .B(n1559), .S(n1174), .Z(n1558) );
  NAND2_X2 U524 ( .A1(n1560), .A2(n1561), .ZN(B[14]) );
  MUX2_X1 U525 ( .A(n1562), .B(n1563), .S(n1184), .Z(n1561) );
  NAND2_X2 U526 ( .A1(n1197), .A2(n1564), .ZN(n1563) );
  NAND2_X2 U527 ( .A1(n1199), .A2(n1539), .ZN(n1562) );
  MUX2_X1 U528 ( .A(n1565), .B(n1566), .S(n1184), .Z(n1560) );
  NAND2_X2 U529 ( .A1(n1552), .A2(n1194), .ZN(n1566) );
  NAND2_X2 U530 ( .A1(n1525), .A2(n1194), .ZN(n1565) );
  INV_X2 U531 ( .A(n1567), .ZN(n1525) );
  MUX2_X1 U532 ( .A(n1568), .B(n1569), .S(n1180), .Z(n1567) );
  NAND2_X2 U533 ( .A1(n1309), .A2(n1164), .ZN(n1569) );
  NAND2_X2 U534 ( .A1(n1310), .A2(n1164), .ZN(n1568) );
  INV_X2 U535 ( .A(n1570), .ZN(n1310) );
  MUX2_X1 U536 ( .A(n1456), .B(n1571), .S(n1174), .Z(n1570) );
  NAND2_X2 U537 ( .A1(n1572), .A2(n1573), .ZN(B[13]) );
  MUX2_X1 U538 ( .A(n1574), .B(n1575), .S(n1184), .Z(n1573) );
  NAND2_X2 U539 ( .A1(n1197), .A2(n1576), .ZN(n1575) );
  NAND2_X2 U540 ( .A1(n1198), .A2(n1552), .ZN(n1574) );
  MUX2_X1 U541 ( .A(n1577), .B(n1578), .S(n1184), .Z(n1572) );
  NAND2_X2 U542 ( .A1(n1564), .A2(n1194), .ZN(n1578) );
  NAND2_X2 U543 ( .A1(n1539), .A2(n1194), .ZN(n1577) );
  INV_X2 U544 ( .A(n1579), .ZN(n1539) );
  MUX2_X1 U545 ( .A(n1580), .B(n1581), .S(n1180), .Z(n1579) );
  NAND2_X2 U546 ( .A1(n1331), .A2(n1164), .ZN(n1581) );
  NAND2_X2 U547 ( .A1(n1332), .A2(n1165), .ZN(n1580) );
  INV_X2 U548 ( .A(n1582), .ZN(n1332) );
  MUX2_X1 U549 ( .A(n1473), .B(n1583), .S(n1174), .Z(n1582) );
  NAND2_X2 U550 ( .A1(n1584), .A2(n1585), .ZN(B[12]) );
  MUX2_X1 U551 ( .A(n1586), .B(n1587), .S(n1184), .Z(n1585) );
  NAND2_X2 U552 ( .A1(n1197), .A2(n1219), .ZN(n1587) );
  NAND2_X2 U553 ( .A1(n1199), .A2(n1564), .ZN(n1586) );
  MUX2_X1 U554 ( .A(n1588), .B(n1589), .S(n1184), .Z(n1584) );
  NAND2_X2 U555 ( .A1(n1576), .A2(n1193), .ZN(n1589) );
  NAND2_X2 U556 ( .A1(n1552), .A2(n1194), .ZN(n1588) );
  INV_X2 U557 ( .A(n1590), .ZN(n1552) );
  MUX2_X1 U558 ( .A(n1591), .B(n1592), .S(n1180), .Z(n1590) );
  NAND2_X2 U559 ( .A1(n1348), .A2(n1164), .ZN(n1592) );
  NAND2_X2 U560 ( .A1(n1349), .A2(n1164), .ZN(n1591) );
  INV_X2 U561 ( .A(n1593), .ZN(n1349) );
  MUX2_X1 U562 ( .A(n1490), .B(n1594), .S(n1174), .Z(n1593) );
  NAND2_X2 U563 ( .A1(n1595), .A2(n1596), .ZN(B[11]) );
  MUX2_X1 U564 ( .A(n1597), .B(n1598), .S(n1184), .Z(n1596) );
  NAND2_X2 U565 ( .A1(n1196), .A2(n1215), .ZN(n1598) );
  NAND2_X2 U566 ( .A1(n1198), .A2(n1576), .ZN(n1597) );
  MUX2_X1 U567 ( .A(n1599), .B(n1600), .S(n1184), .Z(n1595) );
  NAND2_X2 U568 ( .A1(n1219), .A2(n1194), .ZN(n1600) );
  NAND2_X2 U569 ( .A1(n1564), .A2(n1194), .ZN(n1599) );
  INV_X2 U570 ( .A(n1601), .ZN(n1564) );
  MUX2_X1 U571 ( .A(n1602), .B(n1603), .S(n1180), .Z(n1601) );
  NAND2_X2 U572 ( .A1(n1365), .A2(n1165), .ZN(n1603) );
  NAND2_X2 U573 ( .A1(n1296), .A2(n1164), .ZN(n1602) );
  INV_X2 U574 ( .A(n1604), .ZN(n1296) );
  MUX2_X1 U575 ( .A(n1504), .B(n1605), .S(n1174), .Z(n1604) );
  NAND2_X2 U576 ( .A1(n1606), .A2(n1607), .ZN(B[10]) );
  MUX2_X1 U577 ( .A(n1608), .B(n1609), .S(n1184), .Z(n1607) );
  NAND2_X2 U578 ( .A1(n1196), .A2(n1218), .ZN(n1609) );
  INV_X2 U579 ( .A(n1610), .ZN(n1218) );
  MUX2_X1 U580 ( .A(n1611), .B(n1612), .S(n1180), .Z(n1610) );
  NAND2_X2 U581 ( .A1(n1278), .A2(n1165), .ZN(n1612) );
  INV_X2 U582 ( .A(n1613), .ZN(n1278) );
  NAND2_X2 U583 ( .A1(n1365), .A2(n1165), .ZN(n1611) );
  INV_X2 U584 ( .A(n1614), .ZN(n1365) );
  NAND2_X2 U585 ( .A1(n1203), .A2(n1219), .ZN(n1608) );
  INV_X2 U586 ( .A(n1615), .ZN(n1219) );
  MUX2_X1 U587 ( .A(n1616), .B(n1617), .S(n1180), .Z(n1615) );
  NAND2_X2 U588 ( .A1(n1257), .A2(n1165), .ZN(n1617) );
  INV_X2 U589 ( .A(n1618), .ZN(n1257) );
  NAND2_X2 U590 ( .A1(n1331), .A2(n1165), .ZN(n1616) );
  INV_X2 U591 ( .A(n1619), .ZN(n1331) );
  MUX2_X1 U592 ( .A(n1531), .B(n1620), .S(n1174), .Z(n1619) );
  MUX2_X1 U593 ( .A(n1621), .B(n1622), .S(n1185), .Z(n1606) );
  NAND2_X2 U594 ( .A1(n1215), .A2(n1194), .ZN(n1622) );
  INV_X2 U595 ( .A(n1623), .ZN(n1215) );
  MUX2_X1 U596 ( .A(n1624), .B(n1625), .S(n1180), .Z(n1623) );
  NAND2_X2 U597 ( .A1(n1269), .A2(n1165), .ZN(n1625) );
  INV_X2 U598 ( .A(n1626), .ZN(n1269) );
  NAND2_X2 U599 ( .A1(n1348), .A2(n1165), .ZN(n1624) );
  INV_X2 U600 ( .A(n1627), .ZN(n1348) );
  MUX2_X1 U601 ( .A(n1545), .B(n1628), .S(n1174), .Z(n1627) );
  NAND2_X2 U602 ( .A1(n1576), .A2(n1194), .ZN(n1621) );
  INV_X2 U603 ( .A(n1629), .ZN(n1576) );
  MUX2_X1 U604 ( .A(n1630), .B(n1631), .S(n1181), .Z(n1629) );
  NAND2_X2 U605 ( .A1(n1245), .A2(n1165), .ZN(n1631) );
  INV_X2 U606 ( .A(n1632), .ZN(n1245) );
  NAND2_X2 U607 ( .A1(n1309), .A2(n1165), .ZN(n1630) );
  INV_X2 U608 ( .A(n1633), .ZN(n1309) );
  MUX2_X1 U609 ( .A(n1517), .B(n1634), .S(n1174), .Z(n1633) );
  AND3_X2 U610 ( .A1(n1194), .A2(n1189), .A3(n1274), .ZN(B[0]) );
  INV_X2 U611 ( .A(n1635), .ZN(n1274) );
  NAND3_X1 U612 ( .A1(n1183), .A2(n1166), .A3(n1268), .ZN(n1635) );
  INV_X2 U613 ( .A(n1636), .ZN(n1268) );
endmodule


module up_island_DW01_bsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671;

  INV_X1 U169 ( .A(A[29]), .ZN(n1611) );
  NAND2_X1 U170 ( .A1(n1393), .A2(n1394), .ZN(B[21]) );
  NAND2_X1 U171 ( .A1(n1367), .A2(n1368), .ZN(B[23]) );
  INV_X1 U172 ( .A(A[2]), .ZN(n1460) );
  INV_X1 U173 ( .A(A[30]), .ZN(n1623) );
  INV_X1 U174 ( .A(A[1]), .ZN(n1479) );
  INV_X1 U175 ( .A(A[28]), .ZN(n1591) );
  INV_X1 U176 ( .A(A[3]), .ZN(n1572) );
  INV_X1 U177 ( .A(A[4]), .ZN(n1590) );
  INV_X1 U178 ( .A(A[26]), .ZN(n1461) );
  INV_X1 U179 ( .A(A[0]), .ZN(n1599) );
  INV_X1 U180 ( .A(A[27]), .ZN(n1573) );
  INV_X1 U181 ( .A(A[23]), .ZN(n1577) );
  INV_X1 U182 ( .A(A[22]), .ZN(n1619) );
  INV_X1 U183 ( .A(A[24]), .ZN(n1595) );
  INV_X1 U184 ( .A(A[25]), .ZN(n1480) );
  INV_X1 U185 ( .A(A[31]), .ZN(n1581) );
  INV_X1 U186 ( .A(A[19]), .ZN(n1569) );
  INV_X1 U187 ( .A(A[21]), .ZN(n1607) );
  INV_X1 U188 ( .A(A[15]), .ZN(n1578) );
  INV_X1 U189 ( .A(A[18]), .ZN(n1463) );
  INV_X1 U190 ( .A(A[17]), .ZN(n1482) );
  INV_X1 U191 ( .A(A[13]), .ZN(n1608) );
  INV_X1 U192 ( .A(A[7]), .ZN(n1580) );
  INV_X1 U193 ( .A(A[11]), .ZN(n1570) );
  INV_X1 U194 ( .A(A[20]), .ZN(n1587) );
  INV_X1 U195 ( .A(A[16]), .ZN(n1596) );
  INV_X1 U196 ( .A(A[9]), .ZN(n1483) );
  INV_X1 U197 ( .A(A[12]), .ZN(n1588) );
  INV_X1 U198 ( .A(A[6]), .ZN(n1622) );
  INV_X1 U199 ( .A(A[14]), .ZN(n1620) );
  INV_X1 U200 ( .A(A[8]), .ZN(n1598) );
  INV_X1 U201 ( .A(A[10]), .ZN(n1464) );
  INV_X1 U202 ( .A(A[5]), .ZN(n1610) );
  CLKBUF_X3 U203 ( .A(SH[4]), .Z(n1105) );
  CLKBUF_X3 U204 ( .A(SH[4]), .Z(n1106) );
  CLKBUF_X3 U205 ( .A(SH[4]), .Z(n1107) );
  CLKBUF_X3 U206 ( .A(SH[4]), .Z(n1108) );
  CLKBUF_X3 U207 ( .A(SH[4]), .Z(n1109) );
  CLKBUF_X3 U208 ( .A(SH[4]), .Z(n1110) );
  CLKBUF_X3 U209 ( .A(SH[3]), .Z(n1111) );
  CLKBUF_X3 U210 ( .A(SH[3]), .Z(n1112) );
  CLKBUF_X3 U211 ( .A(SH[3]), .Z(n1113) );
  INV_X1 U212 ( .A(n1132), .ZN(n1114) );
  INV_X1 U213 ( .A(n1132), .ZN(n1115) );
  INV_X1 U214 ( .A(n1133), .ZN(n1116) );
  INV_X1 U215 ( .A(n1133), .ZN(n1117) );
  INV_X1 U216 ( .A(n1133), .ZN(n1118) );
  INV_X1 U217 ( .A(n1133), .ZN(n1119) );
  CLKBUF_X3 U218 ( .A(SH[2]), .Z(n1120) );
  CLKBUF_X3 U219 ( .A(SH[2]), .Z(n1121) );
  CLKBUF_X3 U220 ( .A(SH[2]), .Z(n1122) );
  CLKBUF_X3 U221 ( .A(SH[2]), .Z(n1123) );
  CLKBUF_X3 U222 ( .A(SH[2]), .Z(n1124) );
  CLKBUF_X3 U223 ( .A(SH[2]), .Z(n1125) );
  CLKBUF_X3 U224 ( .A(SH[2]), .Z(n1126) );
  CLKBUF_X3 U225 ( .A(SH[2]), .Z(n1127) );
  CLKBUF_X3 U226 ( .A(SH[2]), .Z(n1128) );
  CLKBUF_X3 U227 ( .A(SH[2]), .Z(n1129) );
  CLKBUF_X3 U228 ( .A(SH[2]), .Z(n1130) );
  CLKBUF_X3 U229 ( .A(SH[2]), .Z(n1131) );
  CLKBUF_X3 U230 ( .A(SH[2]), .Z(n1132) );
  CLKBUF_X3 U231 ( .A(SH[2]), .Z(n1133) );
  INV_X1 U232 ( .A(n1152), .ZN(n1134) );
  INV_X1 U233 ( .A(n1152), .ZN(n1135) );
  INV_X1 U234 ( .A(n1153), .ZN(n1136) );
  INV_X1 U235 ( .A(n1153), .ZN(n1137) );
  INV_X1 U236 ( .A(n1153), .ZN(n1138) );
  INV_X1 U237 ( .A(n1153), .ZN(n1139) );
  CLKBUF_X3 U238 ( .A(SH[1]), .Z(n1140) );
  CLKBUF_X3 U239 ( .A(SH[1]), .Z(n1141) );
  CLKBUF_X3 U240 ( .A(SH[1]), .Z(n1142) );
  CLKBUF_X3 U241 ( .A(SH[1]), .Z(n1143) );
  CLKBUF_X3 U242 ( .A(SH[1]), .Z(n1144) );
  CLKBUF_X3 U243 ( .A(SH[1]), .Z(n1145) );
  CLKBUF_X3 U244 ( .A(SH[1]), .Z(n1146) );
  CLKBUF_X3 U245 ( .A(SH[1]), .Z(n1147) );
  CLKBUF_X3 U246 ( .A(SH[1]), .Z(n1148) );
  CLKBUF_X3 U247 ( .A(SH[1]), .Z(n1149) );
  CLKBUF_X3 U248 ( .A(SH[1]), .Z(n1150) );
  CLKBUF_X3 U249 ( .A(SH[1]), .Z(n1151) );
  CLKBUF_X3 U250 ( .A(SH[1]), .Z(n1152) );
  CLKBUF_X3 U251 ( .A(SH[1]), .Z(n1153) );
  CLKBUF_X3 U252 ( .A(SH[0]), .Z(n1154) );
  CLKBUF_X3 U253 ( .A(SH[0]), .Z(n1155) );
  CLKBUF_X3 U254 ( .A(SH[0]), .Z(n1156) );
  CLKBUF_X3 U255 ( .A(SH[0]), .Z(n1157) );
  CLKBUF_X3 U256 ( .A(SH[0]), .Z(n1158) );
  CLKBUF_X3 U257 ( .A(SH[0]), .Z(n1159) );
  NAND2_X2 U258 ( .A1(n1160), .A2(n1161), .ZN(B[9]) );
  MUX2_X1 U259 ( .A(n1162), .B(n1163), .S(n1154), .Z(n1161) );
  NAND2_X2 U260 ( .A1(n1152), .A2(n1164), .ZN(n1163) );
  NAND2_X2 U261 ( .A1(n1152), .A2(n1165), .ZN(n1162) );
  MUX2_X1 U262 ( .A(n1166), .B(n1167), .S(n1154), .Z(n1160) );
  NAND2_X2 U263 ( .A1(n1168), .A2(n1139), .ZN(n1167) );
  NAND2_X2 U264 ( .A1(n1169), .A2(n1139), .ZN(n1166) );
  NAND2_X2 U265 ( .A1(n1170), .A2(n1171), .ZN(B[8]) );
  MUX2_X1 U266 ( .A(n1172), .B(n1173), .S(n1154), .Z(n1171) );
  NAND2_X2 U267 ( .A1(n1152), .A2(n1174), .ZN(n1173) );
  NAND2_X2 U268 ( .A1(n1152), .A2(n1164), .ZN(n1172) );
  MUX2_X1 U269 ( .A(n1175), .B(n1176), .S(n1154), .Z(n1170) );
  NAND2_X2 U270 ( .A1(n1165), .A2(n1139), .ZN(n1176) );
  NAND2_X2 U271 ( .A1(n1168), .A2(n1139), .ZN(n1175) );
  NAND2_X2 U272 ( .A1(n1177), .A2(n1178), .ZN(B[7]) );
  MUX2_X1 U273 ( .A(n1179), .B(n1180), .S(n1154), .Z(n1178) );
  NAND2_X2 U274 ( .A1(n1151), .A2(n1181), .ZN(n1180) );
  NAND2_X2 U275 ( .A1(n1151), .A2(n1174), .ZN(n1179) );
  MUX2_X1 U276 ( .A(n1182), .B(n1183), .S(n1154), .Z(n1177) );
  NAND2_X2 U277 ( .A1(n1164), .A2(n1138), .ZN(n1183) );
  NAND2_X2 U278 ( .A1(n1165), .A2(n1138), .ZN(n1182) );
  NAND2_X2 U279 ( .A1(n1184), .A2(n1185), .ZN(B[6]) );
  MUX2_X1 U280 ( .A(n1186), .B(n1187), .S(n1154), .Z(n1185) );
  NAND2_X2 U281 ( .A1(n1151), .A2(n1188), .ZN(n1187) );
  NAND2_X2 U282 ( .A1(n1151), .A2(n1181), .ZN(n1186) );
  MUX2_X1 U283 ( .A(n1189), .B(n1190), .S(n1154), .Z(n1184) );
  NAND2_X2 U284 ( .A1(n1174), .A2(n1138), .ZN(n1190) );
  NAND2_X2 U285 ( .A1(n1164), .A2(n1138), .ZN(n1189) );
  NAND2_X2 U286 ( .A1(n1191), .A2(n1192), .ZN(n1164) );
  MUX2_X1 U287 ( .A(n1193), .B(n1194), .S(n1105), .Z(n1192) );
  NAND2_X2 U288 ( .A1(n1132), .A2(n1195), .ZN(n1194) );
  NAND2_X2 U289 ( .A1(n1132), .A2(n1196), .ZN(n1193) );
  MUX2_X1 U290 ( .A(n1197), .B(n1198), .S(n1105), .Z(n1191) );
  NAND2_X2 U291 ( .A1(n1199), .A2(n1119), .ZN(n1198) );
  NAND2_X2 U292 ( .A1(n1200), .A2(n1119), .ZN(n1197) );
  NAND2_X2 U293 ( .A1(n1201), .A2(n1202), .ZN(B[5]) );
  MUX2_X1 U294 ( .A(n1203), .B(n1204), .S(n1154), .Z(n1202) );
  NAND2_X2 U295 ( .A1(n1151), .A2(n1205), .ZN(n1204) );
  NAND2_X2 U296 ( .A1(n1150), .A2(n1188), .ZN(n1203) );
  MUX2_X1 U297 ( .A(n1206), .B(n1207), .S(n1154), .Z(n1201) );
  NAND2_X2 U298 ( .A1(n1181), .A2(n1138), .ZN(n1207) );
  NAND2_X2 U299 ( .A1(n1174), .A2(n1138), .ZN(n1206) );
  NAND2_X2 U300 ( .A1(n1208), .A2(n1209), .ZN(n1174) );
  MUX2_X1 U301 ( .A(n1210), .B(n1211), .S(n1105), .Z(n1209) );
  NAND2_X2 U302 ( .A1(n1132), .A2(n1212), .ZN(n1211) );
  NAND2_X2 U303 ( .A1(n1132), .A2(n1213), .ZN(n1210) );
  MUX2_X1 U304 ( .A(n1214), .B(n1215), .S(n1105), .Z(n1208) );
  NAND2_X2 U305 ( .A1(n1216), .A2(n1119), .ZN(n1215) );
  NAND2_X2 U306 ( .A1(n1217), .A2(n1119), .ZN(n1214) );
  NAND2_X2 U307 ( .A1(n1218), .A2(n1219), .ZN(B[4]) );
  MUX2_X1 U308 ( .A(n1220), .B(n1221), .S(n1154), .Z(n1219) );
  NAND2_X2 U309 ( .A1(n1150), .A2(n1222), .ZN(n1221) );
  NAND2_X2 U310 ( .A1(n1150), .A2(n1205), .ZN(n1220) );
  MUX2_X1 U311 ( .A(n1223), .B(n1224), .S(n1154), .Z(n1218) );
  NAND2_X2 U312 ( .A1(n1188), .A2(n1138), .ZN(n1224) );
  NAND2_X2 U313 ( .A1(n1181), .A2(n1138), .ZN(n1223) );
  NAND2_X2 U314 ( .A1(n1225), .A2(n1226), .ZN(n1181) );
  MUX2_X1 U315 ( .A(n1227), .B(n1228), .S(n1105), .Z(n1226) );
  NAND2_X2 U316 ( .A1(n1131), .A2(n1229), .ZN(n1228) );
  NAND2_X2 U317 ( .A1(n1131), .A2(n1230), .ZN(n1227) );
  MUX2_X1 U318 ( .A(n1231), .B(n1232), .S(n1105), .Z(n1225) );
  NAND2_X2 U319 ( .A1(n1233), .A2(n1118), .ZN(n1232) );
  NAND2_X2 U320 ( .A1(n1234), .A2(n1118), .ZN(n1231) );
  NAND2_X2 U321 ( .A1(n1235), .A2(n1236), .ZN(B[3]) );
  MUX2_X1 U322 ( .A(n1237), .B(n1238), .S(n1155), .Z(n1236) );
  NAND2_X2 U323 ( .A1(n1150), .A2(n1239), .ZN(n1238) );
  NAND2_X2 U324 ( .A1(n1150), .A2(n1222), .ZN(n1237) );
  MUX2_X1 U325 ( .A(n1240), .B(n1241), .S(n1155), .Z(n1235) );
  NAND2_X2 U326 ( .A1(n1205), .A2(n1138), .ZN(n1241) );
  NAND2_X2 U327 ( .A1(n1188), .A2(n1138), .ZN(n1240) );
  NAND2_X2 U328 ( .A1(n1242), .A2(n1243), .ZN(n1188) );
  MUX2_X1 U329 ( .A(n1244), .B(n1245), .S(n1105), .Z(n1243) );
  NAND2_X2 U330 ( .A1(n1131), .A2(n1246), .ZN(n1245) );
  NAND2_X2 U331 ( .A1(n1131), .A2(n1247), .ZN(n1244) );
  MUX2_X1 U332 ( .A(n1248), .B(n1249), .S(n1105), .Z(n1242) );
  NAND2_X2 U333 ( .A1(n1250), .A2(n1118), .ZN(n1249) );
  NAND2_X2 U334 ( .A1(n1251), .A2(n1118), .ZN(n1248) );
  NAND2_X2 U335 ( .A1(n1252), .A2(n1253), .ZN(B[31]) );
  MUX2_X1 U336 ( .A(n1254), .B(n1255), .S(n1155), .Z(n1253) );
  NAND2_X2 U337 ( .A1(n1149), .A2(n1256), .ZN(n1255) );
  NAND2_X2 U338 ( .A1(n1149), .A2(n1257), .ZN(n1254) );
  MUX2_X1 U339 ( .A(n1258), .B(n1259), .S(n1155), .Z(n1252) );
  NAND2_X2 U340 ( .A1(n1260), .A2(n1138), .ZN(n1259) );
  NAND2_X2 U341 ( .A1(n1261), .A2(n1138), .ZN(n1258) );
  NAND2_X2 U342 ( .A1(n1262), .A2(n1263), .ZN(B[30]) );
  MUX2_X1 U343 ( .A(n1264), .B(n1265), .S(n1155), .Z(n1263) );
  NAND2_X2 U344 ( .A1(n1149), .A2(n1266), .ZN(n1265) );
  NAND2_X2 U345 ( .A1(n1149), .A2(n1256), .ZN(n1264) );
  MUX2_X1 U346 ( .A(n1267), .B(n1268), .S(n1155), .Z(n1262) );
  NAND2_X2 U347 ( .A1(n1257), .A2(n1137), .ZN(n1268) );
  NAND2_X2 U348 ( .A1(n1260), .A2(n1137), .ZN(n1267) );
  NAND2_X2 U349 ( .A1(n1269), .A2(n1270), .ZN(B[2]) );
  MUX2_X1 U350 ( .A(n1271), .B(n1272), .S(n1155), .Z(n1270) );
  NAND2_X2 U351 ( .A1(n1149), .A2(n1261), .ZN(n1272) );
  NAND2_X2 U352 ( .A1(n1148), .A2(n1239), .ZN(n1271) );
  MUX2_X1 U353 ( .A(n1273), .B(n1274), .S(n1155), .Z(n1269) );
  NAND2_X2 U354 ( .A1(n1222), .A2(n1137), .ZN(n1274) );
  NAND2_X2 U355 ( .A1(n1205), .A2(n1137), .ZN(n1273) );
  NAND2_X2 U356 ( .A1(n1275), .A2(n1276), .ZN(n1205) );
  MUX2_X1 U357 ( .A(n1277), .B(n1278), .S(n1105), .Z(n1276) );
  NAND2_X2 U358 ( .A1(n1131), .A2(n1279), .ZN(n1278) );
  NAND2_X2 U359 ( .A1(n1130), .A2(n1280), .ZN(n1277) );
  MUX2_X1 U360 ( .A(n1281), .B(n1282), .S(n1105), .Z(n1275) );
  NAND2_X2 U361 ( .A1(n1195), .A2(n1118), .ZN(n1282) );
  NAND2_X2 U362 ( .A1(n1196), .A2(n1118), .ZN(n1281) );
  NAND2_X2 U363 ( .A1(n1283), .A2(n1284), .ZN(B[29]) );
  MUX2_X1 U364 ( .A(n1285), .B(n1286), .S(n1155), .Z(n1284) );
  NAND2_X2 U365 ( .A1(n1148), .A2(n1287), .ZN(n1286) );
  NAND2_X2 U366 ( .A1(n1148), .A2(n1266), .ZN(n1285) );
  MUX2_X1 U367 ( .A(n1288), .B(n1289), .S(n1155), .Z(n1283) );
  NAND2_X2 U368 ( .A1(n1256), .A2(n1137), .ZN(n1289) );
  NAND2_X2 U369 ( .A1(n1257), .A2(n1137), .ZN(n1288) );
  NAND2_X2 U370 ( .A1(n1290), .A2(n1291), .ZN(B[28]) );
  MUX2_X1 U371 ( .A(n1292), .B(n1293), .S(n1155), .Z(n1291) );
  NAND2_X2 U372 ( .A1(n1148), .A2(n1294), .ZN(n1293) );
  NAND2_X2 U373 ( .A1(n1148), .A2(n1287), .ZN(n1292) );
  MUX2_X1 U374 ( .A(n1295), .B(n1296), .S(n1155), .Z(n1290) );
  NAND2_X2 U375 ( .A1(n1266), .A2(n1137), .ZN(n1296) );
  NAND2_X2 U376 ( .A1(n1256), .A2(n1137), .ZN(n1295) );
  NAND2_X2 U377 ( .A1(n1297), .A2(n1298), .ZN(n1256) );
  MUX2_X1 U378 ( .A(n1299), .B(n1300), .S(n1105), .Z(n1298) );
  NAND2_X2 U379 ( .A1(n1130), .A2(n1301), .ZN(n1300) );
  NAND2_X2 U380 ( .A1(n1130), .A2(n1302), .ZN(n1299) );
  MUX2_X1 U381 ( .A(n1303), .B(n1304), .S(n1105), .Z(n1297) );
  NAND2_X2 U382 ( .A1(n1305), .A2(n1118), .ZN(n1304) );
  NAND2_X2 U383 ( .A1(n1306), .A2(n1118), .ZN(n1303) );
  NAND2_X2 U384 ( .A1(n1307), .A2(n1308), .ZN(B[27]) );
  MUX2_X1 U385 ( .A(n1309), .B(n1310), .S(n1156), .Z(n1308) );
  NAND2_X2 U386 ( .A1(n1147), .A2(n1311), .ZN(n1310) );
  NAND2_X2 U387 ( .A1(n1147), .A2(n1294), .ZN(n1309) );
  MUX2_X1 U388 ( .A(n1312), .B(n1313), .S(n1156), .Z(n1307) );
  NAND2_X2 U389 ( .A1(n1287), .A2(n1137), .ZN(n1313) );
  NAND2_X2 U390 ( .A1(n1266), .A2(n1137), .ZN(n1312) );
  NAND2_X2 U391 ( .A1(n1314), .A2(n1315), .ZN(n1266) );
  MUX2_X1 U392 ( .A(n1316), .B(n1317), .S(n1106), .Z(n1315) );
  NAND2_X2 U393 ( .A1(n1130), .A2(n1318), .ZN(n1317) );
  NAND2_X2 U394 ( .A1(n1130), .A2(n1319), .ZN(n1316) );
  MUX2_X1 U395 ( .A(n1320), .B(n1321), .S(n1106), .Z(n1314) );
  NAND2_X2 U396 ( .A1(n1322), .A2(n1118), .ZN(n1321) );
  NAND2_X2 U397 ( .A1(n1323), .A2(n1118), .ZN(n1320) );
  NAND2_X2 U398 ( .A1(n1324), .A2(n1325), .ZN(B[26]) );
  MUX2_X1 U399 ( .A(n1326), .B(n1327), .S(n1156), .Z(n1325) );
  NAND2_X2 U400 ( .A1(n1147), .A2(n1328), .ZN(n1327) );
  NAND2_X2 U401 ( .A1(n1147), .A2(n1311), .ZN(n1326) );
  MUX2_X1 U402 ( .A(n1329), .B(n1330), .S(n1156), .Z(n1324) );
  NAND2_X2 U403 ( .A1(n1294), .A2(n1137), .ZN(n1330) );
  NAND2_X2 U404 ( .A1(n1287), .A2(n1137), .ZN(n1329) );
  NAND2_X2 U405 ( .A1(n1331), .A2(n1332), .ZN(n1287) );
  MUX2_X1 U406 ( .A(n1333), .B(n1334), .S(n1106), .Z(n1332) );
  NAND2_X2 U407 ( .A1(n1129), .A2(n1200), .ZN(n1334) );
  NAND2_X2 U408 ( .A1(n1129), .A2(n1199), .ZN(n1333) );
  MUX2_X1 U409 ( .A(n1335), .B(n1336), .S(n1106), .Z(n1331) );
  NAND2_X2 U410 ( .A1(n1337), .A2(n1118), .ZN(n1336) );
  NAND2_X2 U411 ( .A1(n1338), .A2(n1118), .ZN(n1335) );
  NAND2_X2 U412 ( .A1(n1339), .A2(n1340), .ZN(B[25]) );
  MUX2_X1 U413 ( .A(n1341), .B(n1342), .S(n1156), .Z(n1340) );
  NAND2_X2 U414 ( .A1(n1147), .A2(n1343), .ZN(n1342) );
  NAND2_X2 U415 ( .A1(n1146), .A2(n1328), .ZN(n1341) );
  MUX2_X1 U416 ( .A(n1344), .B(n1345), .S(n1156), .Z(n1339) );
  NAND2_X2 U417 ( .A1(n1311), .A2(n1136), .ZN(n1345) );
  NAND2_X2 U418 ( .A1(n1294), .A2(n1136), .ZN(n1344) );
  NAND2_X2 U419 ( .A1(n1346), .A2(n1347), .ZN(n1294) );
  MUX2_X1 U420 ( .A(n1348), .B(n1349), .S(n1106), .Z(n1347) );
  NAND2_X2 U421 ( .A1(n1129), .A2(n1217), .ZN(n1349) );
  NAND2_X2 U422 ( .A1(n1129), .A2(n1216), .ZN(n1348) );
  MUX2_X1 U423 ( .A(n1350), .B(n1351), .S(n1106), .Z(n1346) );
  NAND2_X2 U424 ( .A1(n1352), .A2(n1117), .ZN(n1351) );
  NAND2_X2 U425 ( .A1(n1353), .A2(n1117), .ZN(n1350) );
  NAND2_X2 U426 ( .A1(n1354), .A2(n1355), .ZN(B[24]) );
  MUX2_X1 U427 ( .A(n1356), .B(n1357), .S(n1156), .Z(n1355) );
  NAND2_X2 U428 ( .A1(n1146), .A2(n1358), .ZN(n1357) );
  NAND2_X2 U429 ( .A1(n1146), .A2(n1343), .ZN(n1356) );
  MUX2_X1 U430 ( .A(n1359), .B(n1360), .S(n1156), .Z(n1354) );
  NAND2_X2 U431 ( .A1(n1328), .A2(n1136), .ZN(n1360) );
  NAND2_X2 U432 ( .A1(n1311), .A2(n1136), .ZN(n1359) );
  NAND2_X2 U433 ( .A1(n1361), .A2(n1362), .ZN(n1311) );
  MUX2_X1 U434 ( .A(n1363), .B(n1364), .S(n1106), .Z(n1362) );
  NAND2_X2 U435 ( .A1(n1129), .A2(n1234), .ZN(n1364) );
  NAND2_X2 U436 ( .A1(n1128), .A2(n1233), .ZN(n1363) );
  MUX2_X1 U437 ( .A(n1365), .B(n1366), .S(n1106), .Z(n1361) );
  NAND2_X2 U438 ( .A1(n1301), .A2(n1117), .ZN(n1366) );
  NAND2_X2 U439 ( .A1(n1302), .A2(n1117), .ZN(n1365) );
  MUX2_X1 U440 ( .A(n1369), .B(n1370), .S(n1156), .Z(n1368) );
  NAND2_X2 U441 ( .A1(n1146), .A2(n1371), .ZN(n1370) );
  NAND2_X2 U442 ( .A1(n1146), .A2(n1358), .ZN(n1369) );
  MUX2_X1 U443 ( .A(n1372), .B(n1373), .S(n1156), .Z(n1367) );
  NAND2_X2 U444 ( .A1(n1343), .A2(n1136), .ZN(n1373) );
  NAND2_X2 U445 ( .A1(n1328), .A2(n1136), .ZN(n1372) );
  NAND2_X2 U446 ( .A1(n1374), .A2(n1375), .ZN(n1328) );
  MUX2_X1 U447 ( .A(n1376), .B(n1377), .S(n1106), .Z(n1375) );
  NAND2_X2 U448 ( .A1(n1128), .A2(n1251), .ZN(n1377) );
  NAND2_X2 U449 ( .A1(n1128), .A2(n1250), .ZN(n1376) );
  MUX2_X1 U450 ( .A(n1378), .B(n1379), .S(n1106), .Z(n1374) );
  NAND2_X2 U451 ( .A1(n1318), .A2(n1117), .ZN(n1379) );
  NAND2_X2 U452 ( .A1(n1319), .A2(n1117), .ZN(n1378) );
  NAND2_X2 U453 ( .A1(n1380), .A2(n1381), .ZN(B[22]) );
  MUX2_X1 U454 ( .A(n1382), .B(n1383), .S(n1156), .Z(n1381) );
  NAND2_X2 U455 ( .A1(n1145), .A2(n1384), .ZN(n1383) );
  NAND2_X2 U456 ( .A1(n1145), .A2(n1371), .ZN(n1382) );
  MUX2_X1 U457 ( .A(n1385), .B(n1386), .S(n1156), .Z(n1380) );
  NAND2_X2 U458 ( .A1(n1358), .A2(n1136), .ZN(n1386) );
  NAND2_X2 U459 ( .A1(n1343), .A2(n1136), .ZN(n1385) );
  NAND2_X2 U460 ( .A1(n1387), .A2(n1388), .ZN(n1343) );
  MUX2_X1 U461 ( .A(n1389), .B(n1390), .S(n1106), .Z(n1388) );
  NAND2_X2 U462 ( .A1(n1128), .A2(n1196), .ZN(n1390) );
  NAND2_X2 U463 ( .A1(n1128), .A2(n1195), .ZN(n1389) );
  MUX2_X1 U464 ( .A(n1391), .B(n1392), .S(n1106), .Z(n1387) );
  NAND2_X2 U465 ( .A1(n1200), .A2(n1117), .ZN(n1392) );
  NAND2_X2 U466 ( .A1(n1199), .A2(n1117), .ZN(n1391) );
  MUX2_X1 U467 ( .A(n1395), .B(n1396), .S(n1157), .Z(n1394) );
  NAND2_X2 U468 ( .A1(n1145), .A2(n1397), .ZN(n1396) );
  NAND2_X2 U469 ( .A1(n1145), .A2(n1384), .ZN(n1395) );
  MUX2_X1 U470 ( .A(n1398), .B(n1399), .S(n1157), .Z(n1393) );
  NAND2_X2 U471 ( .A1(n1371), .A2(n1136), .ZN(n1399) );
  NAND2_X2 U472 ( .A1(n1358), .A2(n1136), .ZN(n1398) );
  NAND2_X2 U473 ( .A1(n1400), .A2(n1401), .ZN(n1358) );
  MUX2_X1 U474 ( .A(n1402), .B(n1403), .S(n1107), .Z(n1401) );
  NAND2_X2 U475 ( .A1(n1127), .A2(n1213), .ZN(n1403) );
  NAND2_X2 U476 ( .A1(n1127), .A2(n1212), .ZN(n1402) );
  MUX2_X1 U477 ( .A(n1404), .B(n1405), .S(n1107), .Z(n1400) );
  NAND2_X2 U478 ( .A1(n1217), .A2(n1117), .ZN(n1405) );
  NAND2_X2 U479 ( .A1(n1216), .A2(n1117), .ZN(n1404) );
  NAND2_X2 U480 ( .A1(n1406), .A2(n1407), .ZN(B[20]) );
  MUX2_X1 U481 ( .A(n1408), .B(n1409), .S(n1157), .Z(n1407) );
  NAND2_X2 U482 ( .A1(n1145), .A2(n1410), .ZN(n1409) );
  NAND2_X2 U483 ( .A1(n1144), .A2(n1397), .ZN(n1408) );
  MUX2_X1 U484 ( .A(n1411), .B(n1412), .S(n1157), .Z(n1406) );
  NAND2_X2 U485 ( .A1(n1384), .A2(n1136), .ZN(n1412) );
  NAND2_X2 U486 ( .A1(n1371), .A2(n1136), .ZN(n1411) );
  NAND2_X2 U487 ( .A1(n1413), .A2(n1414), .ZN(n1371) );
  MUX2_X1 U488 ( .A(n1415), .B(n1416), .S(n1107), .Z(n1414) );
  NAND2_X2 U489 ( .A1(n1127), .A2(n1230), .ZN(n1416) );
  NAND2_X2 U490 ( .A1(n1127), .A2(n1229), .ZN(n1415) );
  MUX2_X1 U491 ( .A(n1417), .B(n1418), .S(n1107), .Z(n1413) );
  NAND2_X2 U492 ( .A1(n1234), .A2(n1117), .ZN(n1418) );
  NAND2_X2 U493 ( .A1(n1233), .A2(n1117), .ZN(n1417) );
  NAND2_X2 U494 ( .A1(n1419), .A2(n1420), .ZN(B[1]) );
  MUX2_X1 U495 ( .A(n1421), .B(n1422), .S(n1157), .Z(n1420) );
  NAND2_X2 U496 ( .A1(n1144), .A2(n1260), .ZN(n1422) );
  NAND2_X2 U497 ( .A1(n1144), .A2(n1261), .ZN(n1421) );
  MUX2_X1 U498 ( .A(n1423), .B(n1424), .S(n1157), .Z(n1419) );
  NAND2_X2 U499 ( .A1(n1239), .A2(n1135), .ZN(n1424) );
  NAND2_X2 U500 ( .A1(n1222), .A2(n1135), .ZN(n1423) );
  NAND2_X2 U501 ( .A1(n1425), .A2(n1426), .ZN(n1222) );
  MUX2_X1 U502 ( .A(n1427), .B(n1428), .S(n1107), .Z(n1426) );
  NAND2_X2 U503 ( .A1(n1127), .A2(n1429), .ZN(n1428) );
  NAND2_X2 U504 ( .A1(n1126), .A2(n1430), .ZN(n1427) );
  MUX2_X1 U505 ( .A(n1431), .B(n1432), .S(n1107), .Z(n1425) );
  NAND2_X2 U506 ( .A1(n1212), .A2(n1116), .ZN(n1432) );
  NAND2_X2 U507 ( .A1(n1213), .A2(n1116), .ZN(n1431) );
  NAND2_X2 U508 ( .A1(n1433), .A2(n1434), .ZN(B[19]) );
  MUX2_X1 U509 ( .A(n1435), .B(n1436), .S(n1157), .Z(n1434) );
  NAND2_X2 U510 ( .A1(n1144), .A2(n1437), .ZN(n1436) );
  NAND2_X2 U511 ( .A1(n1144), .A2(n1410), .ZN(n1435) );
  MUX2_X1 U512 ( .A(n1438), .B(n1439), .S(n1157), .Z(n1433) );
  NAND2_X2 U513 ( .A1(n1397), .A2(n1135), .ZN(n1439) );
  NAND2_X2 U514 ( .A1(n1384), .A2(n1135), .ZN(n1438) );
  NAND2_X2 U515 ( .A1(n1440), .A2(n1441), .ZN(n1384) );
  MUX2_X1 U516 ( .A(n1442), .B(n1443), .S(n1107), .Z(n1441) );
  NAND2_X2 U517 ( .A1(n1126), .A2(n1247), .ZN(n1443) );
  NAND2_X2 U518 ( .A1(n1126), .A2(n1246), .ZN(n1442) );
  MUX2_X1 U519 ( .A(n1444), .B(n1445), .S(n1107), .Z(n1440) );
  NAND2_X2 U520 ( .A1(n1251), .A2(n1116), .ZN(n1445) );
  NAND2_X2 U521 ( .A1(n1250), .A2(n1116), .ZN(n1444) );
  NAND2_X2 U522 ( .A1(n1446), .A2(n1447), .ZN(B[18]) );
  MUX2_X1 U523 ( .A(n1448), .B(n1449), .S(n1157), .Z(n1447) );
  NAND2_X2 U524 ( .A1(n1143), .A2(n1450), .ZN(n1449) );
  NAND2_X2 U525 ( .A1(n1143), .A2(n1437), .ZN(n1448) );
  MUX2_X1 U526 ( .A(n1451), .B(n1452), .S(n1157), .Z(n1446) );
  NAND2_X2 U527 ( .A1(n1410), .A2(n1135), .ZN(n1452) );
  NAND2_X2 U528 ( .A1(n1397), .A2(n1135), .ZN(n1451) );
  NAND2_X2 U529 ( .A1(n1453), .A2(n1454), .ZN(n1397) );
  MUX2_X1 U530 ( .A(n1455), .B(n1456), .S(n1107), .Z(n1454) );
  NAND2_X2 U531 ( .A1(n1126), .A2(n1280), .ZN(n1456) );
  NAND2_X2 U532 ( .A1(n1126), .A2(n1279), .ZN(n1455) );
  MUX2_X1 U533 ( .A(n1457), .B(n1458), .S(n1107), .Z(n1453) );
  NAND2_X2 U534 ( .A1(n1196), .A2(n1116), .ZN(n1458) );
  INV_X2 U535 ( .A(n1459), .ZN(n1196) );
  MUX2_X1 U536 ( .A(n1460), .B(n1461), .S(n1111), .Z(n1459) );
  NAND2_X2 U537 ( .A1(n1195), .A2(n1116), .ZN(n1457) );
  INV_X2 U538 ( .A(n1462), .ZN(n1195) );
  MUX2_X1 U539 ( .A(n1463), .B(n1464), .S(n1111), .Z(n1462) );
  NAND2_X2 U540 ( .A1(n1465), .A2(n1466), .ZN(B[17]) );
  MUX2_X1 U541 ( .A(n1467), .B(n1468), .S(n1157), .Z(n1466) );
  NAND2_X2 U542 ( .A1(n1143), .A2(n1469), .ZN(n1468) );
  NAND2_X2 U543 ( .A1(n1143), .A2(n1450), .ZN(n1467) );
  MUX2_X1 U544 ( .A(n1470), .B(n1471), .S(n1157), .Z(n1465) );
  NAND2_X2 U545 ( .A1(n1437), .A2(n1135), .ZN(n1471) );
  NAND2_X2 U546 ( .A1(n1410), .A2(n1135), .ZN(n1470) );
  NAND2_X2 U547 ( .A1(n1472), .A2(n1473), .ZN(n1410) );
  MUX2_X1 U548 ( .A(n1474), .B(n1475), .S(n1107), .Z(n1473) );
  NAND2_X2 U549 ( .A1(n1125), .A2(n1430), .ZN(n1475) );
  NAND2_X2 U550 ( .A1(n1125), .A2(n1429), .ZN(n1474) );
  MUX2_X1 U551 ( .A(n1476), .B(n1477), .S(n1107), .Z(n1472) );
  NAND2_X2 U552 ( .A1(n1213), .A2(n1116), .ZN(n1477) );
  INV_X2 U553 ( .A(n1478), .ZN(n1213) );
  MUX2_X1 U554 ( .A(n1479), .B(n1480), .S(n1111), .Z(n1478) );
  NAND2_X2 U555 ( .A1(n1212), .A2(n1116), .ZN(n1476) );
  INV_X2 U556 ( .A(n1481), .ZN(n1212) );
  MUX2_X1 U557 ( .A(n1482), .B(n1483), .S(n1111), .Z(n1481) );
  NAND2_X2 U558 ( .A1(n1484), .A2(n1485), .ZN(B[16]) );
  MUX2_X1 U559 ( .A(n1486), .B(n1487), .S(n1158), .Z(n1485) );
  NAND2_X2 U560 ( .A1(n1143), .A2(n1488), .ZN(n1487) );
  NAND2_X2 U561 ( .A1(n1142), .A2(n1469), .ZN(n1486) );
  MUX2_X1 U562 ( .A(n1489), .B(n1490), .S(n1158), .Z(n1484) );
  NAND2_X2 U563 ( .A1(n1450), .A2(n1135), .ZN(n1490) );
  NAND2_X2 U564 ( .A1(n1437), .A2(n1135), .ZN(n1489) );
  NAND2_X2 U565 ( .A1(n1491), .A2(n1492), .ZN(n1437) );
  MUX2_X1 U566 ( .A(n1493), .B(n1494), .S(n1108), .Z(n1492) );
  NAND2_X2 U567 ( .A1(n1125), .A2(n1306), .ZN(n1494) );
  NAND2_X2 U568 ( .A1(n1125), .A2(n1305), .ZN(n1493) );
  MUX2_X1 U569 ( .A(n1495), .B(n1496), .S(n1108), .Z(n1491) );
  NAND2_X2 U570 ( .A1(n1230), .A2(n1116), .ZN(n1496) );
  NAND2_X2 U571 ( .A1(n1229), .A2(n1116), .ZN(n1495) );
  NAND2_X2 U572 ( .A1(n1497), .A2(n1498), .ZN(B[15]) );
  MUX2_X1 U573 ( .A(n1499), .B(n1500), .S(n1158), .Z(n1498) );
  NAND2_X2 U574 ( .A1(n1142), .A2(n1501), .ZN(n1500) );
  NAND2_X2 U575 ( .A1(n1142), .A2(n1488), .ZN(n1499) );
  MUX2_X1 U576 ( .A(n1502), .B(n1503), .S(n1158), .Z(n1497) );
  NAND2_X2 U577 ( .A1(n1469), .A2(n1135), .ZN(n1503) );
  NAND2_X2 U578 ( .A1(n1450), .A2(n1135), .ZN(n1502) );
  NAND2_X2 U579 ( .A1(n1504), .A2(n1505), .ZN(n1450) );
  MUX2_X1 U580 ( .A(n1506), .B(n1507), .S(n1108), .Z(n1505) );
  NAND2_X2 U581 ( .A1(n1125), .A2(n1323), .ZN(n1507) );
  NAND2_X2 U582 ( .A1(n1124), .A2(n1322), .ZN(n1506) );
  MUX2_X1 U583 ( .A(n1508), .B(n1509), .S(n1108), .Z(n1504) );
  NAND2_X2 U584 ( .A1(n1247), .A2(n1116), .ZN(n1509) );
  NAND2_X2 U585 ( .A1(n1246), .A2(n1116), .ZN(n1508) );
  NAND2_X2 U586 ( .A1(n1510), .A2(n1511), .ZN(B[14]) );
  MUX2_X1 U587 ( .A(n1512), .B(n1513), .S(n1158), .Z(n1511) );
  NAND2_X2 U588 ( .A1(n1142), .A2(n1514), .ZN(n1513) );
  NAND2_X2 U589 ( .A1(n1142), .A2(n1501), .ZN(n1512) );
  MUX2_X1 U590 ( .A(n1515), .B(n1516), .S(n1158), .Z(n1510) );
  NAND2_X2 U591 ( .A1(n1488), .A2(n1134), .ZN(n1516) );
  NAND2_X2 U592 ( .A1(n1469), .A2(n1134), .ZN(n1515) );
  NAND2_X2 U593 ( .A1(n1517), .A2(n1518), .ZN(n1469) );
  MUX2_X1 U594 ( .A(n1519), .B(n1520), .S(n1108), .Z(n1518) );
  NAND2_X2 U595 ( .A1(n1124), .A2(n1338), .ZN(n1520) );
  NAND2_X2 U596 ( .A1(n1124), .A2(n1337), .ZN(n1519) );
  MUX2_X1 U597 ( .A(n1521), .B(n1522), .S(n1108), .Z(n1517) );
  NAND2_X2 U598 ( .A1(n1280), .A2(n1115), .ZN(n1522) );
  NAND2_X2 U599 ( .A1(n1279), .A2(n1115), .ZN(n1521) );
  NAND2_X2 U600 ( .A1(n1523), .A2(n1524), .ZN(B[13]) );
  MUX2_X1 U601 ( .A(n1525), .B(n1526), .S(n1158), .Z(n1524) );
  NAND2_X2 U602 ( .A1(n1141), .A2(n1527), .ZN(n1526) );
  NAND2_X2 U603 ( .A1(n1141), .A2(n1514), .ZN(n1525) );
  MUX2_X1 U604 ( .A(n1528), .B(n1529), .S(n1158), .Z(n1523) );
  NAND2_X2 U605 ( .A1(n1501), .A2(n1134), .ZN(n1529) );
  NAND2_X2 U606 ( .A1(n1488), .A2(n1134), .ZN(n1528) );
  NAND2_X2 U607 ( .A1(n1530), .A2(n1531), .ZN(n1488) );
  MUX2_X1 U608 ( .A(n1532), .B(n1533), .S(n1108), .Z(n1531) );
  NAND2_X2 U609 ( .A1(n1124), .A2(n1353), .ZN(n1533) );
  NAND2_X2 U610 ( .A1(n1124), .A2(n1352), .ZN(n1532) );
  MUX2_X1 U611 ( .A(n1534), .B(n1535), .S(n1108), .Z(n1530) );
  NAND2_X2 U612 ( .A1(n1430), .A2(n1115), .ZN(n1535) );
  NAND2_X2 U613 ( .A1(n1429), .A2(n1115), .ZN(n1534) );
  NAND2_X2 U614 ( .A1(n1536), .A2(n1537), .ZN(B[12]) );
  MUX2_X1 U615 ( .A(n1538), .B(n1539), .S(n1158), .Z(n1537) );
  NAND2_X2 U616 ( .A1(n1141), .A2(n1169), .ZN(n1539) );
  NAND2_X2 U617 ( .A1(n1141), .A2(n1527), .ZN(n1538) );
  MUX2_X1 U618 ( .A(n1540), .B(n1541), .S(n1158), .Z(n1536) );
  NAND2_X2 U619 ( .A1(n1514), .A2(n1134), .ZN(n1541) );
  NAND2_X2 U620 ( .A1(n1501), .A2(n1134), .ZN(n1540) );
  NAND2_X2 U621 ( .A1(n1542), .A2(n1543), .ZN(n1501) );
  MUX2_X1 U622 ( .A(n1544), .B(n1545), .S(n1108), .Z(n1543) );
  NAND2_X2 U623 ( .A1(n1123), .A2(n1302), .ZN(n1545) );
  NAND2_X2 U624 ( .A1(n1123), .A2(n1301), .ZN(n1544) );
  MUX2_X1 U625 ( .A(n1546), .B(n1547), .S(n1108), .Z(n1542) );
  NAND2_X2 U626 ( .A1(n1306), .A2(n1115), .ZN(n1547) );
  NAND2_X2 U627 ( .A1(n1305), .A2(n1115), .ZN(n1546) );
  NAND2_X2 U628 ( .A1(n1548), .A2(n1549), .ZN(B[11]) );
  MUX2_X1 U629 ( .A(n1550), .B(n1551), .S(n1158), .Z(n1549) );
  NAND2_X2 U630 ( .A1(n1141), .A2(n1168), .ZN(n1551) );
  NAND2_X2 U631 ( .A1(n1140), .A2(n1169), .ZN(n1550) );
  MUX2_X1 U632 ( .A(n1552), .B(n1553), .S(n1158), .Z(n1548) );
  NAND2_X2 U633 ( .A1(n1527), .A2(n1134), .ZN(n1553) );
  NAND2_X2 U634 ( .A1(n1514), .A2(n1134), .ZN(n1552) );
  NAND2_X2 U635 ( .A1(n1554), .A2(n1555), .ZN(n1514) );
  MUX2_X1 U636 ( .A(n1556), .B(n1557), .S(n1108), .Z(n1555) );
  NAND2_X2 U637 ( .A1(n1123), .A2(n1319), .ZN(n1557) );
  NAND2_X2 U638 ( .A1(n1123), .A2(n1318), .ZN(n1556) );
  MUX2_X1 U639 ( .A(n1558), .B(n1559), .S(n1108), .Z(n1554) );
  NAND2_X2 U640 ( .A1(n1323), .A2(n1115), .ZN(n1559) );
  NAND2_X2 U641 ( .A1(n1322), .A2(n1115), .ZN(n1558) );
  NAND2_X2 U642 ( .A1(n1560), .A2(n1561), .ZN(B[10]) );
  MUX2_X1 U643 ( .A(n1562), .B(n1563), .S(n1159), .Z(n1561) );
  NAND2_X2 U644 ( .A1(n1140), .A2(n1165), .ZN(n1563) );
  NAND2_X2 U645 ( .A1(n1564), .A2(n1565), .ZN(n1165) );
  MUX2_X1 U646 ( .A(n1566), .B(n1567), .S(n1109), .Z(n1565) );
  NAND2_X2 U647 ( .A1(n1123), .A2(n1250), .ZN(n1567) );
  INV_X2 U648 ( .A(n1568), .ZN(n1250) );
  MUX2_X1 U649 ( .A(n1569), .B(n1570), .S(n1111), .Z(n1568) );
  NAND2_X2 U650 ( .A1(n1122), .A2(n1251), .ZN(n1566) );
  INV_X2 U651 ( .A(n1571), .ZN(n1251) );
  MUX2_X1 U652 ( .A(n1572), .B(n1573), .S(n1111), .Z(n1571) );
  MUX2_X1 U653 ( .A(n1574), .B(n1575), .S(n1109), .Z(n1564) );
  NAND2_X2 U654 ( .A1(n1319), .A2(n1115), .ZN(n1575) );
  INV_X2 U655 ( .A(n1576), .ZN(n1319) );
  MUX2_X1 U656 ( .A(n1577), .B(n1578), .S(n1111), .Z(n1576) );
  NAND2_X2 U657 ( .A1(n1318), .A2(n1115), .ZN(n1574) );
  INV_X2 U658 ( .A(n1579), .ZN(n1318) );
  MUX2_X1 U659 ( .A(n1580), .B(n1581), .S(n1111), .Z(n1579) );
  NAND2_X2 U660 ( .A1(n1140), .A2(n1168), .ZN(n1562) );
  NAND2_X2 U661 ( .A1(n1582), .A2(n1583), .ZN(n1168) );
  MUX2_X1 U662 ( .A(n1584), .B(n1585), .S(n1109), .Z(n1583) );
  NAND2_X2 U663 ( .A1(n1122), .A2(n1233), .ZN(n1585) );
  INV_X2 U664 ( .A(n1586), .ZN(n1233) );
  MUX2_X1 U665 ( .A(n1587), .B(n1588), .S(n1111), .Z(n1586) );
  NAND2_X2 U666 ( .A1(n1122), .A2(n1234), .ZN(n1584) );
  INV_X2 U667 ( .A(n1589), .ZN(n1234) );
  MUX2_X1 U668 ( .A(n1590), .B(n1591), .S(n1111), .Z(n1589) );
  MUX2_X1 U669 ( .A(n1592), .B(n1593), .S(n1109), .Z(n1582) );
  NAND2_X2 U670 ( .A1(n1302), .A2(n1115), .ZN(n1593) );
  INV_X2 U671 ( .A(n1594), .ZN(n1302) );
  MUX2_X1 U672 ( .A(n1595), .B(n1596), .S(n1111), .Z(n1594) );
  NAND2_X2 U673 ( .A1(n1301), .A2(n1115), .ZN(n1592) );
  INV_X2 U674 ( .A(n1597), .ZN(n1301) );
  MUX2_X1 U675 ( .A(n1598), .B(n1599), .S(n1111), .Z(n1597) );
  MUX2_X1 U676 ( .A(n1600), .B(n1601), .S(n1159), .Z(n1560) );
  NAND2_X2 U677 ( .A1(n1169), .A2(n1134), .ZN(n1601) );
  NAND2_X2 U678 ( .A1(n1602), .A2(n1603), .ZN(n1169) );
  MUX2_X1 U679 ( .A(n1604), .B(n1605), .S(n1109), .Z(n1603) );
  NAND2_X2 U680 ( .A1(n1122), .A2(n1216), .ZN(n1605) );
  INV_X2 U681 ( .A(n1606), .ZN(n1216) );
  MUX2_X1 U682 ( .A(n1607), .B(n1608), .S(n1112), .Z(n1606) );
  NAND2_X2 U683 ( .A1(n1122), .A2(n1217), .ZN(n1604) );
  INV_X2 U684 ( .A(n1609), .ZN(n1217) );
  MUX2_X1 U685 ( .A(n1610), .B(n1611), .S(n1112), .Z(n1609) );
  MUX2_X1 U686 ( .A(n1612), .B(n1613), .S(n1109), .Z(n1602) );
  NAND2_X2 U687 ( .A1(n1353), .A2(n1114), .ZN(n1613) );
  NAND2_X2 U688 ( .A1(n1352), .A2(n1114), .ZN(n1612) );
  NAND2_X2 U689 ( .A1(n1527), .A2(n1134), .ZN(n1600) );
  NAND2_X2 U690 ( .A1(n1614), .A2(n1615), .ZN(n1527) );
  MUX2_X1 U691 ( .A(n1616), .B(n1617), .S(n1109), .Z(n1615) );
  NAND2_X2 U692 ( .A1(n1121), .A2(n1199), .ZN(n1617) );
  INV_X2 U693 ( .A(n1618), .ZN(n1199) );
  MUX2_X1 U694 ( .A(n1619), .B(n1620), .S(n1112), .Z(n1618) );
  NAND2_X2 U695 ( .A1(n1121), .A2(n1200), .ZN(n1616) );
  INV_X2 U696 ( .A(n1621), .ZN(n1200) );
  MUX2_X1 U697 ( .A(n1622), .B(n1623), .S(n1112), .Z(n1621) );
  MUX2_X1 U698 ( .A(n1624), .B(n1625), .S(n1109), .Z(n1614) );
  NAND2_X2 U699 ( .A1(n1338), .A2(n1114), .ZN(n1625) );
  NAND2_X2 U700 ( .A1(n1337), .A2(n1114), .ZN(n1624) );
  NAND2_X2 U701 ( .A1(n1626), .A2(n1627), .ZN(B[0]) );
  MUX2_X1 U702 ( .A(n1628), .B(n1629), .S(n1159), .Z(n1627) );
  NAND2_X2 U703 ( .A1(n1140), .A2(n1257), .ZN(n1629) );
  NAND2_X2 U704 ( .A1(n1630), .A2(n1631), .ZN(n1257) );
  MUX2_X1 U705 ( .A(n1632), .B(n1633), .S(n1109), .Z(n1631) );
  NAND2_X2 U706 ( .A1(n1121), .A2(n1352), .ZN(n1633) );
  INV_X2 U707 ( .A(n1634), .ZN(n1352) );
  MUX2_X1 U708 ( .A(n1483), .B(n1479), .S(n1112), .Z(n1634) );
  NAND2_X2 U709 ( .A1(n1121), .A2(n1353), .ZN(n1632) );
  INV_X2 U710 ( .A(n1635), .ZN(n1353) );
  MUX2_X1 U711 ( .A(n1480), .B(n1482), .S(n1112), .Z(n1635) );
  MUX2_X1 U712 ( .A(n1636), .B(n1637), .S(n1109), .Z(n1630) );
  NAND2_X2 U713 ( .A1(n1429), .A2(n1114), .ZN(n1637) );
  INV_X2 U714 ( .A(n1638), .ZN(n1429) );
  MUX2_X1 U715 ( .A(n1608), .B(n1610), .S(n1112), .Z(n1638) );
  NAND2_X2 U716 ( .A1(n1430), .A2(n1114), .ZN(n1636) );
  INV_X2 U717 ( .A(n1639), .ZN(n1430) );
  MUX2_X1 U718 ( .A(n1611), .B(n1607), .S(n1112), .Z(n1639) );
  NAND2_X2 U719 ( .A1(n1140), .A2(n1260), .ZN(n1628) );
  NAND2_X2 U720 ( .A1(n1640), .A2(n1641), .ZN(n1260) );
  MUX2_X1 U721 ( .A(n1642), .B(n1643), .S(n1109), .Z(n1641) );
  NAND2_X2 U722 ( .A1(n1121), .A2(n1337), .ZN(n1643) );
  INV_X2 U723 ( .A(n1644), .ZN(n1337) );
  MUX2_X1 U724 ( .A(n1464), .B(n1460), .S(n1112), .Z(n1644) );
  NAND2_X2 U725 ( .A1(n1120), .A2(n1338), .ZN(n1642) );
  INV_X2 U726 ( .A(n1645), .ZN(n1338) );
  MUX2_X1 U727 ( .A(n1461), .B(n1463), .S(n1112), .Z(n1645) );
  MUX2_X1 U728 ( .A(n1646), .B(n1647), .S(n1109), .Z(n1640) );
  NAND2_X2 U729 ( .A1(n1279), .A2(n1114), .ZN(n1647) );
  INV_X2 U730 ( .A(n1648), .ZN(n1279) );
  MUX2_X1 U731 ( .A(n1620), .B(n1622), .S(n1112), .Z(n1648) );
  NAND2_X2 U732 ( .A1(n1280), .A2(n1114), .ZN(n1646) );
  INV_X2 U733 ( .A(n1649), .ZN(n1280) );
  MUX2_X1 U734 ( .A(n1623), .B(n1619), .S(n1112), .Z(n1649) );
  MUX2_X1 U735 ( .A(n1650), .B(n1651), .S(n1159), .Z(n1626) );
  NAND2_X2 U736 ( .A1(n1261), .A2(n1134), .ZN(n1651) );
  NAND2_X2 U737 ( .A1(n1652), .A2(n1653), .ZN(n1261) );
  MUX2_X1 U738 ( .A(n1654), .B(n1655), .S(n1110), .Z(n1653) );
  NAND2_X2 U739 ( .A1(n1120), .A2(n1322), .ZN(n1655) );
  INV_X2 U740 ( .A(n1656), .ZN(n1322) );
  MUX2_X1 U741 ( .A(n1570), .B(n1572), .S(n1113), .Z(n1656) );
  NAND2_X2 U742 ( .A1(n1120), .A2(n1323), .ZN(n1654) );
  INV_X2 U743 ( .A(n1657), .ZN(n1323) );
  MUX2_X1 U744 ( .A(n1573), .B(n1569), .S(n1113), .Z(n1657) );
  MUX2_X1 U745 ( .A(n1658), .B(n1659), .S(n1110), .Z(n1652) );
  NAND2_X2 U746 ( .A1(n1246), .A2(n1114), .ZN(n1659) );
  INV_X2 U747 ( .A(n1660), .ZN(n1246) );
  MUX2_X1 U748 ( .A(n1578), .B(n1580), .S(n1113), .Z(n1660) );
  NAND2_X2 U749 ( .A1(n1247), .A2(n1114), .ZN(n1658) );
  INV_X2 U750 ( .A(n1661), .ZN(n1247) );
  MUX2_X1 U751 ( .A(n1581), .B(n1577), .S(n1113), .Z(n1661) );
  NAND2_X2 U752 ( .A1(n1239), .A2(n1134), .ZN(n1650) );
  NAND2_X2 U753 ( .A1(n1662), .A2(n1663), .ZN(n1239) );
  MUX2_X1 U754 ( .A(n1664), .B(n1665), .S(n1110), .Z(n1663) );
  NAND2_X2 U755 ( .A1(n1120), .A2(n1305), .ZN(n1665) );
  INV_X2 U756 ( .A(n1666), .ZN(n1305) );
  MUX2_X1 U757 ( .A(n1588), .B(n1590), .S(n1113), .Z(n1666) );
  NAND2_X2 U758 ( .A1(n1120), .A2(n1306), .ZN(n1664) );
  INV_X2 U759 ( .A(n1667), .ZN(n1306) );
  MUX2_X1 U760 ( .A(n1591), .B(n1587), .S(n1113), .Z(n1667) );
  MUX2_X1 U761 ( .A(n1668), .B(n1669), .S(n1110), .Z(n1662) );
  NAND2_X2 U762 ( .A1(n1229), .A2(n1114), .ZN(n1669) );
  INV_X2 U763 ( .A(n1670), .ZN(n1229) );
  MUX2_X1 U764 ( .A(n1596), .B(n1598), .S(n1113), .Z(n1670) );
  NAND2_X2 U765 ( .A1(n1230), .A2(n1114), .ZN(n1668) );
  INV_X2 U766 ( .A(n1671), .ZN(n1230) );
  MUX2_X1 U767 ( .A(n1599), .B(n1595), .S(n1113), .Z(n1671) );
endmodule


module up_island_DW_rbsh_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672;

  NAND2_X1 U170 ( .A1(n1171), .A2(n1172), .ZN(B[8]) );
  NAND2_X1 U171 ( .A1(n1178), .A2(n1179), .ZN(B[7]) );
  NAND2_X1 U172 ( .A1(n1153), .A2(n1354), .ZN(n1357) );
  NAND2_X1 U173 ( .A1(n1354), .A2(n1143), .ZN(n1352) );
  NAND2_X1 U174 ( .A1(n1152), .A2(n1354), .ZN(n1384) );
  NAND2_X1 U175 ( .A1(n1354), .A2(n1143), .ZN(n1379) );
  MUX2_X1 U176 ( .A(n1576), .B(n1570), .S(n1127), .Z(n1645) );
  NAND2_X1 U177 ( .A1(n1381), .A2(n1382), .ZN(B[22]) );
  INV_X1 U178 ( .A(A[29]), .ZN(n1570) );
  NAND2_X1 U179 ( .A1(n1406), .A2(n1142), .ZN(n1445) );
  NAND2_X1 U180 ( .A1(n1150), .A2(n1406), .ZN(n1450) );
  NAND2_X1 U181 ( .A1(n1151), .A2(n1406), .ZN(n1409) );
  NAND2_X1 U182 ( .A1(n1406), .A2(n1143), .ZN(n1404) );
  NAND2_X1 U183 ( .A1(n1368), .A2(n1369), .ZN(B[23]) );
  INV_X1 U184 ( .A(A[30]), .ZN(n1614) );
  INV_X1 U185 ( .A(A[1]), .ZN(n1462) );
  INV_X1 U186 ( .A(A[2]), .ZN(n1618) );
  NAND2_X1 U187 ( .A1(n1253), .A2(n1254), .ZN(B[31]) );
  INV_X1 U188 ( .A(A[28]), .ZN(n1602) );
  INV_X1 U189 ( .A(A[3]), .ZN(n1586) );
  INV_X1 U190 ( .A(A[4]), .ZN(n1603) );
  INV_X1 U191 ( .A(A[26]), .ZN(n1617) );
  INV_X1 U192 ( .A(A[0]), .ZN(n1481) );
  INV_X1 U193 ( .A(A[27]), .ZN(n1585) );
  INV_X1 U194 ( .A(A[23]), .ZN(n1591) );
  INV_X1 U195 ( .A(A[22]), .ZN(n1623) );
  INV_X1 U196 ( .A(A[24]), .ZN(n1480) );
  INV_X1 U197 ( .A(A[25]), .ZN(n1461) );
  INV_X1 U198 ( .A(A[31]), .ZN(n1582) );
  INV_X1 U199 ( .A(A[19]), .ZN(n1594) );
  INV_X1 U200 ( .A(A[21]), .ZN(n1576) );
  INV_X1 U201 ( .A(A[15]), .ZN(n1590) );
  INV_X1 U202 ( .A(A[18]), .ZN(n1626) );
  INV_X1 U203 ( .A(A[17]), .ZN(n1457) );
  INV_X1 U204 ( .A(A[13]), .ZN(n1575) );
  INV_X1 U205 ( .A(A[7]), .ZN(n1583) );
  INV_X1 U206 ( .A(A[11]), .ZN(n1593) );
  INV_X1 U207 ( .A(A[20]), .ZN(n1608) );
  INV_X1 U208 ( .A(A[16]), .ZN(n1476) );
  INV_X1 U209 ( .A(A[9]), .ZN(n1456) );
  INV_X1 U210 ( .A(A[12]), .ZN(n1607) );
  INV_X1 U211 ( .A(A[6]), .ZN(n1615) );
  INV_X1 U212 ( .A(A[14]), .ZN(n1622) );
  INV_X1 U213 ( .A(A[8]), .ZN(n1475) );
  INV_X1 U214 ( .A(A[10]), .ZN(n1625) );
  INV_X1 U215 ( .A(A[5]), .ZN(n1571) );
  INV_X1 U216 ( .A(n1124), .ZN(n1106) );
  INV_X1 U217 ( .A(n1124), .ZN(n1107) );
  INV_X1 U218 ( .A(n1125), .ZN(n1108) );
  INV_X1 U219 ( .A(n1125), .ZN(n1109) );
  INV_X1 U220 ( .A(n1125), .ZN(n1110) );
  INV_X1 U221 ( .A(n1125), .ZN(n1111) );
  CLKBUF_X3 U222 ( .A(SH[4]), .Z(n1112) );
  CLKBUF_X3 U223 ( .A(SH[4]), .Z(n1113) );
  CLKBUF_X3 U224 ( .A(SH[4]), .Z(n1114) );
  CLKBUF_X3 U225 ( .A(SH[4]), .Z(n1115) );
  CLKBUF_X3 U226 ( .A(SH[4]), .Z(n1116) );
  CLKBUF_X3 U227 ( .A(SH[4]), .Z(n1117) );
  CLKBUF_X3 U228 ( .A(SH[4]), .Z(n1118) );
  CLKBUF_X3 U229 ( .A(SH[4]), .Z(n1119) );
  CLKBUF_X3 U230 ( .A(SH[4]), .Z(n1120) );
  CLKBUF_X3 U231 ( .A(SH[4]), .Z(n1121) );
  CLKBUF_X3 U232 ( .A(SH[4]), .Z(n1122) );
  CLKBUF_X3 U233 ( .A(SH[4]), .Z(n1123) );
  CLKBUF_X3 U234 ( .A(SH[4]), .Z(n1124) );
  CLKBUF_X3 U235 ( .A(SH[4]), .Z(n1125) );
  CLKBUF_X3 U236 ( .A(SH[3]), .Z(n1126) );
  CLKBUF_X3 U237 ( .A(SH[3]), .Z(n1127) );
  CLKBUF_X3 U238 ( .A(SH[3]), .Z(n1128) );
  CLKBUF_X3 U239 ( .A(SH[2]), .Z(n1129) );
  CLKBUF_X3 U240 ( .A(SH[2]), .Z(n1130) );
  CLKBUF_X3 U241 ( .A(SH[2]), .Z(n1131) );
  CLKBUF_X3 U242 ( .A(SH[2]), .Z(n1132) );
  CLKBUF_X3 U243 ( .A(SH[2]), .Z(n1133) );
  CLKBUF_X3 U244 ( .A(SH[2]), .Z(n1134) );
  CLKBUF_X3 U245 ( .A(SH[1]), .Z(n1135) );
  CLKBUF_X3 U246 ( .A(SH[1]), .Z(n1136) );
  CLKBUF_X3 U247 ( .A(SH[1]), .Z(n1137) );
  CLKBUF_X3 U248 ( .A(SH[1]), .Z(n1138) );
  CLKBUF_X3 U249 ( .A(SH[1]), .Z(n1139) );
  CLKBUF_X3 U250 ( .A(SH[1]), .Z(n1140) );
  INV_X1 U251 ( .A(n1159), .ZN(n1141) );
  INV_X1 U252 ( .A(n1159), .ZN(n1142) );
  INV_X1 U253 ( .A(n1160), .ZN(n1143) );
  INV_X1 U254 ( .A(n1160), .ZN(n1144) );
  INV_X1 U255 ( .A(n1160), .ZN(n1145) );
  INV_X1 U256 ( .A(n1160), .ZN(n1146) );
  CLKBUF_X3 U257 ( .A(SH[0]), .Z(n1147) );
  CLKBUF_X3 U258 ( .A(SH[0]), .Z(n1148) );
  CLKBUF_X3 U259 ( .A(SH[0]), .Z(n1149) );
  CLKBUF_X3 U260 ( .A(SH[0]), .Z(n1150) );
  CLKBUF_X3 U261 ( .A(SH[0]), .Z(n1151) );
  CLKBUF_X3 U262 ( .A(SH[0]), .Z(n1152) );
  CLKBUF_X3 U263 ( .A(SH[0]), .Z(n1153) );
  CLKBUF_X3 U264 ( .A(SH[0]), .Z(n1154) );
  CLKBUF_X3 U265 ( .A(SH[0]), .Z(n1155) );
  CLKBUF_X3 U266 ( .A(SH[0]), .Z(n1156) );
  CLKBUF_X3 U267 ( .A(SH[0]), .Z(n1157) );
  CLKBUF_X3 U268 ( .A(SH[0]), .Z(n1158) );
  CLKBUF_X3 U269 ( .A(SH[0]), .Z(n1159) );
  CLKBUF_X3 U270 ( .A(SH[0]), .Z(n1160) );
  NAND2_X2 U271 ( .A1(n1161), .A2(n1162), .ZN(B[9]) );
  MUX2_X1 U272 ( .A(n1163), .B(n1164), .S(n1135), .Z(n1162) );
  NAND2_X2 U273 ( .A1(n1159), .A2(n1165), .ZN(n1164) );
  NAND2_X2 U274 ( .A1(n1159), .A2(n1166), .ZN(n1163) );
  MUX2_X1 U275 ( .A(n1167), .B(n1168), .S(n1135), .Z(n1161) );
  NAND2_X2 U276 ( .A1(n1169), .A2(n1146), .ZN(n1168) );
  NAND2_X2 U277 ( .A1(n1170), .A2(n1146), .ZN(n1167) );
  MUX2_X1 U278 ( .A(n1173), .B(n1174), .S(n1135), .Z(n1172) );
  NAND2_X2 U279 ( .A1(n1159), .A2(n1169), .ZN(n1174) );
  NAND2_X2 U280 ( .A1(n1159), .A2(n1170), .ZN(n1173) );
  MUX2_X1 U281 ( .A(n1175), .B(n1176), .S(n1135), .Z(n1171) );
  NAND2_X2 U282 ( .A1(n1166), .A2(n1146), .ZN(n1176) );
  NAND2_X2 U283 ( .A1(n1177), .A2(n1146), .ZN(n1175) );
  MUX2_X1 U284 ( .A(n1180), .B(n1181), .S(n1135), .Z(n1179) );
  NAND2_X2 U285 ( .A1(n1158), .A2(n1166), .ZN(n1181) );
  NAND2_X2 U286 ( .A1(n1158), .A2(n1177), .ZN(n1180) );
  MUX2_X1 U287 ( .A(n1182), .B(n1183), .S(n1135), .Z(n1178) );
  NAND2_X2 U288 ( .A1(n1170), .A2(n1145), .ZN(n1183) );
  NAND2_X2 U289 ( .A1(n1184), .A2(n1145), .ZN(n1182) );
  NAND2_X2 U290 ( .A1(n1185), .A2(n1186), .ZN(B[6]) );
  MUX2_X1 U291 ( .A(n1187), .B(n1188), .S(n1135), .Z(n1186) );
  NAND2_X2 U292 ( .A1(n1158), .A2(n1170), .ZN(n1188) );
  NAND2_X2 U293 ( .A1(n1189), .A2(n1190), .ZN(n1170) );
  MUX2_X1 U294 ( .A(n1191), .B(n1192), .S(n1129), .Z(n1190) );
  NAND2_X2 U295 ( .A1(n1124), .A2(n1193), .ZN(n1192) );
  NAND2_X2 U296 ( .A1(n1124), .A2(n1194), .ZN(n1191) );
  MUX2_X1 U297 ( .A(n1195), .B(n1196), .S(n1129), .Z(n1189) );
  NAND2_X2 U298 ( .A1(n1197), .A2(n1111), .ZN(n1196) );
  NAND2_X2 U299 ( .A1(n1198), .A2(n1111), .ZN(n1195) );
  NAND2_X2 U300 ( .A1(n1158), .A2(n1184), .ZN(n1187) );
  MUX2_X1 U301 ( .A(n1199), .B(n1200), .S(n1135), .Z(n1185) );
  NAND2_X2 U302 ( .A1(n1177), .A2(n1145), .ZN(n1200) );
  NAND2_X2 U303 ( .A1(n1201), .A2(n1145), .ZN(n1199) );
  NAND2_X2 U304 ( .A1(n1202), .A2(n1203), .ZN(B[5]) );
  MUX2_X1 U305 ( .A(n1204), .B(n1205), .S(n1135), .Z(n1203) );
  NAND2_X2 U306 ( .A1(n1158), .A2(n1177), .ZN(n1205) );
  NAND2_X2 U307 ( .A1(n1206), .A2(n1207), .ZN(n1177) );
  MUX2_X1 U308 ( .A(n1208), .B(n1209), .S(n1129), .Z(n1207) );
  NAND2_X2 U309 ( .A1(n1124), .A2(n1210), .ZN(n1209) );
  NAND2_X2 U310 ( .A1(n1124), .A2(n1211), .ZN(n1208) );
  MUX2_X1 U311 ( .A(n1212), .B(n1213), .S(n1129), .Z(n1206) );
  NAND2_X2 U312 ( .A1(n1214), .A2(n1111), .ZN(n1213) );
  NAND2_X2 U313 ( .A1(n1215), .A2(n1111), .ZN(n1212) );
  NAND2_X2 U314 ( .A1(n1157), .A2(n1201), .ZN(n1204) );
  MUX2_X1 U315 ( .A(n1216), .B(n1217), .S(n1135), .Z(n1202) );
  NAND2_X2 U316 ( .A1(n1184), .A2(n1145), .ZN(n1217) );
  NAND2_X2 U317 ( .A1(n1218), .A2(n1145), .ZN(n1216) );
  NAND2_X2 U318 ( .A1(n1219), .A2(n1220), .ZN(B[4]) );
  MUX2_X1 U319 ( .A(n1221), .B(n1222), .S(n1135), .Z(n1220) );
  NAND2_X2 U320 ( .A1(n1157), .A2(n1184), .ZN(n1222) );
  NAND2_X2 U321 ( .A1(n1223), .A2(n1224), .ZN(n1184) );
  MUX2_X1 U322 ( .A(n1225), .B(n1226), .S(n1129), .Z(n1224) );
  NAND2_X2 U323 ( .A1(n1123), .A2(n1227), .ZN(n1226) );
  NAND2_X2 U324 ( .A1(n1123), .A2(n1228), .ZN(n1225) );
  MUX2_X1 U325 ( .A(n1229), .B(n1230), .S(n1129), .Z(n1223) );
  NAND2_X2 U326 ( .A1(n1231), .A2(n1110), .ZN(n1230) );
  NAND2_X2 U327 ( .A1(n1232), .A2(n1110), .ZN(n1229) );
  NAND2_X2 U328 ( .A1(n1157), .A2(n1218), .ZN(n1221) );
  MUX2_X1 U329 ( .A(n1233), .B(n1234), .S(n1135), .Z(n1219) );
  NAND2_X2 U330 ( .A1(n1201), .A2(n1145), .ZN(n1234) );
  NAND2_X2 U331 ( .A1(n1235), .A2(n1145), .ZN(n1233) );
  NAND2_X2 U332 ( .A1(n1236), .A2(n1237), .ZN(B[3]) );
  MUX2_X1 U333 ( .A(n1238), .B(n1239), .S(n1136), .Z(n1237) );
  NAND2_X2 U334 ( .A1(n1157), .A2(n1201), .ZN(n1239) );
  NAND2_X2 U335 ( .A1(n1240), .A2(n1241), .ZN(n1201) );
  MUX2_X1 U336 ( .A(n1242), .B(n1243), .S(n1129), .Z(n1241) );
  NAND2_X2 U337 ( .A1(n1123), .A2(n1244), .ZN(n1243) );
  NAND2_X2 U338 ( .A1(n1123), .A2(n1245), .ZN(n1242) );
  MUX2_X1 U339 ( .A(n1246), .B(n1247), .S(n1129), .Z(n1240) );
  NAND2_X2 U340 ( .A1(n1248), .A2(n1110), .ZN(n1247) );
  NAND2_X2 U341 ( .A1(n1249), .A2(n1110), .ZN(n1246) );
  NAND2_X2 U342 ( .A1(n1157), .A2(n1235), .ZN(n1238) );
  MUX2_X1 U343 ( .A(n1250), .B(n1251), .S(n1136), .Z(n1236) );
  NAND2_X2 U344 ( .A1(n1218), .A2(n1145), .ZN(n1251) );
  NAND2_X2 U345 ( .A1(n1252), .A2(n1145), .ZN(n1250) );
  MUX2_X1 U346 ( .A(n1255), .B(n1256), .S(n1136), .Z(n1254) );
  NAND2_X2 U347 ( .A1(n1156), .A2(n1257), .ZN(n1256) );
  NAND2_X2 U348 ( .A1(n1156), .A2(n1258), .ZN(n1255) );
  MUX2_X1 U349 ( .A(n1259), .B(n1260), .S(n1136), .Z(n1253) );
  NAND2_X2 U350 ( .A1(n1261), .A2(n1145), .ZN(n1260) );
  NAND2_X2 U351 ( .A1(n1262), .A2(n1145), .ZN(n1259) );
  NAND2_X2 U352 ( .A1(n1263), .A2(n1264), .ZN(B[30]) );
  MUX2_X1 U353 ( .A(n1265), .B(n1266), .S(n1136), .Z(n1264) );
  NAND2_X2 U354 ( .A1(n1156), .A2(n1261), .ZN(n1266) );
  NAND2_X2 U355 ( .A1(n1156), .A2(n1262), .ZN(n1265) );
  MUX2_X1 U356 ( .A(n1267), .B(n1268), .S(n1136), .Z(n1263) );
  NAND2_X2 U357 ( .A1(n1258), .A2(n1144), .ZN(n1268) );
  NAND2_X2 U358 ( .A1(n1269), .A2(n1144), .ZN(n1267) );
  NAND2_X2 U359 ( .A1(n1270), .A2(n1271), .ZN(B[2]) );
  MUX2_X1 U360 ( .A(n1272), .B(n1273), .S(n1136), .Z(n1271) );
  NAND2_X2 U361 ( .A1(n1156), .A2(n1218), .ZN(n1273) );
  NAND2_X2 U362 ( .A1(n1274), .A2(n1275), .ZN(n1218) );
  MUX2_X1 U363 ( .A(n1276), .B(n1277), .S(n1129), .Z(n1275) );
  NAND2_X2 U364 ( .A1(n1123), .A2(n1194), .ZN(n1277) );
  NAND2_X2 U365 ( .A1(n1122), .A2(n1278), .ZN(n1276) );
  MUX2_X1 U366 ( .A(n1279), .B(n1280), .S(n1129), .Z(n1274) );
  NAND2_X2 U367 ( .A1(n1198), .A2(n1110), .ZN(n1280) );
  NAND2_X2 U368 ( .A1(n1281), .A2(n1110), .ZN(n1279) );
  NAND2_X2 U369 ( .A1(n1155), .A2(n1252), .ZN(n1272) );
  MUX2_X1 U370 ( .A(n1282), .B(n1283), .S(n1136), .Z(n1270) );
  NAND2_X2 U371 ( .A1(n1235), .A2(n1144), .ZN(n1283) );
  NAND2_X2 U372 ( .A1(n1257), .A2(n1144), .ZN(n1282) );
  NAND2_X2 U373 ( .A1(n1284), .A2(n1285), .ZN(B[29]) );
  MUX2_X1 U374 ( .A(n1286), .B(n1287), .S(n1136), .Z(n1285) );
  NAND2_X2 U375 ( .A1(n1155), .A2(n1258), .ZN(n1287) );
  NAND2_X2 U376 ( .A1(n1155), .A2(n1269), .ZN(n1286) );
  MUX2_X1 U377 ( .A(n1288), .B(n1289), .S(n1136), .Z(n1284) );
  NAND2_X2 U378 ( .A1(n1262), .A2(n1144), .ZN(n1289) );
  NAND2_X2 U379 ( .A1(n1290), .A2(n1144), .ZN(n1288) );
  NAND2_X2 U380 ( .A1(n1291), .A2(n1292), .ZN(B[28]) );
  MUX2_X1 U381 ( .A(n1293), .B(n1294), .S(n1136), .Z(n1292) );
  NAND2_X2 U382 ( .A1(n1155), .A2(n1262), .ZN(n1294) );
  NAND2_X2 U383 ( .A1(n1295), .A2(n1296), .ZN(n1262) );
  MUX2_X1 U384 ( .A(n1297), .B(n1298), .S(n1129), .Z(n1296) );
  NAND2_X2 U385 ( .A1(n1122), .A2(n1299), .ZN(n1298) );
  NAND2_X2 U386 ( .A1(n1122), .A2(n1300), .ZN(n1297) );
  MUX2_X1 U387 ( .A(n1301), .B(n1302), .S(n1129), .Z(n1295) );
  NAND2_X2 U388 ( .A1(n1303), .A2(n1110), .ZN(n1302) );
  NAND2_X2 U389 ( .A1(n1304), .A2(n1110), .ZN(n1301) );
  NAND2_X2 U390 ( .A1(n1155), .A2(n1290), .ZN(n1293) );
  MUX2_X1 U391 ( .A(n1305), .B(n1306), .S(n1136), .Z(n1291) );
  NAND2_X2 U392 ( .A1(n1269), .A2(n1144), .ZN(n1306) );
  NAND2_X2 U393 ( .A1(n1307), .A2(n1144), .ZN(n1305) );
  NAND2_X2 U394 ( .A1(n1308), .A2(n1309), .ZN(B[27]) );
  MUX2_X1 U395 ( .A(n1310), .B(n1311), .S(n1137), .Z(n1309) );
  NAND2_X2 U396 ( .A1(n1154), .A2(n1269), .ZN(n1311) );
  NAND2_X2 U397 ( .A1(n1312), .A2(n1313), .ZN(n1269) );
  MUX2_X1 U398 ( .A(n1314), .B(n1315), .S(n1130), .Z(n1313) );
  NAND2_X2 U399 ( .A1(n1122), .A2(n1316), .ZN(n1315) );
  NAND2_X2 U400 ( .A1(n1122), .A2(n1317), .ZN(n1314) );
  MUX2_X1 U401 ( .A(n1318), .B(n1319), .S(n1130), .Z(n1312) );
  NAND2_X2 U402 ( .A1(n1320), .A2(n1110), .ZN(n1319) );
  NAND2_X2 U403 ( .A1(n1321), .A2(n1110), .ZN(n1318) );
  NAND2_X2 U404 ( .A1(n1154), .A2(n1307), .ZN(n1310) );
  MUX2_X1 U405 ( .A(n1322), .B(n1323), .S(n1137), .Z(n1308) );
  NAND2_X2 U406 ( .A1(n1290), .A2(n1144), .ZN(n1323) );
  NAND2_X2 U407 ( .A1(n1324), .A2(n1144), .ZN(n1322) );
  NAND2_X2 U408 ( .A1(n1325), .A2(n1326), .ZN(B[26]) );
  MUX2_X1 U409 ( .A(n1327), .B(n1328), .S(n1137), .Z(n1326) );
  NAND2_X2 U410 ( .A1(n1154), .A2(n1290), .ZN(n1328) );
  NAND2_X2 U411 ( .A1(n1329), .A2(n1330), .ZN(n1290) );
  MUX2_X1 U412 ( .A(n1331), .B(n1332), .S(n1130), .Z(n1330) );
  NAND2_X2 U413 ( .A1(n1121), .A2(n1333), .ZN(n1332) );
  NAND2_X2 U414 ( .A1(n1121), .A2(n1197), .ZN(n1331) );
  MUX2_X1 U415 ( .A(n1334), .B(n1335), .S(n1130), .Z(n1329) );
  NAND2_X2 U416 ( .A1(n1336), .A2(n1110), .ZN(n1335) );
  NAND2_X2 U417 ( .A1(n1193), .A2(n1110), .ZN(n1334) );
  NAND2_X2 U418 ( .A1(n1154), .A2(n1324), .ZN(n1327) );
  MUX2_X1 U419 ( .A(n1337), .B(n1338), .S(n1137), .Z(n1325) );
  NAND2_X2 U420 ( .A1(n1307), .A2(n1144), .ZN(n1338) );
  NAND2_X2 U421 ( .A1(n1339), .A2(n1144), .ZN(n1337) );
  NAND2_X2 U422 ( .A1(n1340), .A2(n1341), .ZN(B[25]) );
  MUX2_X1 U423 ( .A(n1342), .B(n1343), .S(n1137), .Z(n1341) );
  NAND2_X2 U424 ( .A1(n1154), .A2(n1307), .ZN(n1343) );
  NAND2_X2 U425 ( .A1(n1344), .A2(n1345), .ZN(n1307) );
  MUX2_X1 U426 ( .A(n1346), .B(n1347), .S(n1130), .Z(n1345) );
  NAND2_X2 U427 ( .A1(n1121), .A2(n1348), .ZN(n1347) );
  NAND2_X2 U428 ( .A1(n1121), .A2(n1214), .ZN(n1346) );
  MUX2_X1 U429 ( .A(n1349), .B(n1350), .S(n1130), .Z(n1344) );
  NAND2_X2 U430 ( .A1(n1351), .A2(n1109), .ZN(n1350) );
  NAND2_X2 U431 ( .A1(n1210), .A2(n1109), .ZN(n1349) );
  NAND2_X2 U432 ( .A1(n1153), .A2(n1339), .ZN(n1342) );
  MUX2_X1 U433 ( .A(n1352), .B(n1353), .S(n1137), .Z(n1340) );
  NAND2_X2 U434 ( .A1(n1324), .A2(n1143), .ZN(n1353) );
  NAND2_X2 U435 ( .A1(n1355), .A2(n1356), .ZN(B[24]) );
  MUX2_X1 U436 ( .A(n1357), .B(n1358), .S(n1137), .Z(n1356) );
  NAND2_X2 U437 ( .A1(n1153), .A2(n1324), .ZN(n1358) );
  NAND2_X2 U438 ( .A1(n1359), .A2(n1360), .ZN(n1324) );
  MUX2_X1 U439 ( .A(n1361), .B(n1362), .S(n1130), .Z(n1360) );
  NAND2_X2 U440 ( .A1(n1121), .A2(n1300), .ZN(n1362) );
  NAND2_X2 U441 ( .A1(n1120), .A2(n1231), .ZN(n1361) );
  MUX2_X1 U442 ( .A(n1363), .B(n1364), .S(n1130), .Z(n1359) );
  NAND2_X2 U443 ( .A1(n1304), .A2(n1109), .ZN(n1364) );
  NAND2_X2 U444 ( .A1(n1227), .A2(n1109), .ZN(n1363) );
  MUX2_X1 U445 ( .A(n1365), .B(n1366), .S(n1137), .Z(n1355) );
  NAND2_X2 U446 ( .A1(n1339), .A2(n1143), .ZN(n1366) );
  NAND2_X2 U447 ( .A1(n1367), .A2(n1143), .ZN(n1365) );
  MUX2_X1 U448 ( .A(n1370), .B(n1371), .S(n1137), .Z(n1369) );
  NAND2_X2 U449 ( .A1(n1153), .A2(n1339), .ZN(n1371) );
  NAND2_X2 U450 ( .A1(n1372), .A2(n1373), .ZN(n1339) );
  MUX2_X1 U451 ( .A(n1374), .B(n1375), .S(n1130), .Z(n1373) );
  NAND2_X2 U452 ( .A1(n1120), .A2(n1317), .ZN(n1375) );
  NAND2_X2 U453 ( .A1(n1120), .A2(n1248), .ZN(n1374) );
  MUX2_X1 U454 ( .A(n1376), .B(n1377), .S(n1130), .Z(n1372) );
  NAND2_X2 U455 ( .A1(n1321), .A2(n1109), .ZN(n1377) );
  NAND2_X2 U456 ( .A1(n1244), .A2(n1109), .ZN(n1376) );
  NAND2_X2 U457 ( .A1(n1153), .A2(n1367), .ZN(n1370) );
  MUX2_X1 U458 ( .A(n1378), .B(n1379), .S(n1137), .Z(n1368) );
  NAND2_X2 U459 ( .A1(n1380), .A2(n1143), .ZN(n1378) );
  MUX2_X1 U460 ( .A(n1383), .B(n1384), .S(n1137), .Z(n1382) );
  NAND2_X2 U461 ( .A1(n1385), .A2(n1386), .ZN(n1354) );
  MUX2_X1 U462 ( .A(n1387), .B(n1388), .S(n1130), .Z(n1386) );
  NAND2_X2 U463 ( .A1(n1120), .A2(n1197), .ZN(n1388) );
  NAND2_X2 U464 ( .A1(n1120), .A2(n1198), .ZN(n1387) );
  MUX2_X1 U465 ( .A(n1389), .B(n1390), .S(n1130), .Z(n1385) );
  NAND2_X2 U466 ( .A1(n1193), .A2(n1109), .ZN(n1390) );
  NAND2_X2 U467 ( .A1(n1194), .A2(n1109), .ZN(n1389) );
  NAND2_X2 U468 ( .A1(n1152), .A2(n1380), .ZN(n1383) );
  MUX2_X1 U469 ( .A(n1391), .B(n1392), .S(n1137), .Z(n1381) );
  NAND2_X2 U470 ( .A1(n1367), .A2(n1143), .ZN(n1392) );
  NAND2_X2 U471 ( .A1(n1393), .A2(n1143), .ZN(n1391) );
  NAND2_X2 U472 ( .A1(n1394), .A2(n1395), .ZN(B[21]) );
  MUX2_X1 U473 ( .A(n1396), .B(n1397), .S(n1138), .Z(n1395) );
  NAND2_X2 U474 ( .A1(n1152), .A2(n1367), .ZN(n1397) );
  NAND2_X2 U475 ( .A1(n1398), .A2(n1399), .ZN(n1367) );
  MUX2_X1 U476 ( .A(n1400), .B(n1401), .S(n1131), .Z(n1399) );
  NAND2_X2 U477 ( .A1(n1119), .A2(n1214), .ZN(n1401) );
  NAND2_X2 U478 ( .A1(n1119), .A2(n1215), .ZN(n1400) );
  MUX2_X1 U479 ( .A(n1402), .B(n1403), .S(n1131), .Z(n1398) );
  NAND2_X2 U480 ( .A1(n1210), .A2(n1109), .ZN(n1403) );
  NAND2_X2 U481 ( .A1(n1211), .A2(n1109), .ZN(n1402) );
  NAND2_X2 U482 ( .A1(n1152), .A2(n1393), .ZN(n1396) );
  MUX2_X1 U483 ( .A(n1404), .B(n1405), .S(n1138), .Z(n1394) );
  NAND2_X2 U484 ( .A1(n1380), .A2(n1143), .ZN(n1405) );
  NAND2_X2 U485 ( .A1(n1407), .A2(n1408), .ZN(B[20]) );
  MUX2_X1 U486 ( .A(n1409), .B(n1410), .S(n1138), .Z(n1408) );
  NAND2_X2 U487 ( .A1(n1152), .A2(n1380), .ZN(n1410) );
  NAND2_X2 U488 ( .A1(n1411), .A2(n1412), .ZN(n1380) );
  MUX2_X1 U489 ( .A(n1413), .B(n1414), .S(n1131), .Z(n1412) );
  NAND2_X2 U490 ( .A1(n1119), .A2(n1231), .ZN(n1414) );
  NAND2_X2 U491 ( .A1(n1119), .A2(n1232), .ZN(n1413) );
  MUX2_X1 U492 ( .A(n1415), .B(n1416), .S(n1131), .Z(n1411) );
  NAND2_X2 U493 ( .A1(n1227), .A2(n1109), .ZN(n1416) );
  NAND2_X2 U494 ( .A1(n1228), .A2(n1109), .ZN(n1415) );
  MUX2_X1 U495 ( .A(n1417), .B(n1418), .S(n1138), .Z(n1407) );
  NAND2_X2 U496 ( .A1(n1393), .A2(n1143), .ZN(n1418) );
  NAND2_X2 U497 ( .A1(n1419), .A2(n1143), .ZN(n1417) );
  NAND2_X2 U498 ( .A1(n1420), .A2(n1421), .ZN(B[1]) );
  MUX2_X1 U499 ( .A(n1422), .B(n1423), .S(n1138), .Z(n1421) );
  NAND2_X2 U500 ( .A1(n1151), .A2(n1235), .ZN(n1423) );
  NAND2_X2 U501 ( .A1(n1424), .A2(n1425), .ZN(n1235) );
  MUX2_X1 U502 ( .A(n1426), .B(n1427), .S(n1131), .Z(n1425) );
  NAND2_X2 U503 ( .A1(n1119), .A2(n1211), .ZN(n1427) );
  NAND2_X2 U504 ( .A1(n1118), .A2(n1428), .ZN(n1426) );
  MUX2_X1 U505 ( .A(n1429), .B(n1430), .S(n1131), .Z(n1424) );
  NAND2_X2 U506 ( .A1(n1215), .A2(n1108), .ZN(n1430) );
  NAND2_X2 U507 ( .A1(n1431), .A2(n1108), .ZN(n1429) );
  NAND2_X2 U508 ( .A1(n1151), .A2(n1257), .ZN(n1422) );
  MUX2_X1 U509 ( .A(n1432), .B(n1433), .S(n1138), .Z(n1420) );
  NAND2_X2 U510 ( .A1(n1252), .A2(n1142), .ZN(n1433) );
  NAND2_X2 U511 ( .A1(n1261), .A2(n1142), .ZN(n1432) );
  NAND2_X2 U512 ( .A1(n1434), .A2(n1435), .ZN(B[19]) );
  MUX2_X1 U513 ( .A(n1436), .B(n1437), .S(n1138), .Z(n1435) );
  NAND2_X2 U514 ( .A1(n1151), .A2(n1393), .ZN(n1437) );
  NAND2_X2 U515 ( .A1(n1438), .A2(n1439), .ZN(n1393) );
  MUX2_X1 U516 ( .A(n1440), .B(n1441), .S(n1131), .Z(n1439) );
  NAND2_X2 U517 ( .A1(n1118), .A2(n1248), .ZN(n1441) );
  NAND2_X2 U518 ( .A1(n1118), .A2(n1249), .ZN(n1440) );
  MUX2_X1 U519 ( .A(n1442), .B(n1443), .S(n1131), .Z(n1438) );
  NAND2_X2 U520 ( .A1(n1244), .A2(n1108), .ZN(n1443) );
  NAND2_X2 U521 ( .A1(n1245), .A2(n1108), .ZN(n1442) );
  NAND2_X2 U522 ( .A1(n1151), .A2(n1419), .ZN(n1436) );
  MUX2_X1 U523 ( .A(n1444), .B(n1445), .S(n1138), .Z(n1434) );
  NAND2_X2 U524 ( .A1(n1446), .A2(n1142), .ZN(n1444) );
  NAND2_X2 U525 ( .A1(n1447), .A2(n1448), .ZN(B[18]) );
  MUX2_X1 U526 ( .A(n1449), .B(n1450), .S(n1138), .Z(n1448) );
  NAND2_X2 U527 ( .A1(n1451), .A2(n1452), .ZN(n1406) );
  MUX2_X1 U528 ( .A(n1453), .B(n1454), .S(n1131), .Z(n1452) );
  NAND2_X2 U529 ( .A1(n1118), .A2(n1198), .ZN(n1454) );
  INV_X2 U530 ( .A(n1455), .ZN(n1198) );
  MUX2_X1 U531 ( .A(n1456), .B(n1457), .S(n1126), .Z(n1455) );
  NAND2_X2 U532 ( .A1(n1118), .A2(n1281), .ZN(n1453) );
  MUX2_X1 U533 ( .A(n1458), .B(n1459), .S(n1131), .Z(n1451) );
  NAND2_X2 U534 ( .A1(n1194), .A2(n1108), .ZN(n1459) );
  INV_X2 U535 ( .A(n1460), .ZN(n1194) );
  MUX2_X1 U536 ( .A(n1461), .B(n1462), .S(n1126), .Z(n1460) );
  NAND2_X2 U537 ( .A1(n1278), .A2(n1108), .ZN(n1458) );
  NAND2_X2 U538 ( .A1(n1150), .A2(n1446), .ZN(n1449) );
  MUX2_X1 U539 ( .A(n1463), .B(n1464), .S(n1138), .Z(n1447) );
  NAND2_X2 U540 ( .A1(n1419), .A2(n1142), .ZN(n1464) );
  NAND2_X2 U541 ( .A1(n1465), .A2(n1142), .ZN(n1463) );
  NAND2_X2 U542 ( .A1(n1466), .A2(n1467), .ZN(B[17]) );
  MUX2_X1 U543 ( .A(n1468), .B(n1469), .S(n1138), .Z(n1467) );
  NAND2_X2 U544 ( .A1(n1150), .A2(n1419), .ZN(n1469) );
  NAND2_X2 U545 ( .A1(n1470), .A2(n1471), .ZN(n1419) );
  MUX2_X1 U546 ( .A(n1472), .B(n1473), .S(n1131), .Z(n1471) );
  NAND2_X2 U547 ( .A1(n1117), .A2(n1215), .ZN(n1473) );
  INV_X2 U548 ( .A(n1474), .ZN(n1215) );
  MUX2_X1 U549 ( .A(n1475), .B(n1476), .S(n1126), .Z(n1474) );
  NAND2_X2 U550 ( .A1(n1117), .A2(n1431), .ZN(n1472) );
  MUX2_X1 U551 ( .A(n1477), .B(n1478), .S(n1131), .Z(n1470) );
  NAND2_X2 U552 ( .A1(n1211), .A2(n1108), .ZN(n1478) );
  INV_X2 U553 ( .A(n1479), .ZN(n1211) );
  MUX2_X1 U554 ( .A(n1480), .B(n1481), .S(n1126), .Z(n1479) );
  NAND2_X2 U555 ( .A1(n1428), .A2(n1108), .ZN(n1477) );
  NAND2_X2 U556 ( .A1(n1150), .A2(n1465), .ZN(n1468) );
  MUX2_X1 U557 ( .A(n1482), .B(n1483), .S(n1138), .Z(n1466) );
  NAND2_X2 U558 ( .A1(n1446), .A2(n1142), .ZN(n1483) );
  NAND2_X2 U559 ( .A1(n1484), .A2(n1142), .ZN(n1482) );
  NAND2_X2 U560 ( .A1(n1485), .A2(n1486), .ZN(B[16]) );
  MUX2_X1 U561 ( .A(n1487), .B(n1488), .S(n1139), .Z(n1486) );
  NAND2_X2 U562 ( .A1(n1150), .A2(n1446), .ZN(n1488) );
  NAND2_X2 U563 ( .A1(n1489), .A2(n1490), .ZN(n1446) );
  MUX2_X1 U564 ( .A(n1491), .B(n1492), .S(n1132), .Z(n1490) );
  NAND2_X2 U565 ( .A1(n1117), .A2(n1232), .ZN(n1492) );
  NAND2_X2 U566 ( .A1(n1117), .A2(n1303), .ZN(n1491) );
  MUX2_X1 U567 ( .A(n1493), .B(n1494), .S(n1132), .Z(n1489) );
  NAND2_X2 U568 ( .A1(n1228), .A2(n1108), .ZN(n1494) );
  NAND2_X2 U569 ( .A1(n1299), .A2(n1108), .ZN(n1493) );
  NAND2_X2 U570 ( .A1(n1149), .A2(n1484), .ZN(n1487) );
  MUX2_X1 U571 ( .A(n1495), .B(n1496), .S(n1139), .Z(n1485) );
  NAND2_X2 U572 ( .A1(n1465), .A2(n1142), .ZN(n1496) );
  NAND2_X2 U573 ( .A1(n1497), .A2(n1142), .ZN(n1495) );
  NAND2_X2 U574 ( .A1(n1498), .A2(n1499), .ZN(B[15]) );
  MUX2_X1 U575 ( .A(n1500), .B(n1501), .S(n1139), .Z(n1499) );
  NAND2_X2 U576 ( .A1(n1149), .A2(n1465), .ZN(n1501) );
  NAND2_X2 U577 ( .A1(n1502), .A2(n1503), .ZN(n1465) );
  MUX2_X1 U578 ( .A(n1504), .B(n1505), .S(n1132), .Z(n1503) );
  NAND2_X2 U579 ( .A1(n1117), .A2(n1249), .ZN(n1505) );
  NAND2_X2 U580 ( .A1(n1116), .A2(n1320), .ZN(n1504) );
  MUX2_X1 U581 ( .A(n1506), .B(n1507), .S(n1132), .Z(n1502) );
  NAND2_X2 U582 ( .A1(n1245), .A2(n1108), .ZN(n1507) );
  NAND2_X2 U583 ( .A1(n1316), .A2(n1108), .ZN(n1506) );
  NAND2_X2 U584 ( .A1(n1149), .A2(n1497), .ZN(n1500) );
  MUX2_X1 U585 ( .A(n1508), .B(n1509), .S(n1139), .Z(n1498) );
  NAND2_X2 U586 ( .A1(n1484), .A2(n1142), .ZN(n1509) );
  NAND2_X2 U587 ( .A1(n1510), .A2(n1142), .ZN(n1508) );
  NAND2_X2 U588 ( .A1(n1511), .A2(n1512), .ZN(B[14]) );
  MUX2_X1 U589 ( .A(n1513), .B(n1514), .S(n1139), .Z(n1512) );
  NAND2_X2 U590 ( .A1(n1149), .A2(n1484), .ZN(n1514) );
  NAND2_X2 U591 ( .A1(n1515), .A2(n1516), .ZN(n1484) );
  MUX2_X1 U592 ( .A(n1517), .B(n1518), .S(n1132), .Z(n1516) );
  NAND2_X2 U593 ( .A1(n1116), .A2(n1281), .ZN(n1518) );
  NAND2_X2 U594 ( .A1(n1116), .A2(n1336), .ZN(n1517) );
  MUX2_X1 U595 ( .A(n1519), .B(n1520), .S(n1132), .Z(n1515) );
  NAND2_X2 U596 ( .A1(n1278), .A2(n1107), .ZN(n1520) );
  NAND2_X2 U597 ( .A1(n1333), .A2(n1107), .ZN(n1519) );
  NAND2_X2 U598 ( .A1(n1149), .A2(n1510), .ZN(n1513) );
  MUX2_X1 U599 ( .A(n1521), .B(n1522), .S(n1139), .Z(n1511) );
  NAND2_X2 U600 ( .A1(n1497), .A2(n1141), .ZN(n1522) );
  NAND2_X2 U601 ( .A1(n1523), .A2(n1141), .ZN(n1521) );
  NAND2_X2 U602 ( .A1(n1524), .A2(n1525), .ZN(B[13]) );
  MUX2_X1 U603 ( .A(n1526), .B(n1527), .S(n1139), .Z(n1525) );
  NAND2_X2 U604 ( .A1(n1148), .A2(n1497), .ZN(n1527) );
  NAND2_X2 U605 ( .A1(n1528), .A2(n1529), .ZN(n1497) );
  MUX2_X1 U606 ( .A(n1530), .B(n1531), .S(n1132), .Z(n1529) );
  NAND2_X2 U607 ( .A1(n1116), .A2(n1431), .ZN(n1531) );
  NAND2_X2 U608 ( .A1(n1116), .A2(n1351), .ZN(n1530) );
  MUX2_X1 U609 ( .A(n1532), .B(n1533), .S(n1132), .Z(n1528) );
  NAND2_X2 U610 ( .A1(n1428), .A2(n1107), .ZN(n1533) );
  NAND2_X2 U611 ( .A1(n1348), .A2(n1107), .ZN(n1532) );
  NAND2_X2 U612 ( .A1(n1148), .A2(n1523), .ZN(n1526) );
  MUX2_X1 U613 ( .A(n1534), .B(n1535), .S(n1139), .Z(n1524) );
  NAND2_X2 U614 ( .A1(n1510), .A2(n1141), .ZN(n1535) );
  NAND2_X2 U615 ( .A1(n1536), .A2(n1141), .ZN(n1534) );
  NAND2_X2 U616 ( .A1(n1537), .A2(n1538), .ZN(B[12]) );
  MUX2_X1 U617 ( .A(n1539), .B(n1540), .S(n1139), .Z(n1538) );
  NAND2_X2 U618 ( .A1(n1148), .A2(n1510), .ZN(n1540) );
  NAND2_X2 U619 ( .A1(n1541), .A2(n1542), .ZN(n1510) );
  MUX2_X1 U620 ( .A(n1543), .B(n1544), .S(n1132), .Z(n1542) );
  NAND2_X2 U621 ( .A1(n1115), .A2(n1303), .ZN(n1544) );
  NAND2_X2 U622 ( .A1(n1115), .A2(n1304), .ZN(n1543) );
  MUX2_X1 U623 ( .A(n1545), .B(n1546), .S(n1132), .Z(n1541) );
  NAND2_X2 U624 ( .A1(n1299), .A2(n1107), .ZN(n1546) );
  NAND2_X2 U625 ( .A1(n1300), .A2(n1107), .ZN(n1545) );
  NAND2_X2 U626 ( .A1(n1148), .A2(n1536), .ZN(n1539) );
  MUX2_X1 U627 ( .A(n1547), .B(n1548), .S(n1139), .Z(n1537) );
  NAND2_X2 U628 ( .A1(n1523), .A2(n1141), .ZN(n1548) );
  NAND2_X2 U629 ( .A1(n1165), .A2(n1141), .ZN(n1547) );
  NAND2_X2 U630 ( .A1(n1549), .A2(n1550), .ZN(B[11]) );
  MUX2_X1 U631 ( .A(n1551), .B(n1552), .S(n1139), .Z(n1550) );
  NAND2_X2 U632 ( .A1(n1148), .A2(n1523), .ZN(n1552) );
  NAND2_X2 U633 ( .A1(n1553), .A2(n1554), .ZN(n1523) );
  MUX2_X1 U634 ( .A(n1555), .B(n1556), .S(n1132), .Z(n1554) );
  NAND2_X2 U635 ( .A1(n1115), .A2(n1320), .ZN(n1556) );
  NAND2_X2 U636 ( .A1(n1115), .A2(n1321), .ZN(n1555) );
  MUX2_X1 U637 ( .A(n1557), .B(n1558), .S(n1132), .Z(n1553) );
  NAND2_X2 U638 ( .A1(n1316), .A2(n1107), .ZN(n1558) );
  NAND2_X2 U639 ( .A1(n1317), .A2(n1107), .ZN(n1557) );
  NAND2_X2 U640 ( .A1(n1147), .A2(n1165), .ZN(n1551) );
  MUX2_X1 U641 ( .A(n1559), .B(n1560), .S(n1139), .Z(n1549) );
  NAND2_X2 U642 ( .A1(n1536), .A2(n1141), .ZN(n1560) );
  NAND2_X2 U643 ( .A1(n1169), .A2(n1141), .ZN(n1559) );
  NAND2_X2 U644 ( .A1(n1561), .A2(n1562), .ZN(B[10]) );
  MUX2_X1 U645 ( .A(n1563), .B(n1564), .S(n1140), .Z(n1562) );
  NAND2_X2 U646 ( .A1(n1147), .A2(n1536), .ZN(n1564) );
  NAND2_X2 U647 ( .A1(n1565), .A2(n1566), .ZN(n1536) );
  MUX2_X1 U648 ( .A(n1567), .B(n1568), .S(n1133), .Z(n1566) );
  NAND2_X2 U649 ( .A1(n1115), .A2(n1336), .ZN(n1568) );
  NAND2_X2 U650 ( .A1(n1114), .A2(n1193), .ZN(n1567) );
  INV_X2 U651 ( .A(n1569), .ZN(n1193) );
  MUX2_X1 U652 ( .A(n1570), .B(n1571), .S(n1126), .Z(n1569) );
  MUX2_X1 U653 ( .A(n1572), .B(n1573), .S(n1133), .Z(n1565) );
  NAND2_X2 U654 ( .A1(n1333), .A2(n1107), .ZN(n1573) );
  NAND2_X2 U655 ( .A1(n1197), .A2(n1107), .ZN(n1572) );
  INV_X2 U656 ( .A(n1574), .ZN(n1197) );
  MUX2_X1 U657 ( .A(n1575), .B(n1576), .S(n1126), .Z(n1574) );
  NAND2_X2 U658 ( .A1(n1147), .A2(n1169), .ZN(n1563) );
  NAND2_X2 U659 ( .A1(n1577), .A2(n1578), .ZN(n1169) );
  MUX2_X1 U660 ( .A(n1579), .B(n1580), .S(n1133), .Z(n1578) );
  NAND2_X2 U661 ( .A1(n1114), .A2(n1304), .ZN(n1580) );
  INV_X2 U662 ( .A(n1581), .ZN(n1304) );
  MUX2_X1 U663 ( .A(n1582), .B(n1583), .S(n1126), .Z(n1581) );
  NAND2_X2 U664 ( .A1(n1114), .A2(n1227), .ZN(n1579) );
  INV_X2 U665 ( .A(n1584), .ZN(n1227) );
  MUX2_X1 U666 ( .A(n1585), .B(n1586), .S(n1126), .Z(n1584) );
  MUX2_X1 U667 ( .A(n1587), .B(n1588), .S(n1133), .Z(n1577) );
  NAND2_X2 U668 ( .A1(n1300), .A2(n1107), .ZN(n1588) );
  INV_X2 U669 ( .A(n1589), .ZN(n1300) );
  MUX2_X1 U670 ( .A(n1590), .B(n1591), .S(n1126), .Z(n1589) );
  NAND2_X2 U671 ( .A1(n1231), .A2(n1107), .ZN(n1587) );
  INV_X2 U672 ( .A(n1592), .ZN(n1231) );
  MUX2_X1 U673 ( .A(n1593), .B(n1594), .S(n1126), .Z(n1592) );
  MUX2_X1 U674 ( .A(n1595), .B(n1596), .S(n1140), .Z(n1561) );
  NAND2_X2 U675 ( .A1(n1165), .A2(n1141), .ZN(n1596) );
  NAND2_X2 U676 ( .A1(n1597), .A2(n1598), .ZN(n1165) );
  MUX2_X1 U677 ( .A(n1599), .B(n1600), .S(n1133), .Z(n1598) );
  NAND2_X2 U678 ( .A1(n1114), .A2(n1351), .ZN(n1600) );
  NAND2_X2 U679 ( .A1(n1114), .A2(n1210), .ZN(n1599) );
  INV_X2 U680 ( .A(n1601), .ZN(n1210) );
  MUX2_X1 U681 ( .A(n1602), .B(n1603), .S(n1126), .Z(n1601) );
  MUX2_X1 U682 ( .A(n1604), .B(n1605), .S(n1133), .Z(n1597) );
  NAND2_X2 U683 ( .A1(n1348), .A2(n1106), .ZN(n1605) );
  NAND2_X2 U684 ( .A1(n1214), .A2(n1106), .ZN(n1604) );
  INV_X2 U685 ( .A(n1606), .ZN(n1214) );
  MUX2_X1 U686 ( .A(n1607), .B(n1608), .S(n1126), .Z(n1606) );
  NAND2_X2 U687 ( .A1(n1166), .A2(n1141), .ZN(n1595) );
  NAND2_X2 U688 ( .A1(n1609), .A2(n1610), .ZN(n1166) );
  MUX2_X1 U689 ( .A(n1611), .B(n1612), .S(n1133), .Z(n1610) );
  NAND2_X2 U690 ( .A1(n1113), .A2(n1321), .ZN(n1612) );
  INV_X2 U691 ( .A(n1613), .ZN(n1321) );
  MUX2_X1 U692 ( .A(n1614), .B(n1615), .S(n1127), .Z(n1613) );
  NAND2_X2 U693 ( .A1(n1113), .A2(n1244), .ZN(n1611) );
  INV_X2 U694 ( .A(n1616), .ZN(n1244) );
  MUX2_X1 U695 ( .A(n1617), .B(n1618), .S(n1127), .Z(n1616) );
  MUX2_X1 U696 ( .A(n1619), .B(n1620), .S(n1133), .Z(n1609) );
  NAND2_X2 U697 ( .A1(n1317), .A2(n1106), .ZN(n1620) );
  INV_X2 U698 ( .A(n1621), .ZN(n1317) );
  MUX2_X1 U699 ( .A(n1622), .B(n1623), .S(n1127), .Z(n1621) );
  NAND2_X2 U700 ( .A1(n1248), .A2(n1106), .ZN(n1619) );
  INV_X2 U701 ( .A(n1624), .ZN(n1248) );
  MUX2_X1 U702 ( .A(n1625), .B(n1626), .S(n1127), .Z(n1624) );
  NAND2_X2 U703 ( .A1(n1627), .A2(n1628), .ZN(B[0]) );
  MUX2_X1 U704 ( .A(n1629), .B(n1630), .S(n1140), .Z(n1628) );
  NAND2_X2 U705 ( .A1(n1147), .A2(n1252), .ZN(n1630) );
  NAND2_X2 U706 ( .A1(n1631), .A2(n1632), .ZN(n1252) );
  MUX2_X1 U707 ( .A(n1633), .B(n1634), .S(n1133), .Z(n1632) );
  NAND2_X2 U708 ( .A1(n1113), .A2(n1228), .ZN(n1634) );
  INV_X2 U709 ( .A(n1635), .ZN(n1228) );
  MUX2_X1 U710 ( .A(n1591), .B(n1582), .S(n1127), .Z(n1635) );
  NAND2_X2 U711 ( .A1(n1113), .A2(n1299), .ZN(n1633) );
  INV_X2 U712 ( .A(n1636), .ZN(n1299) );
  MUX2_X1 U713 ( .A(n1594), .B(n1585), .S(n1127), .Z(n1636) );
  MUX2_X1 U714 ( .A(n1637), .B(n1638), .S(n1133), .Z(n1631) );
  NAND2_X2 U715 ( .A1(n1232), .A2(n1106), .ZN(n1638) );
  INV_X2 U716 ( .A(n1639), .ZN(n1232) );
  MUX2_X1 U717 ( .A(n1583), .B(n1590), .S(n1127), .Z(n1639) );
  NAND2_X2 U718 ( .A1(n1303), .A2(n1106), .ZN(n1637) );
  INV_X2 U719 ( .A(n1640), .ZN(n1303) );
  MUX2_X1 U720 ( .A(n1586), .B(n1593), .S(n1127), .Z(n1640) );
  NAND2_X2 U721 ( .A1(n1147), .A2(n1261), .ZN(n1629) );
  NAND2_X2 U722 ( .A1(n1641), .A2(n1642), .ZN(n1261) );
  MUX2_X1 U723 ( .A(n1643), .B(n1644), .S(n1133), .Z(n1642) );
  NAND2_X2 U724 ( .A1(n1113), .A2(n1278), .ZN(n1644) );
  INV_X2 U725 ( .A(n1645), .ZN(n1278) );
  NAND2_X2 U726 ( .A1(n1112), .A2(n1333), .ZN(n1643) );
  INV_X2 U727 ( .A(n1646), .ZN(n1333) );
  MUX2_X1 U728 ( .A(n1457), .B(n1461), .S(n1127), .Z(n1646) );
  MUX2_X1 U729 ( .A(n1647), .B(n1648), .S(n1133), .Z(n1641) );
  NAND2_X2 U730 ( .A1(n1281), .A2(n1106), .ZN(n1648) );
  INV_X2 U731 ( .A(n1649), .ZN(n1281) );
  MUX2_X1 U732 ( .A(n1571), .B(n1575), .S(n1127), .Z(n1649) );
  NAND2_X2 U733 ( .A1(n1336), .A2(n1106), .ZN(n1647) );
  INV_X2 U734 ( .A(n1650), .ZN(n1336) );
  MUX2_X1 U735 ( .A(n1462), .B(n1456), .S(n1127), .Z(n1650) );
  MUX2_X1 U736 ( .A(n1651), .B(n1652), .S(n1140), .Z(n1627) );
  NAND2_X2 U737 ( .A1(n1257), .A2(n1141), .ZN(n1652) );
  NAND2_X2 U738 ( .A1(n1653), .A2(n1654), .ZN(n1257) );
  MUX2_X1 U739 ( .A(n1655), .B(n1656), .S(n1134), .Z(n1654) );
  NAND2_X2 U740 ( .A1(n1112), .A2(n1245), .ZN(n1656) );
  INV_X2 U741 ( .A(n1657), .ZN(n1245) );
  MUX2_X1 U742 ( .A(n1623), .B(n1614), .S(n1128), .Z(n1657) );
  NAND2_X2 U743 ( .A1(n1112), .A2(n1316), .ZN(n1655) );
  INV_X2 U744 ( .A(n1658), .ZN(n1316) );
  MUX2_X1 U745 ( .A(n1626), .B(n1617), .S(n1128), .Z(n1658) );
  MUX2_X1 U746 ( .A(n1659), .B(n1660), .S(n1134), .Z(n1653) );
  NAND2_X2 U747 ( .A1(n1249), .A2(n1106), .ZN(n1660) );
  INV_X2 U748 ( .A(n1661), .ZN(n1249) );
  MUX2_X1 U749 ( .A(n1615), .B(n1622), .S(n1128), .Z(n1661) );
  NAND2_X2 U750 ( .A1(n1320), .A2(n1106), .ZN(n1659) );
  INV_X2 U751 ( .A(n1662), .ZN(n1320) );
  MUX2_X1 U752 ( .A(n1618), .B(n1625), .S(n1128), .Z(n1662) );
  NAND2_X2 U753 ( .A1(n1258), .A2(n1141), .ZN(n1651) );
  NAND2_X2 U754 ( .A1(n1663), .A2(n1664), .ZN(n1258) );
  MUX2_X1 U755 ( .A(n1665), .B(n1666), .S(n1134), .Z(n1664) );
  NAND2_X2 U756 ( .A1(n1112), .A2(n1428), .ZN(n1666) );
  INV_X2 U757 ( .A(n1667), .ZN(n1428) );
  MUX2_X1 U758 ( .A(n1608), .B(n1602), .S(n1128), .Z(n1667) );
  NAND2_X2 U759 ( .A1(n1112), .A2(n1348), .ZN(n1665) );
  INV_X2 U760 ( .A(n1668), .ZN(n1348) );
  MUX2_X1 U761 ( .A(n1476), .B(n1480), .S(n1128), .Z(n1668) );
  MUX2_X1 U762 ( .A(n1669), .B(n1670), .S(n1134), .Z(n1663) );
  NAND2_X2 U763 ( .A1(n1431), .A2(n1106), .ZN(n1670) );
  INV_X2 U764 ( .A(n1671), .ZN(n1431) );
  MUX2_X1 U765 ( .A(n1603), .B(n1607), .S(n1128), .Z(n1671) );
  NAND2_X2 U766 ( .A1(n1351), .A2(n1106), .ZN(n1669) );
  INV_X2 U767 ( .A(n1672), .ZN(n1351) );
  MUX2_X1 U768 ( .A(n1481), .B(n1475), .S(n1128), .Z(n1672) );
endmodule


module up_island_DW_sra_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  INV_X4 U170 ( .A(n1130), .ZN(n1121) );
  BUF_X4 U171 ( .A(n1133), .Z(n1130) );
  INV_X1 U172 ( .A(A[30]), .ZN(n1527) );
  INV_X1 U173 ( .A(A[29]), .ZN(n1491) );
  NAND2_X1 U174 ( .A1(n1331), .A2(n1332), .ZN(B[22]) );
  INV_X1 U175 ( .A(A[28]), .ZN(n1502) );
  INV_X1 U176 ( .A(A[4]), .ZN(n1587) );
  INV_X1 U177 ( .A(A[26]), .ZN(n1534) );
  INV_X1 U178 ( .A(A[27]), .ZN(n1518) );
  INV_X1 U179 ( .A(A[23]), .ZN(n1514) );
  INV_X1 U180 ( .A(A[22]), .ZN(n1530) );
  INV_X1 U181 ( .A(A[24]), .ZN(n1409) );
  INV_X1 U182 ( .A(A[25]), .ZN(n1397) );
  OAI21_X1 U183 ( .B1(n1253), .B2(n1111), .A(n1316), .ZN(n1293) );
  NAND2_X1 U184 ( .A1(n1147), .A2(\A[31] ), .ZN(n1280) );
  OAI21_X1 U185 ( .B1(n1253), .B2(n1111), .A(n1307), .ZN(n1283) );
  NAND2_X1 U186 ( .A1(n1152), .A2(\A[31] ), .ZN(n1251) );
  NAND2_X1 U187 ( .A1(n1119), .A2(\A[31] ), .ZN(n1511) );
  NAND2_X1 U188 ( .A1(n1119), .A2(\A[31] ), .ZN(n1498) );
  NAND2_X1 U189 ( .A1(n1120), .A2(\A[31] ), .ZN(n1487) );
  NAND2_X1 U190 ( .A1(n1120), .A2(\A[31] ), .ZN(n1474) );
  MUX2_X2 U191 ( .A(n1518), .B(n1253), .S(n1116), .Z(n1517) );
  INV_X4 U192 ( .A(\A[31] ), .ZN(n1253) );
  INV_X1 U193 ( .A(A[19]), .ZN(n1521) );
  INV_X1 U194 ( .A(A[21]), .ZN(n1494) );
  INV_X1 U195 ( .A(A[15]), .ZN(n1513) );
  INV_X1 U196 ( .A(A[18]), .ZN(n1537) );
  INV_X1 U197 ( .A(A[17]), .ZN(n1265) );
  INV_X1 U198 ( .A(A[13]), .ZN(n1493) );
  INV_X1 U199 ( .A(A[7]), .ZN(n1548) );
  INV_X1 U200 ( .A(A[11]), .ZN(n1520) );
  INV_X1 U201 ( .A(A[20]), .ZN(n1505) );
  INV_X1 U202 ( .A(A[16]), .ZN(n1371) );
  INV_X1 U203 ( .A(A[9]), .ZN(n1264) );
  INV_X1 U204 ( .A(A[12]), .ZN(n1504) );
  INV_X1 U205 ( .A(A[6]), .ZN(n1559) );
  INV_X1 U206 ( .A(A[14]), .ZN(n1529) );
  INV_X1 U207 ( .A(A[8]), .ZN(n1370) );
  INV_X1 U208 ( .A(A[10]), .ZN(n1536) );
  INV_X1 U209 ( .A(A[5]), .ZN(n1572) );
  INV_X1 U210 ( .A(n1112), .ZN(n1106) );
  INV_X1 U211 ( .A(n1112), .ZN(n1107) );
  INV_X1 U212 ( .A(n1112), .ZN(n1108) );
  INV_X1 U213 ( .A(n1112), .ZN(n1109) );
  CLKBUF_X3 U214 ( .A(n1115), .Z(n1110) );
  CLKBUF_X3 U215 ( .A(n1115), .Z(n1111) );
  CLKBUF_X3 U216 ( .A(n1115), .Z(n1112) );
  CLKBUF_X3 U217 ( .A(n1115), .Z(n1113) );
  CLKBUF_X3 U218 ( .A(n1115), .Z(n1114) );
  INV_X8 U219 ( .A(SH[4]), .ZN(n1115) );
  CLKBUF_X3 U220 ( .A(SH[3]), .Z(n1116) );
  CLKBUF_X3 U221 ( .A(SH[3]), .Z(n1117) );
  CLKBUF_X3 U222 ( .A(SH[3]), .Z(n1118) );
  INV_X1 U223 ( .A(n1130), .ZN(n1119) );
  INV_X1 U224 ( .A(n1130), .ZN(n1120) );
  INV_X1 U225 ( .A(n1130), .ZN(n1122) );
  CLKBUF_X3 U226 ( .A(n1133), .Z(n1123) );
  CLKBUF_X3 U227 ( .A(n1133), .Z(n1124) );
  CLKBUF_X3 U228 ( .A(n1133), .Z(n1125) );
  CLKBUF_X3 U229 ( .A(n1133), .Z(n1126) );
  CLKBUF_X3 U230 ( .A(n1133), .Z(n1127) );
  CLKBUF_X3 U231 ( .A(n1133), .Z(n1128) );
  CLKBUF_X3 U232 ( .A(n1133), .Z(n1129) );
  CLKBUF_X3 U233 ( .A(n1133), .Z(n1131) );
  CLKBUF_X3 U234 ( .A(n1133), .Z(n1132) );
  INV_X16 U235 ( .A(SH[2]), .ZN(n1133) );
  INV_X1 U236 ( .A(n1150), .ZN(n1134) );
  INV_X1 U237 ( .A(n1151), .ZN(n1135) );
  INV_X1 U238 ( .A(n1151), .ZN(n1136) );
  INV_X1 U239 ( .A(n1151), .ZN(n1137) );
  INV_X1 U240 ( .A(n1151), .ZN(n1138) );
  CLKBUF_X3 U241 ( .A(SH[1]), .Z(n1139) );
  CLKBUF_X3 U242 ( .A(SH[1]), .Z(n1140) );
  CLKBUF_X3 U243 ( .A(SH[1]), .Z(n1141) );
  CLKBUF_X3 U244 ( .A(SH[1]), .Z(n1142) );
  CLKBUF_X3 U245 ( .A(SH[1]), .Z(n1143) );
  CLKBUF_X3 U246 ( .A(SH[1]), .Z(n1144) );
  CLKBUF_X3 U247 ( .A(SH[1]), .Z(n1145) );
  CLKBUF_X3 U248 ( .A(SH[1]), .Z(n1146) );
  CLKBUF_X3 U249 ( .A(SH[1]), .Z(n1147) );
  CLKBUF_X3 U250 ( .A(SH[1]), .Z(n1148) );
  CLKBUF_X3 U251 ( .A(SH[1]), .Z(n1149) );
  CLKBUF_X3 U252 ( .A(SH[1]), .Z(n1150) );
  CLKBUF_X3 U253 ( .A(SH[1]), .Z(n1151) );
  INV_X1 U254 ( .A(n1157), .ZN(n1152) );
  INV_X1 U255 ( .A(n1157), .ZN(n1153) );
  INV_X1 U256 ( .A(n1156), .ZN(n1154) );
  INV_X1 U257 ( .A(n1157), .ZN(n1155) );
  INV_X1 U258 ( .A(SH[0]), .ZN(n1156) );
  INV_X1 U259 ( .A(SH[0]), .ZN(n1157) );
  NAND2_X2 U260 ( .A1(n1158), .A2(n1159), .ZN(B[9]) );
  MUX2_X1 U261 ( .A(n1160), .B(n1161), .S(n1152), .Z(n1159) );
  NAND2_X2 U262 ( .A1(n1150), .A2(n1162), .ZN(n1161) );
  NAND2_X2 U263 ( .A1(n1150), .A2(n1163), .ZN(n1160) );
  MUX2_X1 U264 ( .A(n1164), .B(n1165), .S(n1155), .Z(n1158) );
  NAND2_X2 U265 ( .A1(n1166), .A2(n1136), .ZN(n1165) );
  NAND2_X2 U266 ( .A1(n1167), .A2(n1134), .ZN(n1164) );
  NAND2_X2 U267 ( .A1(n1168), .A2(n1169), .ZN(B[8]) );
  MUX2_X1 U268 ( .A(n1170), .B(n1171), .S(n1155), .Z(n1169) );
  NAND2_X2 U269 ( .A1(n1150), .A2(n1163), .ZN(n1171) );
  NAND2_X2 U270 ( .A1(n1149), .A2(n1166), .ZN(n1170) );
  MUX2_X1 U271 ( .A(n1172), .B(n1173), .S(n1155), .Z(n1168) );
  NAND2_X2 U272 ( .A1(n1167), .A2(n1134), .ZN(n1173) );
  NAND2_X2 U273 ( .A1(n1174), .A2(n1134), .ZN(n1172) );
  NAND2_X2 U274 ( .A1(n1175), .A2(n1176), .ZN(B[7]) );
  MUX2_X1 U275 ( .A(n1177), .B(n1178), .S(n1155), .Z(n1176) );
  NAND2_X2 U276 ( .A1(n1149), .A2(n1166), .ZN(n1178) );
  NAND2_X2 U277 ( .A1(n1149), .A2(n1167), .ZN(n1177) );
  MUX2_X1 U278 ( .A(n1179), .B(n1180), .S(n1155), .Z(n1175) );
  NAND2_X2 U279 ( .A1(n1174), .A2(n1134), .ZN(n1180) );
  NAND2_X2 U280 ( .A1(n1181), .A2(n1134), .ZN(n1179) );
  NAND2_X2 U281 ( .A1(n1182), .A2(n1183), .ZN(B[6]) );
  MUX2_X1 U282 ( .A(n1184), .B(n1185), .S(n1155), .Z(n1183) );
  NAND2_X2 U283 ( .A1(n1149), .A2(n1167), .ZN(n1185) );
  NAND2_X2 U284 ( .A1(n1186), .A2(n1187), .ZN(n1167) );
  MUX2_X1 U285 ( .A(n1188), .B(n1189), .S(n1106), .Z(n1187) );
  NAND2_X2 U286 ( .A1(n1119), .A2(n1190), .ZN(n1189) );
  NAND2_X2 U287 ( .A1(n1121), .A2(n1191), .ZN(n1188) );
  MUX2_X1 U288 ( .A(n1192), .B(n1193), .S(n1106), .Z(n1186) );
  NAND2_X2 U289 ( .A1(n1194), .A2(n1124), .ZN(n1193) );
  NAND2_X2 U290 ( .A1(n1195), .A2(n1123), .ZN(n1192) );
  NAND2_X2 U291 ( .A1(n1148), .A2(n1174), .ZN(n1184) );
  MUX2_X1 U292 ( .A(n1196), .B(n1197), .S(n1155), .Z(n1182) );
  NAND2_X2 U293 ( .A1(n1181), .A2(n1134), .ZN(n1197) );
  NAND2_X2 U294 ( .A1(n1198), .A2(n1134), .ZN(n1196) );
  NAND2_X2 U295 ( .A1(n1199), .A2(n1200), .ZN(B[5]) );
  MUX2_X1 U296 ( .A(n1201), .B(n1202), .S(n1155), .Z(n1200) );
  NAND2_X2 U297 ( .A1(n1149), .A2(n1174), .ZN(n1202) );
  NAND2_X2 U298 ( .A1(n1203), .A2(n1204), .ZN(n1174) );
  MUX2_X1 U299 ( .A(n1205), .B(n1206), .S(n1106), .Z(n1204) );
  NAND2_X2 U300 ( .A1(n1122), .A2(n1207), .ZN(n1206) );
  NAND2_X2 U301 ( .A1(n1122), .A2(n1208), .ZN(n1205) );
  MUX2_X1 U302 ( .A(n1209), .B(n1210), .S(n1106), .Z(n1203) );
  NAND2_X2 U303 ( .A1(n1211), .A2(n1123), .ZN(n1210) );
  NAND2_X2 U304 ( .A1(n1212), .A2(n1123), .ZN(n1209) );
  NAND2_X2 U305 ( .A1(n1148), .A2(n1181), .ZN(n1201) );
  MUX2_X1 U306 ( .A(n1213), .B(n1214), .S(n1155), .Z(n1199) );
  NAND2_X2 U307 ( .A1(n1198), .A2(n1134), .ZN(n1214) );
  NAND2_X2 U308 ( .A1(n1215), .A2(n1134), .ZN(n1213) );
  NAND2_X2 U309 ( .A1(n1216), .A2(n1217), .ZN(B[4]) );
  MUX2_X1 U310 ( .A(n1218), .B(n1219), .S(n1155), .Z(n1217) );
  NAND2_X2 U311 ( .A1(n1148), .A2(n1181), .ZN(n1219) );
  NAND2_X2 U312 ( .A1(n1220), .A2(n1221), .ZN(n1181) );
  MUX2_X1 U313 ( .A(n1222), .B(n1223), .S(n1106), .Z(n1221) );
  NAND2_X2 U314 ( .A1(n1121), .A2(n1224), .ZN(n1223) );
  NAND2_X2 U315 ( .A1(n1122), .A2(n1225), .ZN(n1222) );
  MUX2_X1 U316 ( .A(n1226), .B(n1227), .S(n1106), .Z(n1220) );
  NAND2_X2 U317 ( .A1(n1228), .A2(n1123), .ZN(n1227) );
  NAND2_X2 U318 ( .A1(n1229), .A2(n1124), .ZN(n1226) );
  NAND2_X2 U319 ( .A1(n1148), .A2(n1198), .ZN(n1218) );
  MUX2_X1 U320 ( .A(n1230), .B(n1231), .S(n1154), .Z(n1216) );
  NAND2_X2 U321 ( .A1(n1215), .A2(n1134), .ZN(n1231) );
  NAND2_X2 U322 ( .A1(n1232), .A2(n1134), .ZN(n1230) );
  NAND2_X2 U323 ( .A1(n1233), .A2(n1234), .ZN(B[3]) );
  MUX2_X1 U324 ( .A(n1235), .B(n1236), .S(n1154), .Z(n1234) );
  NAND2_X2 U325 ( .A1(n1148), .A2(n1198), .ZN(n1236) );
  NAND2_X2 U326 ( .A1(n1237), .A2(n1238), .ZN(n1198) );
  MUX2_X1 U327 ( .A(n1239), .B(n1240), .S(n1106), .Z(n1238) );
  NAND2_X2 U328 ( .A1(n1122), .A2(n1241), .ZN(n1240) );
  NAND2_X2 U329 ( .A1(n1121), .A2(n1242), .ZN(n1239) );
  MUX2_X1 U330 ( .A(n1243), .B(n1244), .S(n1106), .Z(n1237) );
  NAND2_X2 U331 ( .A1(n1245), .A2(n1128), .ZN(n1244) );
  NAND2_X2 U332 ( .A1(n1246), .A2(n1128), .ZN(n1243) );
  NAND2_X2 U333 ( .A1(n1147), .A2(n1215), .ZN(n1235) );
  MUX2_X1 U334 ( .A(n1247), .B(n1248), .S(n1154), .Z(n1233) );
  NAND2_X2 U335 ( .A1(n1232), .A2(n1134), .ZN(n1248) );
  NAND2_X2 U336 ( .A1(n1249), .A2(n1135), .ZN(n1247) );
  NAND2_X2 U337 ( .A1(n1250), .A2(n1251), .ZN(B[30]) );
  MUX2_X1 U338 ( .A(n1252), .B(n1253), .S(n1150), .Z(n1250) );
  NAND2_X2 U339 ( .A1(n1254), .A2(n1156), .ZN(n1252) );
  NAND2_X2 U340 ( .A1(n1255), .A2(n1256), .ZN(B[2]) );
  MUX2_X1 U341 ( .A(n1257), .B(n1258), .S(n1154), .Z(n1256) );
  NAND2_X2 U342 ( .A1(n1147), .A2(n1215), .ZN(n1258) );
  NAND2_X2 U343 ( .A1(n1259), .A2(n1260), .ZN(n1215) );
  MUX2_X1 U344 ( .A(n1261), .B(n1262), .S(n1106), .Z(n1260) );
  NAND2_X2 U345 ( .A1(n1121), .A2(n1194), .ZN(n1262) );
  NAND2_X2 U346 ( .A1(n1121), .A2(n1195), .ZN(n1261) );
  INV_X2 U347 ( .A(n1263), .ZN(n1195) );
  MUX2_X1 U348 ( .A(n1264), .B(n1265), .S(n1116), .Z(n1263) );
  MUX2_X1 U349 ( .A(n1266), .B(n1267), .S(n1106), .Z(n1259) );
  NAND2_X2 U350 ( .A1(n1268), .A2(n1129), .ZN(n1267) );
  NAND2_X2 U351 ( .A1(n1269), .A2(n1129), .ZN(n1266) );
  NAND2_X2 U352 ( .A1(n1147), .A2(n1232), .ZN(n1257) );
  MUX2_X1 U353 ( .A(n1270), .B(n1271), .S(n1154), .Z(n1255) );
  NAND2_X2 U354 ( .A1(n1249), .A2(n1135), .ZN(n1271) );
  NAND2_X2 U355 ( .A1(n1272), .A2(n1135), .ZN(n1270) );
  NAND2_X2 U356 ( .A1(n1273), .A2(n1274), .ZN(B[29]) );
  NAND3_X1 U357 ( .A1(n1156), .A2(n1138), .A3(n1275), .ZN(n1274) );
  MUX2_X1 U358 ( .A(n1276), .B(n1253), .S(n1150), .Z(n1273) );
  NAND2_X2 U359 ( .A1(n1152), .A2(n1254), .ZN(n1276) );
  NAND2_X2 U360 ( .A1(n1277), .A2(n1278), .ZN(B[28]) );
  MUX2_X1 U361 ( .A(n1279), .B(n1280), .S(n1154), .Z(n1278) );
  NAND2_X2 U362 ( .A1(n1147), .A2(n1254), .ZN(n1279) );
  MUX2_X1 U363 ( .A(n1281), .B(n1282), .S(n1154), .Z(n1277) );
  NAND2_X2 U364 ( .A1(n1275), .A2(n1135), .ZN(n1282) );
  NAND2_X2 U365 ( .A1(n1283), .A2(n1135), .ZN(n1281) );
  NAND2_X2 U366 ( .A1(n1284), .A2(n1285), .ZN(B[27]) );
  MUX2_X1 U367 ( .A(n1286), .B(n1287), .S(n1154), .Z(n1285) );
  NAND2_X2 U368 ( .A1(n1146), .A2(n1254), .ZN(n1287) );
  OAI21_X2 U369 ( .B1(n1253), .B2(n1111), .A(n1288), .ZN(n1254) );
  MUX2_X1 U370 ( .A(n1289), .B(n1253), .S(n1122), .Z(n1288) );
  NAND2_X2 U371 ( .A1(n1290), .A2(n1110), .ZN(n1289) );
  NAND2_X2 U372 ( .A1(n1146), .A2(n1275), .ZN(n1286) );
  MUX2_X1 U373 ( .A(n1291), .B(n1292), .S(n1154), .Z(n1284) );
  NAND2_X2 U374 ( .A1(n1283), .A2(n1135), .ZN(n1292) );
  NAND2_X2 U375 ( .A1(n1293), .A2(n1135), .ZN(n1291) );
  NAND2_X2 U376 ( .A1(n1294), .A2(n1295), .ZN(B[26]) );
  MUX2_X1 U377 ( .A(n1296), .B(n1297), .S(n1154), .Z(n1295) );
  NAND2_X2 U378 ( .A1(n1146), .A2(n1275), .ZN(n1297) );
  OAI21_X2 U379 ( .B1(n1253), .B2(n1111), .A(n1298), .ZN(n1275) );
  MUX2_X1 U380 ( .A(n1299), .B(n1253), .S(n1122), .Z(n1298) );
  NAND2_X2 U381 ( .A1(n1190), .A2(n1110), .ZN(n1299) );
  NAND2_X2 U382 ( .A1(n1146), .A2(n1283), .ZN(n1296) );
  MUX2_X1 U383 ( .A(n1300), .B(n1301), .S(n1154), .Z(n1294) );
  NAND2_X2 U384 ( .A1(n1293), .A2(n1135), .ZN(n1301) );
  NAND2_X2 U385 ( .A1(n1302), .A2(n1135), .ZN(n1300) );
  NAND2_X2 U386 ( .A1(n1303), .A2(n1304), .ZN(B[25]) );
  MUX2_X1 U387 ( .A(n1305), .B(n1306), .S(n1154), .Z(n1304) );
  NAND2_X2 U388 ( .A1(n1146), .A2(n1283), .ZN(n1306) );
  MUX2_X1 U389 ( .A(n1308), .B(n1253), .S(n1122), .Z(n1307) );
  NAND2_X2 U390 ( .A1(n1207), .A2(n1110), .ZN(n1308) );
  NAND2_X2 U391 ( .A1(n1145), .A2(n1293), .ZN(n1305) );
  MUX2_X1 U392 ( .A(n1309), .B(n1310), .S(n1154), .Z(n1303) );
  NAND2_X2 U393 ( .A1(n1302), .A2(n1135), .ZN(n1310) );
  NAND2_X2 U394 ( .A1(n1311), .A2(n1135), .ZN(n1309) );
  NAND2_X2 U395 ( .A1(n1312), .A2(n1313), .ZN(B[24]) );
  MUX2_X1 U396 ( .A(n1314), .B(n1315), .S(n1154), .Z(n1313) );
  NAND2_X2 U397 ( .A1(n1145), .A2(n1293), .ZN(n1315) );
  MUX2_X1 U398 ( .A(n1317), .B(n1253), .S(n1122), .Z(n1316) );
  NAND2_X2 U399 ( .A1(n1224), .A2(n1110), .ZN(n1317) );
  NAND2_X2 U400 ( .A1(n1145), .A2(n1302), .ZN(n1314) );
  MUX2_X1 U401 ( .A(n1318), .B(n1319), .S(n1154), .Z(n1312) );
  NAND2_X2 U402 ( .A1(n1311), .A2(n1135), .ZN(n1319) );
  NAND2_X2 U403 ( .A1(n1320), .A2(n1136), .ZN(n1318) );
  NAND2_X2 U404 ( .A1(n1321), .A2(n1322), .ZN(B[23]) );
  MUX2_X1 U405 ( .A(n1323), .B(n1324), .S(n1154), .Z(n1322) );
  NAND2_X2 U406 ( .A1(n1145), .A2(n1302), .ZN(n1324) );
  NAND2_X2 U407 ( .A1(n1325), .A2(n1326), .ZN(n1302) );
  NAND3_X1 U408 ( .A1(n1131), .A2(n1113), .A3(n1241), .ZN(n1326) );
  MUX2_X1 U409 ( .A(n1327), .B(n1253), .S(n1106), .Z(n1325) );
  NAND2_X2 U410 ( .A1(n1121), .A2(n1290), .ZN(n1327) );
  NAND2_X2 U411 ( .A1(n1144), .A2(n1311), .ZN(n1323) );
  MUX2_X1 U412 ( .A(n1328), .B(n1329), .S(n1154), .Z(n1321) );
  NAND2_X2 U413 ( .A1(n1320), .A2(n1136), .ZN(n1329) );
  NAND2_X2 U414 ( .A1(n1330), .A2(n1136), .ZN(n1328) );
  MUX2_X1 U415 ( .A(n1333), .B(n1334), .S(n1153), .Z(n1332) );
  NAND2_X2 U416 ( .A1(n1144), .A2(n1311), .ZN(n1334) );
  NAND2_X2 U417 ( .A1(n1335), .A2(n1336), .ZN(n1311) );
  NAND3_X1 U418 ( .A1(n1131), .A2(n1113), .A3(n1194), .ZN(n1336) );
  MUX2_X1 U419 ( .A(n1337), .B(n1253), .S(n1106), .Z(n1335) );
  NAND2_X2 U420 ( .A1(n1121), .A2(n1190), .ZN(n1337) );
  NAND2_X2 U421 ( .A1(n1144), .A2(n1320), .ZN(n1333) );
  MUX2_X1 U422 ( .A(n1338), .B(n1339), .S(n1153), .Z(n1331) );
  NAND2_X2 U423 ( .A1(n1330), .A2(n1136), .ZN(n1339) );
  NAND2_X2 U424 ( .A1(n1340), .A2(n1136), .ZN(n1338) );
  NAND2_X2 U425 ( .A1(n1341), .A2(n1342), .ZN(B[21]) );
  MUX2_X1 U426 ( .A(n1343), .B(n1344), .S(n1153), .Z(n1342) );
  NAND2_X2 U427 ( .A1(n1144), .A2(n1320), .ZN(n1344) );
  NAND2_X2 U428 ( .A1(n1345), .A2(n1346), .ZN(n1320) );
  NAND3_X1 U429 ( .A1(n1131), .A2(n1112), .A3(n1211), .ZN(n1346) );
  MUX2_X1 U430 ( .A(n1347), .B(n1253), .S(n1107), .Z(n1345) );
  NAND2_X2 U431 ( .A1(n1121), .A2(n1207), .ZN(n1347) );
  NAND2_X2 U432 ( .A1(n1144), .A2(n1330), .ZN(n1343) );
  MUX2_X1 U433 ( .A(n1348), .B(n1349), .S(n1153), .Z(n1341) );
  NAND2_X2 U434 ( .A1(n1340), .A2(n1136), .ZN(n1349) );
  NAND2_X2 U435 ( .A1(n1350), .A2(n1136), .ZN(n1348) );
  NAND2_X2 U436 ( .A1(n1351), .A2(n1352), .ZN(B[20]) );
  MUX2_X1 U437 ( .A(n1353), .B(n1354), .S(n1153), .Z(n1352) );
  NAND2_X2 U438 ( .A1(n1143), .A2(n1330), .ZN(n1354) );
  NAND2_X2 U439 ( .A1(n1355), .A2(n1356), .ZN(n1330) );
  NAND3_X1 U440 ( .A1(n1131), .A2(n1112), .A3(n1228), .ZN(n1356) );
  MUX2_X1 U441 ( .A(n1357), .B(n1253), .S(n1107), .Z(n1355) );
  NAND2_X2 U442 ( .A1(n1121), .A2(n1224), .ZN(n1357) );
  NAND2_X2 U443 ( .A1(n1143), .A2(n1340), .ZN(n1353) );
  MUX2_X1 U444 ( .A(n1358), .B(n1359), .S(n1153), .Z(n1351) );
  NAND2_X2 U445 ( .A1(n1350), .A2(n1136), .ZN(n1359) );
  NAND2_X2 U446 ( .A1(n1360), .A2(n1136), .ZN(n1358) );
  NAND2_X2 U447 ( .A1(n1361), .A2(n1362), .ZN(B[1]) );
  MUX2_X1 U448 ( .A(n1363), .B(n1364), .S(n1153), .Z(n1362) );
  NAND2_X2 U449 ( .A1(n1143), .A2(n1232), .ZN(n1364) );
  NAND2_X2 U450 ( .A1(n1365), .A2(n1366), .ZN(n1232) );
  MUX2_X1 U451 ( .A(n1367), .B(n1368), .S(n1107), .Z(n1366) );
  NAND2_X2 U452 ( .A1(n1121), .A2(n1211), .ZN(n1368) );
  NAND2_X2 U453 ( .A1(n1121), .A2(n1212), .ZN(n1367) );
  INV_X2 U454 ( .A(n1369), .ZN(n1212) );
  MUX2_X1 U455 ( .A(n1370), .B(n1371), .S(n1116), .Z(n1369) );
  MUX2_X1 U456 ( .A(n1372), .B(n1373), .S(n1107), .Z(n1365) );
  NAND2_X2 U457 ( .A1(n1374), .A2(n1129), .ZN(n1373) );
  NAND2_X2 U458 ( .A1(n1375), .A2(n1129), .ZN(n1372) );
  NAND2_X2 U459 ( .A1(n1143), .A2(n1249), .ZN(n1363) );
  MUX2_X1 U460 ( .A(n1376), .B(n1377), .S(n1153), .Z(n1361) );
  NAND2_X2 U461 ( .A1(n1272), .A2(n1136), .ZN(n1377) );
  NAND2_X2 U462 ( .A1(n1378), .A2(n1136), .ZN(n1376) );
  NAND2_X2 U463 ( .A1(n1379), .A2(n1380), .ZN(B[19]) );
  MUX2_X1 U464 ( .A(n1381), .B(n1382), .S(n1153), .Z(n1380) );
  NAND2_X2 U465 ( .A1(n1143), .A2(n1340), .ZN(n1382) );
  NAND2_X2 U466 ( .A1(n1383), .A2(n1384), .ZN(n1340) );
  NAND3_X1 U467 ( .A1(n1130), .A2(n1113), .A3(n1245), .ZN(n1384) );
  MUX2_X1 U468 ( .A(n1385), .B(n1253), .S(n1107), .Z(n1383) );
  NAND2_X2 U469 ( .A1(n1121), .A2(n1241), .ZN(n1385) );
  NAND2_X2 U470 ( .A1(n1142), .A2(n1350), .ZN(n1381) );
  MUX2_X1 U471 ( .A(n1386), .B(n1387), .S(n1153), .Z(n1379) );
  NAND2_X2 U472 ( .A1(n1360), .A2(n1137), .ZN(n1387) );
  NAND2_X2 U473 ( .A1(n1388), .A2(n1137), .ZN(n1386) );
  NAND2_X2 U474 ( .A1(n1389), .A2(n1390), .ZN(B[18]) );
  MUX2_X1 U475 ( .A(n1391), .B(n1392), .S(n1153), .Z(n1390) );
  NAND2_X2 U476 ( .A1(n1142), .A2(n1350), .ZN(n1392) );
  NAND2_X2 U477 ( .A1(n1393), .A2(n1394), .ZN(n1350) );
  NAND3_X1 U478 ( .A1(n1131), .A2(n1112), .A3(n1268), .ZN(n1394) );
  MUX2_X1 U479 ( .A(n1395), .B(n1253), .S(n1107), .Z(n1393) );
  NAND2_X2 U480 ( .A1(n1120), .A2(n1194), .ZN(n1395) );
  INV_X2 U481 ( .A(n1396), .ZN(n1194) );
  MUX2_X1 U482 ( .A(n1397), .B(n1253), .S(n1116), .Z(n1396) );
  NAND2_X2 U483 ( .A1(n1142), .A2(n1360), .ZN(n1391) );
  MUX2_X1 U484 ( .A(n1398), .B(n1399), .S(n1153), .Z(n1389) );
  NAND2_X2 U485 ( .A1(n1388), .A2(n1137), .ZN(n1399) );
  NAND2_X2 U486 ( .A1(n1400), .A2(n1137), .ZN(n1398) );
  NAND2_X2 U487 ( .A1(n1401), .A2(n1402), .ZN(B[17]) );
  MUX2_X1 U488 ( .A(n1403), .B(n1404), .S(n1153), .Z(n1402) );
  NAND2_X2 U489 ( .A1(n1142), .A2(n1360), .ZN(n1404) );
  NAND2_X2 U490 ( .A1(n1405), .A2(n1406), .ZN(n1360) );
  NAND3_X1 U491 ( .A1(n1131), .A2(n1113), .A3(n1374), .ZN(n1406) );
  MUX2_X1 U492 ( .A(n1407), .B(n1253), .S(n1107), .Z(n1405) );
  NAND2_X2 U493 ( .A1(n1120), .A2(n1211), .ZN(n1407) );
  INV_X2 U494 ( .A(n1408), .ZN(n1211) );
  MUX2_X1 U495 ( .A(n1409), .B(n1253), .S(n1116), .Z(n1408) );
  NAND2_X2 U496 ( .A1(n1142), .A2(n1388), .ZN(n1403) );
  MUX2_X1 U497 ( .A(n1410), .B(n1411), .S(n1153), .Z(n1401) );
  NAND2_X2 U498 ( .A1(n1400), .A2(n1137), .ZN(n1411) );
  NAND2_X2 U499 ( .A1(n1412), .A2(n1137), .ZN(n1410) );
  NAND2_X2 U500 ( .A1(n1413), .A2(n1414), .ZN(B[16]) );
  MUX2_X1 U501 ( .A(n1415), .B(n1416), .S(n1153), .Z(n1414) );
  NAND2_X2 U502 ( .A1(n1141), .A2(n1388), .ZN(n1416) );
  NAND2_X2 U503 ( .A1(n1417), .A2(n1418), .ZN(n1388) );
  NAND3_X1 U504 ( .A1(n1132), .A2(n1114), .A3(n1419), .ZN(n1418) );
  MUX2_X1 U505 ( .A(n1420), .B(n1253), .S(n1107), .Z(n1417) );
  NAND2_X2 U506 ( .A1(n1120), .A2(n1228), .ZN(n1420) );
  NAND2_X2 U507 ( .A1(n1141), .A2(n1400), .ZN(n1415) );
  MUX2_X1 U508 ( .A(n1421), .B(n1422), .S(n1152), .Z(n1413) );
  NAND2_X2 U509 ( .A1(n1412), .A2(n1137), .ZN(n1422) );
  NAND2_X2 U510 ( .A1(n1423), .A2(n1137), .ZN(n1421) );
  NAND2_X2 U511 ( .A1(n1424), .A2(n1425), .ZN(B[15]) );
  MUX2_X1 U512 ( .A(n1426), .B(n1427), .S(n1152), .Z(n1425) );
  NAND2_X2 U513 ( .A1(n1141), .A2(n1400), .ZN(n1427) );
  NAND2_X2 U514 ( .A1(n1428), .A2(n1429), .ZN(n1400) );
  NAND3_X1 U515 ( .A1(n1131), .A2(n1113), .A3(n1430), .ZN(n1429) );
  MUX2_X1 U516 ( .A(n1431), .B(n1253), .S(n1107), .Z(n1428) );
  NAND2_X2 U517 ( .A1(n1120), .A2(n1245), .ZN(n1431) );
  NAND2_X2 U518 ( .A1(n1141), .A2(n1412), .ZN(n1426) );
  MUX2_X1 U519 ( .A(n1432), .B(n1433), .S(n1152), .Z(n1424) );
  NAND2_X2 U520 ( .A1(n1423), .A2(n1137), .ZN(n1433) );
  NAND2_X2 U521 ( .A1(n1434), .A2(n1137), .ZN(n1432) );
  NAND2_X2 U522 ( .A1(n1435), .A2(n1436), .ZN(B[14]) );
  MUX2_X1 U523 ( .A(n1437), .B(n1438), .S(n1152), .Z(n1436) );
  NAND2_X2 U524 ( .A1(n1141), .A2(n1412), .ZN(n1438) );
  NAND2_X2 U525 ( .A1(n1439), .A2(n1440), .ZN(n1412) );
  NAND3_X1 U526 ( .A1(n1132), .A2(n1113), .A3(n1441), .ZN(n1440) );
  MUX2_X1 U527 ( .A(n1442), .B(n1253), .S(n1107), .Z(n1439) );
  NAND2_X2 U528 ( .A1(n1120), .A2(n1268), .ZN(n1442) );
  NAND2_X2 U529 ( .A1(n1140), .A2(n1423), .ZN(n1437) );
  MUX2_X1 U530 ( .A(n1443), .B(n1444), .S(n1152), .Z(n1435) );
  NAND2_X2 U531 ( .A1(n1434), .A2(n1137), .ZN(n1444) );
  NAND2_X2 U532 ( .A1(n1445), .A2(n1137), .ZN(n1443) );
  NAND2_X2 U533 ( .A1(n1446), .A2(n1447), .ZN(B[13]) );
  MUX2_X1 U534 ( .A(n1448), .B(n1449), .S(n1152), .Z(n1447) );
  NAND2_X2 U535 ( .A1(n1140), .A2(n1423), .ZN(n1449) );
  NAND2_X2 U536 ( .A1(n1450), .A2(n1451), .ZN(n1423) );
  NAND3_X1 U537 ( .A1(n1132), .A2(n1113), .A3(n1452), .ZN(n1451) );
  MUX2_X1 U538 ( .A(n1453), .B(n1253), .S(n1107), .Z(n1450) );
  NAND2_X2 U539 ( .A1(n1120), .A2(n1374), .ZN(n1453) );
  NAND2_X2 U540 ( .A1(n1140), .A2(n1434), .ZN(n1448) );
  MUX2_X1 U541 ( .A(n1454), .B(n1455), .S(n1152), .Z(n1446) );
  NAND2_X2 U542 ( .A1(n1445), .A2(n1138), .ZN(n1455) );
  NAND2_X2 U543 ( .A1(n1456), .A2(n1138), .ZN(n1454) );
  NAND2_X2 U544 ( .A1(n1457), .A2(n1458), .ZN(B[12]) );
  MUX2_X1 U545 ( .A(n1459), .B(n1460), .S(n1152), .Z(n1458) );
  NAND2_X2 U546 ( .A1(n1140), .A2(n1434), .ZN(n1460) );
  NAND2_X2 U547 ( .A1(n1461), .A2(n1462), .ZN(n1434) );
  NAND3_X1 U548 ( .A1(n1132), .A2(n1114), .A3(n1463), .ZN(n1462) );
  MUX2_X1 U549 ( .A(n1464), .B(n1253), .S(n1107), .Z(n1461) );
  NAND2_X2 U550 ( .A1(n1120), .A2(n1419), .ZN(n1464) );
  NAND2_X2 U551 ( .A1(n1140), .A2(n1445), .ZN(n1459) );
  MUX2_X1 U552 ( .A(n1465), .B(n1466), .S(n1152), .Z(n1457) );
  NAND2_X2 U553 ( .A1(n1456), .A2(n1138), .ZN(n1466) );
  NAND2_X2 U554 ( .A1(n1162), .A2(n1138), .ZN(n1465) );
  NAND2_X2 U555 ( .A1(n1467), .A2(n1468), .ZN(B[11]) );
  MUX2_X1 U556 ( .A(n1469), .B(n1470), .S(n1152), .Z(n1468) );
  NAND2_X2 U557 ( .A1(n1139), .A2(n1445), .ZN(n1470) );
  NAND2_X2 U558 ( .A1(n1471), .A2(n1472), .ZN(n1445) );
  MUX2_X1 U559 ( .A(n1473), .B(n1474), .S(n1108), .Z(n1472) );
  NAND2_X2 U560 ( .A1(n1120), .A2(n1430), .ZN(n1473) );
  MUX2_X1 U561 ( .A(n1475), .B(n1476), .S(n1108), .Z(n1471) );
  NAND2_X2 U562 ( .A1(n1290), .A2(n1128), .ZN(n1476) );
  NAND2_X2 U563 ( .A1(n1477), .A2(n1128), .ZN(n1475) );
  NAND2_X2 U564 ( .A1(n1139), .A2(n1456), .ZN(n1469) );
  MUX2_X1 U565 ( .A(n1478), .B(n1479), .S(n1153), .Z(n1467) );
  NAND2_X2 U566 ( .A1(n1162), .A2(n1138), .ZN(n1479) );
  NAND2_X2 U567 ( .A1(n1163), .A2(n1138), .ZN(n1478) );
  NAND2_X2 U568 ( .A1(n1480), .A2(n1481), .ZN(B[10]) );
  MUX2_X1 U569 ( .A(n1482), .B(n1483), .S(n1152), .Z(n1481) );
  NAND2_X2 U570 ( .A1(n1139), .A2(n1456), .ZN(n1483) );
  NAND2_X2 U571 ( .A1(n1484), .A2(n1485), .ZN(n1456) );
  MUX2_X1 U572 ( .A(n1486), .B(n1487), .S(n1108), .Z(n1485) );
  NAND2_X2 U573 ( .A1(n1120), .A2(n1441), .ZN(n1486) );
  MUX2_X1 U574 ( .A(n1488), .B(n1489), .S(n1108), .Z(n1484) );
  NAND2_X2 U575 ( .A1(n1190), .A2(n1127), .ZN(n1489) );
  INV_X2 U576 ( .A(n1490), .ZN(n1190) );
  MUX2_X1 U577 ( .A(n1491), .B(n1253), .S(n1116), .Z(n1490) );
  NAND2_X2 U578 ( .A1(n1191), .A2(n1127), .ZN(n1488) );
  INV_X2 U579 ( .A(n1492), .ZN(n1191) );
  MUX2_X1 U580 ( .A(n1493), .B(n1494), .S(n1116), .Z(n1492) );
  NAND2_X2 U581 ( .A1(n1139), .A2(n1162), .ZN(n1482) );
  NAND2_X2 U582 ( .A1(n1495), .A2(n1496), .ZN(n1162) );
  MUX2_X1 U583 ( .A(n1497), .B(n1498), .S(n1108), .Z(n1496) );
  NAND2_X2 U584 ( .A1(n1119), .A2(n1452), .ZN(n1497) );
  MUX2_X1 U585 ( .A(n1499), .B(n1500), .S(n1108), .Z(n1495) );
  NAND2_X2 U586 ( .A1(n1207), .A2(n1127), .ZN(n1500) );
  INV_X2 U587 ( .A(n1501), .ZN(n1207) );
  MUX2_X1 U588 ( .A(n1502), .B(n1253), .S(n1116), .Z(n1501) );
  NAND2_X2 U589 ( .A1(n1208), .A2(n1127), .ZN(n1499) );
  INV_X2 U590 ( .A(n1503), .ZN(n1208) );
  MUX2_X1 U591 ( .A(n1504), .B(n1505), .S(n1116), .Z(n1503) );
  MUX2_X1 U592 ( .A(n1506), .B(n1507), .S(n1152), .Z(n1480) );
  NAND2_X2 U593 ( .A1(n1163), .A2(n1138), .ZN(n1507) );
  NAND2_X2 U594 ( .A1(n1508), .A2(n1509), .ZN(n1163) );
  MUX2_X1 U595 ( .A(n1510), .B(n1511), .S(n1108), .Z(n1509) );
  NAND2_X2 U596 ( .A1(n1120), .A2(n1463), .ZN(n1510) );
  INV_X2 U597 ( .A(n1512), .ZN(n1463) );
  MUX2_X1 U598 ( .A(n1513), .B(n1514), .S(n1116), .Z(n1512) );
  MUX2_X1 U599 ( .A(n1515), .B(n1516), .S(n1108), .Z(n1508) );
  NAND2_X2 U600 ( .A1(n1224), .A2(n1126), .ZN(n1516) );
  INV_X2 U601 ( .A(n1517), .ZN(n1224) );
  NAND2_X2 U602 ( .A1(n1225), .A2(n1126), .ZN(n1515) );
  INV_X2 U603 ( .A(n1519), .ZN(n1225) );
  MUX2_X1 U604 ( .A(n1520), .B(n1521), .S(n1116), .Z(n1519) );
  NAND2_X2 U605 ( .A1(n1166), .A2(n1138), .ZN(n1506) );
  NAND2_X2 U606 ( .A1(n1522), .A2(n1523), .ZN(n1166) );
  MUX2_X1 U607 ( .A(n1524), .B(n1525), .S(n1108), .Z(n1523) );
  NAND2_X2 U608 ( .A1(n1119), .A2(n1290), .ZN(n1525) );
  INV_X2 U609 ( .A(n1526), .ZN(n1290) );
  MUX2_X1 U610 ( .A(n1527), .B(n1253), .S(n1116), .Z(n1526) );
  NAND2_X2 U611 ( .A1(n1119), .A2(n1477), .ZN(n1524) );
  INV_X2 U612 ( .A(n1528), .ZN(n1477) );
  MUX2_X1 U613 ( .A(n1529), .B(n1530), .S(n1117), .Z(n1528) );
  MUX2_X1 U614 ( .A(n1531), .B(n1532), .S(n1108), .Z(n1522) );
  NAND2_X2 U615 ( .A1(n1241), .A2(n1126), .ZN(n1532) );
  INV_X2 U616 ( .A(n1533), .ZN(n1241) );
  MUX2_X1 U617 ( .A(n1534), .B(n1253), .S(n1117), .Z(n1533) );
  NAND2_X2 U618 ( .A1(n1242), .A2(n1126), .ZN(n1531) );
  INV_X2 U619 ( .A(n1535), .ZN(n1242) );
  MUX2_X1 U620 ( .A(n1536), .B(n1537), .S(n1117), .Z(n1535) );
  NAND2_X2 U621 ( .A1(n1538), .A2(n1539), .ZN(B[0]) );
  MUX2_X1 U622 ( .A(n1540), .B(n1541), .S(n1152), .Z(n1539) );
  NAND2_X2 U623 ( .A1(n1139), .A2(n1249), .ZN(n1541) );
  NAND2_X2 U624 ( .A1(n1542), .A2(n1543), .ZN(n1249) );
  MUX2_X1 U625 ( .A(n1544), .B(n1545), .S(n1108), .Z(n1543) );
  NAND2_X2 U626 ( .A1(n1119), .A2(n1228), .ZN(n1545) );
  INV_X2 U627 ( .A(n1546), .ZN(n1228) );
  MUX2_X1 U628 ( .A(n1514), .B(n1253), .S(n1117), .Z(n1546) );
  NAND2_X2 U629 ( .A1(n1119), .A2(n1229), .ZN(n1544) );
  INV_X2 U630 ( .A(n1547), .ZN(n1229) );
  MUX2_X1 U631 ( .A(n1548), .B(n1513), .S(n1117), .Z(n1547) );
  MUX2_X1 U632 ( .A(n1549), .B(n1550), .S(n1108), .Z(n1542) );
  NAND2_X2 U633 ( .A1(n1419), .A2(n1125), .ZN(n1550) );
  INV_X2 U634 ( .A(n1551), .ZN(n1419) );
  MUX2_X1 U635 ( .A(n1521), .B(n1518), .S(n1117), .Z(n1551) );
  NAND2_X2 U636 ( .A1(n1552), .A2(n1125), .ZN(n1549) );
  MUX2_X1 U637 ( .A(A[3]), .B(A[11]), .S(n1117), .Z(n1552) );
  NAND2_X2 U638 ( .A1(n1145), .A2(n1272), .ZN(n1540) );
  NAND2_X2 U639 ( .A1(n1553), .A2(n1554), .ZN(n1272) );
  MUX2_X1 U640 ( .A(n1555), .B(n1556), .S(n1109), .Z(n1554) );
  NAND2_X2 U641 ( .A1(n1119), .A2(n1245), .ZN(n1556) );
  INV_X2 U642 ( .A(n1557), .ZN(n1245) );
  MUX2_X1 U643 ( .A(n1530), .B(n1527), .S(n1117), .Z(n1557) );
  NAND2_X2 U644 ( .A1(n1119), .A2(n1246), .ZN(n1555) );
  INV_X2 U645 ( .A(n1558), .ZN(n1246) );
  MUX2_X1 U646 ( .A(n1559), .B(n1529), .S(n1117), .Z(n1558) );
  MUX2_X1 U647 ( .A(n1560), .B(n1561), .S(n1109), .Z(n1553) );
  NAND2_X2 U648 ( .A1(n1430), .A2(n1125), .ZN(n1561) );
  INV_X2 U649 ( .A(n1562), .ZN(n1430) );
  MUX2_X1 U650 ( .A(n1537), .B(n1534), .S(n1117), .Z(n1562) );
  NAND2_X2 U651 ( .A1(n1563), .A2(n1125), .ZN(n1560) );
  MUX2_X1 U652 ( .A(A[2]), .B(A[10]), .S(n1117), .Z(n1563) );
  MUX2_X1 U653 ( .A(n1564), .B(n1565), .S(n1153), .Z(n1538) );
  NAND2_X2 U654 ( .A1(n1378), .A2(n1138), .ZN(n1565) );
  NAND2_X2 U655 ( .A1(n1566), .A2(n1567), .ZN(n1378) );
  MUX2_X1 U656 ( .A(n1568), .B(n1569), .S(n1109), .Z(n1567) );
  NAND2_X2 U657 ( .A1(n1119), .A2(n1268), .ZN(n1569) );
  INV_X2 U658 ( .A(n1570), .ZN(n1268) );
  MUX2_X1 U659 ( .A(n1494), .B(n1491), .S(n1117), .Z(n1570) );
  NAND2_X2 U660 ( .A1(n1119), .A2(n1269), .ZN(n1568) );
  INV_X2 U661 ( .A(n1571), .ZN(n1269) );
  MUX2_X1 U662 ( .A(n1572), .B(n1493), .S(n1118), .Z(n1571) );
  MUX2_X1 U663 ( .A(n1573), .B(n1574), .S(n1109), .Z(n1566) );
  NAND2_X2 U664 ( .A1(n1441), .A2(n1124), .ZN(n1574) );
  INV_X2 U665 ( .A(n1575), .ZN(n1441) );
  MUX2_X1 U666 ( .A(n1265), .B(n1397), .S(n1118), .Z(n1575) );
  NAND2_X2 U667 ( .A1(n1576), .A2(n1124), .ZN(n1573) );
  MUX2_X1 U668 ( .A(A[1]), .B(A[9]), .S(n1118), .Z(n1576) );
  OAI21_X2 U669 ( .B1(n1577), .B2(n1578), .A(n1138), .ZN(n1564) );
  MUX2_X1 U670 ( .A(n1579), .B(n1580), .S(n1109), .Z(n1578) );
  AND2_X2 U671 ( .A1(n1452), .A2(n1130), .ZN(n1580) );
  INV_X2 U672 ( .A(n1581), .ZN(n1452) );
  MUX2_X1 U673 ( .A(n1371), .B(n1409), .S(n1118), .Z(n1581) );
  AND2_X2 U674 ( .A1(n1582), .A2(n1130), .ZN(n1579) );
  MUX2_X1 U675 ( .A(A[0]), .B(A[8]), .S(n1118), .Z(n1582) );
  MUX2_X1 U676 ( .A(n1583), .B(n1584), .S(n1109), .Z(n1577) );
  AND2_X2 U677 ( .A1(n1122), .A2(n1374), .ZN(n1584) );
  INV_X2 U678 ( .A(n1585), .ZN(n1374) );
  MUX2_X1 U679 ( .A(n1505), .B(n1502), .S(n1118), .Z(n1585) );
  AND2_X2 U680 ( .A1(n1122), .A2(n1375), .ZN(n1583) );
  INV_X2 U681 ( .A(n1586), .ZN(n1375) );
  MUX2_X1 U682 ( .A(n1587), .B(n1504), .S(n1118), .Z(n1586) );
endmodule


module up_island_DW_rightsh_1 ( A, SH, B, DATA_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633;

  NAND2_X1 U108 ( .A1(A[29]), .A2(n1180), .ZN(n1535) );
  INV_X1 U109 ( .A(A[29]), .ZN(n1584) );
  INV_X1 U110 ( .A(A[2]), .ZN(n1626) );
  INV_X4 U111 ( .A(SH[2]), .ZN(n1186) );
  NAND2_X1 U112 ( .A1(A[30]), .A2(n1179), .ZN(n1530) );
  INV_X1 U113 ( .A(A[30]), .ZN(n1588) );
  INV_X1 U114 ( .A(A[1]), .ZN(n1633) );
  INV_X1 U115 ( .A(A[28]), .ZN(n1590) );
  NAND2_X1 U116 ( .A1(A[28]), .A2(n1181), .ZN(n1539) );
  INV_X1 U117 ( .A(A[3]), .ZN(n1631) );
  INV_X1 U118 ( .A(A[4]), .ZN(n1620) );
  NAND2_X1 U119 ( .A1(A[26]), .A2(n1181), .ZN(n1540) );
  INV_X1 U120 ( .A(A[26]), .ZN(n1602) );
  NAND2_X1 U121 ( .A1(A[27]), .A2(n1180), .ZN(n1536) );
  INV_X1 U122 ( .A(A[27]), .ZN(n1596) );
  INV_X1 U123 ( .A(A[23]), .ZN(n1549) );
  INV_X1 U124 ( .A(A[22]), .ZN(n1554) );
  INV_X1 U125 ( .A(A[24]), .ZN(n1604) );
  NAND2_X1 U126 ( .A1(A[24]), .A2(n1178), .ZN(n1420) );
  INV_X1 U127 ( .A(A[25]), .ZN(n1598) );
  NAND2_X1 U128 ( .A1(A[25]), .A2(n1178), .ZN(n1410) );
  INV_X1 U129 ( .A(A[31]), .ZN(n1582) );
  NAND2_X1 U130 ( .A1(A[31]), .A2(n1179), .ZN(n1528) );
  INV_X1 U131 ( .A(A[19]), .ZN(n1564) );
  INV_X1 U132 ( .A(A[21]), .ZN(n1561) );
  INV_X1 U133 ( .A(A[15]), .ZN(n1548) );
  INV_X1 U134 ( .A(A[18]), .ZN(n1572) );
  INV_X1 U135 ( .A(A[17]), .ZN(n1324) );
  INV_X1 U136 ( .A(A[13]), .ZN(n1560) );
  INV_X1 U137 ( .A(A[7]), .ZN(n1612) );
  INV_X1 U138 ( .A(A[11]), .ZN(n1563) );
  INV_X1 U139 ( .A(A[20]), .ZN(n1569) );
  INV_X1 U140 ( .A(A[16]), .ZN(n1385) );
  INV_X1 U141 ( .A(A[9]), .ZN(n1323) );
  INV_X1 U142 ( .A(A[12]), .ZN(n1568) );
  INV_X1 U143 ( .A(A[6]), .ZN(n1618) );
  INV_X1 U144 ( .A(A[14]), .ZN(n1553) );
  INV_X1 U145 ( .A(A[8]), .ZN(n1384) );
  INV_X1 U146 ( .A(A[10]), .ZN(n1571) );
  INV_X1 U147 ( .A(A[5]), .ZN(n1614) );
  INV_X1 U148 ( .A(n1168), .ZN(n1163) );
  INV_X1 U149 ( .A(n1173), .ZN(n1164) );
  INV_X1 U150 ( .A(n1174), .ZN(n1165) );
  INV_X1 U151 ( .A(n1175), .ZN(n1166) );
  CLKBUF_X3 U152 ( .A(SH[4]), .Z(n1167) );
  CLKBUF_X3 U153 ( .A(SH[4]), .Z(n1168) );
  CLKBUF_X3 U154 ( .A(SH[4]), .Z(n1169) );
  CLKBUF_X3 U155 ( .A(SH[4]), .Z(n1170) );
  CLKBUF_X3 U156 ( .A(SH[4]), .Z(n1171) );
  CLKBUF_X3 U157 ( .A(SH[4]), .Z(n1172) );
  CLKBUF_X3 U158 ( .A(SH[4]), .Z(n1173) );
  CLKBUF_X3 U159 ( .A(SH[4]), .Z(n1174) );
  CLKBUF_X3 U160 ( .A(SH[4]), .Z(n1175) );
  INV_X1 U161 ( .A(n1182), .ZN(n1176) );
  INV_X1 U162 ( .A(n1182), .ZN(n1177) );
  INV_X1 U163 ( .A(SH[3]), .ZN(n1178) );
  INV_X1 U164 ( .A(SH[3]), .ZN(n1179) );
  INV_X1 U165 ( .A(SH[3]), .ZN(n1180) );
  INV_X1 U166 ( .A(SH[3]), .ZN(n1181) );
  INV_X1 U167 ( .A(SH[3]), .ZN(n1182) );
  INV_X1 U168 ( .A(n1186), .ZN(n1183) );
  INV_X1 U169 ( .A(n1186), .ZN(n1184) );
  INV_X1 U170 ( .A(n1186), .ZN(n1185) );
  INV_X1 U171 ( .A(n1192), .ZN(n1187) );
  INV_X1 U172 ( .A(n1192), .ZN(n1188) );
  INV_X1 U173 ( .A(n1192), .ZN(n1189) );
  INV_X1 U174 ( .A(n1192), .ZN(n1190) );
  INV_X2 U175 ( .A(SH[1]), .ZN(n1191) );
  INV_X2 U176 ( .A(SH[1]), .ZN(n1192) );
  INV_X1 U177 ( .A(n1206), .ZN(n1193) );
  INV_X1 U178 ( .A(n1204), .ZN(n1194) );
  INV_X1 U179 ( .A(n1207), .ZN(n1195) );
  INV_X1 U180 ( .A(n1205), .ZN(n1196) );
  INV_X1 U181 ( .A(n1203), .ZN(n1197) );
  CLKBUF_X3 U182 ( .A(SH[0]), .Z(n1198) );
  CLKBUF_X3 U183 ( .A(SH[0]), .Z(n1199) );
  CLKBUF_X3 U184 ( .A(SH[0]), .Z(n1200) );
  CLKBUF_X3 U185 ( .A(SH[0]), .Z(n1201) );
  CLKBUF_X3 U186 ( .A(SH[0]), .Z(n1202) );
  CLKBUF_X3 U187 ( .A(SH[0]), .Z(n1203) );
  CLKBUF_X3 U188 ( .A(SH[0]), .Z(n1204) );
  CLKBUF_X3 U189 ( .A(SH[0]), .Z(n1205) );
  CLKBUF_X3 U190 ( .A(SH[0]), .Z(n1206) );
  CLKBUF_X3 U191 ( .A(SH[0]), .Z(n1207) );
  CLKBUF_X3 U192 ( .A(SH[0]), .Z(n1208) );
  CLKBUF_X3 U193 ( .A(SH[0]), .Z(n1209) );
  CLKBUF_X3 U194 ( .A(SH[0]), .Z(n1210) );
  CLKBUF_X3 U195 ( .A(SH[0]), .Z(n1211) );
  NAND2_X2 U196 ( .A1(n1212), .A2(n1213), .ZN(B[9]) );
  MUX2_X1 U197 ( .A(n1214), .B(n1215), .S(n1183), .Z(n1213) );
  NAND2_X2 U198 ( .A1(n1174), .A2(n1216), .ZN(n1215) );
  NAND2_X2 U199 ( .A1(n1175), .A2(n1217), .ZN(n1214) );
  MUX2_X1 U200 ( .A(n1218), .B(n1219), .S(n1185), .Z(n1212) );
  NAND2_X2 U201 ( .A1(n1220), .A2(n1163), .ZN(n1219) );
  NAND2_X2 U202 ( .A1(n1221), .A2(n1163), .ZN(n1218) );
  NAND2_X2 U203 ( .A1(n1222), .A2(n1223), .ZN(B[8]) );
  MUX2_X1 U204 ( .A(n1224), .B(n1225), .S(n1185), .Z(n1223) );
  NAND2_X2 U205 ( .A1(n1174), .A2(n1226), .ZN(n1225) );
  NAND2_X2 U206 ( .A1(n1174), .A2(n1227), .ZN(n1224) );
  MUX2_X1 U207 ( .A(n1228), .B(n1229), .S(n1185), .Z(n1222) );
  NAND2_X2 U208 ( .A1(n1230), .A2(n1163), .ZN(n1229) );
  NAND2_X2 U209 ( .A1(n1231), .A2(n1163), .ZN(n1228) );
  NAND2_X2 U210 ( .A1(n1232), .A2(n1233), .ZN(B[7]) );
  MUX2_X1 U211 ( .A(n1234), .B(n1235), .S(n1185), .Z(n1233) );
  NAND2_X2 U212 ( .A1(n1174), .A2(n1236), .ZN(n1235) );
  NAND2_X2 U213 ( .A1(n1173), .A2(n1237), .ZN(n1234) );
  MUX2_X1 U214 ( .A(n1238), .B(n1239), .S(n1185), .Z(n1232) );
  NAND2_X2 U215 ( .A1(n1240), .A2(n1163), .ZN(n1239) );
  NAND2_X2 U216 ( .A1(n1241), .A2(n1163), .ZN(n1238) );
  NAND2_X2 U217 ( .A1(n1242), .A2(n1243), .ZN(B[6]) );
  MUX2_X1 U218 ( .A(n1244), .B(n1245), .S(n1185), .Z(n1243) );
  NAND2_X2 U219 ( .A1(n1173), .A2(n1246), .ZN(n1245) );
  NAND2_X2 U220 ( .A1(n1173), .A2(n1247), .ZN(n1244) );
  MUX2_X1 U221 ( .A(n1248), .B(n1249), .S(n1185), .Z(n1242) );
  NAND2_X2 U222 ( .A1(n1250), .A2(n1163), .ZN(n1249) );
  NAND2_X2 U223 ( .A1(n1251), .A2(n1164), .ZN(n1248) );
  NAND2_X2 U224 ( .A1(n1252), .A2(n1253), .ZN(B[5]) );
  MUX2_X1 U225 ( .A(n1254), .B(n1255), .S(n1185), .Z(n1253) );
  NAND2_X2 U226 ( .A1(n1173), .A2(n1217), .ZN(n1255) );
  NAND2_X2 U227 ( .A1(n1172), .A2(n1256), .ZN(n1254) );
  MUX2_X1 U228 ( .A(n1257), .B(n1258), .S(n1184), .Z(n1252) );
  NAND2_X2 U229 ( .A1(n1221), .A2(n1164), .ZN(n1258) );
  NAND2_X2 U230 ( .A1(n1259), .A2(n1260), .ZN(n1221) );
  MUX2_X1 U231 ( .A(n1261), .B(n1262), .S(n1187), .Z(n1260) );
  NAND2_X2 U232 ( .A1(n1209), .A2(n1263), .ZN(n1262) );
  NAND2_X2 U233 ( .A1(n1210), .A2(n1264), .ZN(n1261) );
  MUX2_X1 U234 ( .A(n1265), .B(n1266), .S(n1190), .Z(n1259) );
  NAND2_X2 U235 ( .A1(n1267), .A2(n1195), .ZN(n1266) );
  NAND2_X2 U236 ( .A1(n1268), .A2(n1193), .ZN(n1265) );
  NAND2_X2 U237 ( .A1(n1269), .A2(n1164), .ZN(n1257) );
  NAND2_X2 U238 ( .A1(n1270), .A2(n1271), .ZN(B[4]) );
  MUX2_X1 U239 ( .A(n1272), .B(n1273), .S(n1184), .Z(n1271) );
  NAND2_X2 U240 ( .A1(n1172), .A2(n1227), .ZN(n1273) );
  NAND2_X2 U241 ( .A1(n1172), .A2(n1274), .ZN(n1272) );
  MUX2_X1 U242 ( .A(n1275), .B(n1276), .S(n1184), .Z(n1270) );
  NAND2_X2 U243 ( .A1(n1231), .A2(n1164), .ZN(n1276) );
  NAND2_X2 U244 ( .A1(n1277), .A2(n1278), .ZN(n1231) );
  MUX2_X1 U245 ( .A(n1279), .B(n1280), .S(n1190), .Z(n1278) );
  NAND2_X2 U246 ( .A1(n1209), .A2(n1267), .ZN(n1280) );
  NAND2_X2 U247 ( .A1(n1210), .A2(n1268), .ZN(n1279) );
  MUX2_X1 U248 ( .A(n1281), .B(n1282), .S(n1190), .Z(n1277) );
  NAND2_X2 U249 ( .A1(n1264), .A2(n1193), .ZN(n1282) );
  NAND2_X2 U250 ( .A1(n1283), .A2(n1193), .ZN(n1281) );
  NAND2_X2 U251 ( .A1(n1284), .A2(n1164), .ZN(n1275) );
  NAND2_X2 U252 ( .A1(n1285), .A2(n1286), .ZN(B[3]) );
  MUX2_X1 U253 ( .A(n1287), .B(n1288), .S(n1184), .Z(n1286) );
  NAND2_X2 U254 ( .A1(n1172), .A2(n1237), .ZN(n1288) );
  NAND2_X2 U255 ( .A1(n1171), .A2(n1289), .ZN(n1287) );
  MUX2_X1 U256 ( .A(n1290), .B(n1291), .S(n1184), .Z(n1285) );
  NAND2_X2 U257 ( .A1(n1241), .A2(n1164), .ZN(n1291) );
  NAND2_X2 U258 ( .A1(n1292), .A2(n1293), .ZN(n1241) );
  MUX2_X1 U259 ( .A(n1294), .B(n1295), .S(n1190), .Z(n1293) );
  NAND2_X2 U260 ( .A1(n1208), .A2(n1264), .ZN(n1295) );
  NAND2_X2 U261 ( .A1(n1209), .A2(n1283), .ZN(n1294) );
  MUX2_X1 U262 ( .A(n1296), .B(n1297), .S(n1190), .Z(n1292) );
  NAND2_X2 U263 ( .A1(n1268), .A2(n1193), .ZN(n1297) );
  NAND2_X2 U264 ( .A1(n1298), .A2(n1193), .ZN(n1296) );
  OAI21_X2 U265 ( .B1(n1299), .B2(n1300), .A(n1164), .ZN(n1290) );
  MUX2_X1 U266 ( .A(n1301), .B(n1302), .S(n1190), .Z(n1300) );
  AND2_X2 U267 ( .A1(n1303), .A2(n1197), .ZN(n1302) );
  AND2_X2 U268 ( .A1(n1304), .A2(n1197), .ZN(n1301) );
  MUX2_X1 U269 ( .A(n1305), .B(n1306), .S(n1190), .Z(n1299) );
  AND2_X2 U270 ( .A1(n1210), .A2(n1307), .ZN(n1306) );
  AND2_X2 U271 ( .A1(n1211), .A2(n1308), .ZN(n1305) );
  AND3_X2 U272 ( .A1(n1186), .A2(n1165), .A3(n1309), .ZN(B[31]) );
  AND3_X2 U273 ( .A1(n1186), .A2(n1165), .A3(n1310), .ZN(B[30]) );
  NAND2_X2 U274 ( .A1(n1311), .A2(n1312), .ZN(B[2]) );
  MUX2_X1 U275 ( .A(n1313), .B(n1314), .S(n1184), .Z(n1312) );
  NAND2_X2 U276 ( .A1(n1171), .A2(n1247), .ZN(n1314) );
  NAND2_X2 U277 ( .A1(n1171), .A2(n1315), .ZN(n1313) );
  MUX2_X1 U278 ( .A(n1316), .B(n1317), .S(n1184), .Z(n1311) );
  NAND2_X2 U279 ( .A1(n1251), .A2(n1164), .ZN(n1317) );
  NAND2_X2 U280 ( .A1(n1318), .A2(n1319), .ZN(n1251) );
  MUX2_X1 U281 ( .A(n1320), .B(n1321), .S(n1190), .Z(n1319) );
  NAND2_X2 U282 ( .A1(n1209), .A2(n1268), .ZN(n1321) );
  INV_X2 U283 ( .A(n1322), .ZN(n1268) );
  MUX2_X1 U284 ( .A(n1323), .B(n1324), .S(n1176), .Z(n1322) );
  NAND2_X2 U285 ( .A1(n1208), .A2(n1298), .ZN(n1320) );
  MUX2_X1 U286 ( .A(n1325), .B(n1326), .S(n1190), .Z(n1318) );
  NAND2_X2 U287 ( .A1(n1283), .A2(n1193), .ZN(n1326) );
  NAND2_X2 U288 ( .A1(n1307), .A2(n1193), .ZN(n1325) );
  OAI21_X2 U289 ( .B1(n1327), .B2(n1328), .A(n1164), .ZN(n1316) );
  MUX2_X1 U290 ( .A(n1329), .B(n1330), .S(n1189), .Z(n1328) );
  AND2_X2 U291 ( .A1(n1308), .A2(n1197), .ZN(n1330) );
  AND2_X2 U292 ( .A1(n1331), .A2(n1197), .ZN(n1329) );
  MUX2_X1 U293 ( .A(n1332), .B(n1333), .S(n1189), .Z(n1327) );
  AND2_X2 U294 ( .A1(n1209), .A2(n1303), .ZN(n1333) );
  AND2_X2 U295 ( .A1(n1210), .A2(n1304), .ZN(n1332) );
  AND3_X2 U296 ( .A1(n1186), .A2(n1165), .A3(n1216), .ZN(B[29]) );
  AND3_X2 U297 ( .A1(n1186), .A2(n1165), .A3(n1226), .ZN(B[28]) );
  MUX2_X1 U298 ( .A(n1334), .B(n1335), .S(n1184), .Z(B[27]) );
  AND2_X2 U299 ( .A1(n1309), .A2(n1165), .ZN(n1335) );
  NOR2_X2 U300 ( .A1(n1169), .A2(n1336), .ZN(n1334) );
  MUX2_X1 U301 ( .A(n1337), .B(n1338), .S(n1184), .Z(B[26]) );
  AND2_X2 U302 ( .A1(n1310), .A2(n1165), .ZN(n1338) );
  NOR2_X2 U303 ( .A1(n1168), .A2(n1339), .ZN(n1337) );
  MUX2_X1 U304 ( .A(n1340), .B(n1341), .S(n1184), .Z(B[25]) );
  AND2_X2 U305 ( .A1(n1216), .A2(n1165), .ZN(n1341) );
  NOR2_X2 U306 ( .A1(n1169), .A2(n1342), .ZN(n1340) );
  MUX2_X1 U307 ( .A(n1343), .B(n1344), .S(n1184), .Z(B[24]) );
  NOR2_X2 U308 ( .A1(n1168), .A2(n1345), .ZN(n1344) );
  INV_X2 U309 ( .A(n1226), .ZN(n1345) );
  NOR2_X2 U310 ( .A1(n1167), .A2(n1346), .ZN(n1343) );
  MUX2_X1 U311 ( .A(n1347), .B(n1348), .S(n1184), .Z(B[23]) );
  NOR2_X2 U312 ( .A1(n1167), .A2(n1336), .ZN(n1348) );
  INV_X2 U313 ( .A(n1236), .ZN(n1336) );
  AND2_X2 U314 ( .A1(n1237), .A2(n1165), .ZN(n1347) );
  MUX2_X1 U315 ( .A(n1349), .B(n1350), .S(n1184), .Z(B[22]) );
  NOR2_X2 U316 ( .A1(n1168), .A2(n1339), .ZN(n1350) );
  INV_X2 U317 ( .A(n1246), .ZN(n1339) );
  AND2_X2 U318 ( .A1(n1247), .A2(n1165), .ZN(n1349) );
  MUX2_X1 U319 ( .A(n1351), .B(n1352), .S(n1184), .Z(B[21]) );
  NOR2_X2 U320 ( .A1(n1167), .A2(n1342), .ZN(n1352) );
  INV_X2 U321 ( .A(n1217), .ZN(n1342) );
  NAND2_X2 U322 ( .A1(n1353), .A2(n1354), .ZN(n1217) );
  MUX2_X1 U323 ( .A(n1355), .B(n1356), .S(n1189), .Z(n1354) );
  NAND2_X2 U324 ( .A1(n1357), .A2(n1198), .ZN(n1356) );
  NAND2_X2 U325 ( .A1(n1358), .A2(n1198), .ZN(n1355) );
  MUX2_X1 U326 ( .A(n1359), .B(n1360), .S(n1189), .Z(n1353) );
  NAND2_X2 U327 ( .A1(n1361), .A2(n1193), .ZN(n1360) );
  NAND2_X2 U328 ( .A1(n1362), .A2(n1193), .ZN(n1359) );
  AND2_X2 U329 ( .A1(n1256), .A2(n1165), .ZN(n1351) );
  MUX2_X1 U330 ( .A(n1363), .B(n1364), .S(n1184), .Z(B[20]) );
  NOR2_X2 U331 ( .A1(n1168), .A2(n1346), .ZN(n1364) );
  INV_X2 U332 ( .A(n1227), .ZN(n1346) );
  NAND2_X2 U333 ( .A1(n1365), .A2(n1366), .ZN(n1227) );
  MUX2_X1 U334 ( .A(n1367), .B(n1368), .S(n1189), .Z(n1366) );
  NAND2_X2 U335 ( .A1(n1361), .A2(n1199), .ZN(n1368) );
  NAND2_X2 U336 ( .A1(n1362), .A2(n1200), .ZN(n1367) );
  MUX2_X1 U337 ( .A(n1369), .B(n1370), .S(n1189), .Z(n1365) );
  NAND2_X2 U338 ( .A1(n1358), .A2(n1193), .ZN(n1370) );
  NAND2_X2 U339 ( .A1(n1371), .A2(n1193), .ZN(n1369) );
  AND2_X2 U340 ( .A1(n1274), .A2(n1165), .ZN(n1363) );
  NAND2_X2 U341 ( .A1(n1372), .A2(n1373), .ZN(B[1]) );
  MUX2_X1 U342 ( .A(n1374), .B(n1375), .S(n1184), .Z(n1373) );
  NAND2_X2 U343 ( .A1(n1170), .A2(n1256), .ZN(n1375) );
  NAND2_X2 U344 ( .A1(n1170), .A2(n1376), .ZN(n1374) );
  MUX2_X1 U345 ( .A(n1377), .B(n1378), .S(n1183), .Z(n1372) );
  NAND2_X2 U346 ( .A1(n1269), .A2(n1164), .ZN(n1378) );
  NAND2_X2 U347 ( .A1(n1379), .A2(n1380), .ZN(n1269) );
  MUX2_X1 U348 ( .A(n1381), .B(n1382), .S(n1189), .Z(n1380) );
  NAND2_X2 U349 ( .A1(n1208), .A2(n1283), .ZN(n1382) );
  INV_X2 U350 ( .A(n1383), .ZN(n1283) );
  MUX2_X1 U351 ( .A(n1384), .B(n1385), .S(n1176), .Z(n1383) );
  NAND2_X2 U352 ( .A1(n1207), .A2(n1307), .ZN(n1381) );
  MUX2_X1 U353 ( .A(n1386), .B(n1387), .S(n1189), .Z(n1379) );
  NAND2_X2 U354 ( .A1(n1298), .A2(n1193), .ZN(n1387) );
  NAND2_X2 U355 ( .A1(n1303), .A2(n1194), .ZN(n1386) );
  OAI21_X2 U356 ( .B1(n1388), .B2(n1389), .A(n1164), .ZN(n1377) );
  MUX2_X1 U357 ( .A(n1390), .B(n1391), .S(n1189), .Z(n1389) );
  AND2_X2 U358 ( .A1(n1304), .A2(n1197), .ZN(n1391) );
  AND2_X2 U359 ( .A1(n1392), .A2(n1197), .ZN(n1390) );
  MUX2_X1 U360 ( .A(n1393), .B(n1394), .S(n1189), .Z(n1388) );
  AND2_X2 U361 ( .A1(n1208), .A2(n1308), .ZN(n1394) );
  AND2_X2 U362 ( .A1(n1210), .A2(n1331), .ZN(n1393) );
  MUX2_X1 U363 ( .A(n1395), .B(n1396), .S(n1183), .Z(B[19]) );
  AND2_X2 U364 ( .A1(n1237), .A2(n1165), .ZN(n1396) );
  NAND2_X2 U365 ( .A1(n1397), .A2(n1398), .ZN(n1237) );
  MUX2_X1 U366 ( .A(n1399), .B(n1400), .S(n1189), .Z(n1398) );
  NAND2_X2 U367 ( .A1(n1358), .A2(n1199), .ZN(n1400) );
  NAND2_X2 U368 ( .A1(n1371), .A2(n1201), .ZN(n1399) );
  MUX2_X1 U369 ( .A(n1401), .B(n1402), .S(n1189), .Z(n1397) );
  NAND2_X2 U370 ( .A1(n1362), .A2(n1194), .ZN(n1402) );
  NAND2_X2 U371 ( .A1(n1403), .A2(n1194), .ZN(n1401) );
  AND2_X2 U372 ( .A1(n1289), .A2(n1165), .ZN(n1395) );
  MUX2_X1 U373 ( .A(n1404), .B(n1405), .S(n1183), .Z(B[18]) );
  AND2_X2 U374 ( .A1(n1247), .A2(n1165), .ZN(n1405) );
  NAND2_X2 U375 ( .A1(n1406), .A2(n1407), .ZN(n1247) );
  MUX2_X1 U376 ( .A(n1408), .B(n1409), .S(n1189), .Z(n1407) );
  NAND2_X2 U377 ( .A1(n1362), .A2(n1198), .ZN(n1409) );
  INV_X2 U378 ( .A(n1410), .ZN(n1362) );
  NAND2_X2 U379 ( .A1(n1208), .A2(n1403), .ZN(n1408) );
  MUX2_X1 U380 ( .A(n1411), .B(n1412), .S(n1189), .Z(n1406) );
  NAND2_X2 U381 ( .A1(n1371), .A2(n1194), .ZN(n1412) );
  NAND2_X2 U382 ( .A1(n1413), .A2(n1194), .ZN(n1411) );
  AND2_X2 U383 ( .A1(n1315), .A2(n1165), .ZN(n1404) );
  MUX2_X1 U384 ( .A(n1414), .B(n1415), .S(n1183), .Z(B[17]) );
  AND2_X2 U385 ( .A1(n1256), .A2(n1165), .ZN(n1415) );
  NAND2_X2 U386 ( .A1(n1416), .A2(n1417), .ZN(n1256) );
  MUX2_X1 U387 ( .A(n1418), .B(n1419), .S(n1189), .Z(n1417) );
  NAND2_X2 U388 ( .A1(n1371), .A2(n1200), .ZN(n1419) );
  INV_X2 U389 ( .A(n1420), .ZN(n1371) );
  NAND2_X2 U390 ( .A1(n1207), .A2(n1413), .ZN(n1418) );
  MUX2_X1 U391 ( .A(n1421), .B(n1422), .S(n1189), .Z(n1416) );
  NAND2_X2 U392 ( .A1(n1403), .A2(n1194), .ZN(n1422) );
  NAND2_X2 U393 ( .A1(n1423), .A2(n1194), .ZN(n1421) );
  AND2_X2 U394 ( .A1(n1376), .A2(n1165), .ZN(n1414) );
  MUX2_X1 U395 ( .A(n1424), .B(n1425), .S(n1183), .Z(B[16]) );
  AND2_X2 U396 ( .A1(n1274), .A2(n1165), .ZN(n1425) );
  AND2_X2 U397 ( .A1(n1426), .A2(n1165), .ZN(n1424) );
  NAND2_X2 U398 ( .A1(n1427), .A2(n1428), .ZN(B[15]) );
  NAND3_X1 U399 ( .A1(n1186), .A2(n1165), .A3(n1429), .ZN(n1428) );
  MUX2_X1 U400 ( .A(n1430), .B(n1431), .S(n1169), .Z(n1427) );
  NAND2_X2 U401 ( .A1(n1309), .A2(n1186), .ZN(n1431) );
  NAND2_X2 U402 ( .A1(n1183), .A2(n1289), .ZN(n1430) );
  NAND2_X2 U403 ( .A1(n1432), .A2(n1433), .ZN(n1289) );
  MUX2_X1 U404 ( .A(n1434), .B(n1435), .S(n1189), .Z(n1433) );
  NAND2_X2 U405 ( .A1(n1207), .A2(n1413), .ZN(n1435) );
  NAND2_X2 U406 ( .A1(n1206), .A2(n1436), .ZN(n1434) );
  MUX2_X1 U407 ( .A(n1437), .B(n1438), .S(n1188), .Z(n1432) );
  NAND2_X2 U408 ( .A1(n1423), .A2(n1194), .ZN(n1438) );
  NAND2_X2 U409 ( .A1(n1439), .A2(n1194), .ZN(n1437) );
  NAND2_X2 U410 ( .A1(n1440), .A2(n1441), .ZN(B[14]) );
  NAND3_X1 U411 ( .A1(n1186), .A2(n1166), .A3(n1442), .ZN(n1441) );
  MUX2_X1 U412 ( .A(n1443), .B(n1444), .S(n1172), .Z(n1440) );
  NAND2_X2 U413 ( .A1(n1310), .A2(n1186), .ZN(n1444) );
  NAND2_X2 U414 ( .A1(n1183), .A2(n1315), .ZN(n1443) );
  NAND2_X2 U415 ( .A1(n1445), .A2(n1446), .ZN(n1315) );
  MUX2_X1 U416 ( .A(n1447), .B(n1448), .S(n1188), .Z(n1446) );
  NAND2_X2 U417 ( .A1(n1207), .A2(n1423), .ZN(n1448) );
  NAND2_X2 U418 ( .A1(n1206), .A2(n1439), .ZN(n1447) );
  MUX2_X1 U419 ( .A(n1449), .B(n1450), .S(n1188), .Z(n1445) );
  NAND2_X2 U420 ( .A1(n1436), .A2(n1194), .ZN(n1450) );
  NAND2_X2 U421 ( .A1(n1451), .A2(n1194), .ZN(n1449) );
  NAND2_X2 U422 ( .A1(n1452), .A2(n1453), .ZN(B[13]) );
  NAND3_X1 U423 ( .A1(n1186), .A2(n1166), .A3(n1220), .ZN(n1453) );
  NAND2_X2 U424 ( .A1(n1454), .A2(n1455), .ZN(n1220) );
  MUX2_X1 U425 ( .A(n1456), .B(n1457), .S(n1188), .Z(n1455) );
  NAND2_X2 U426 ( .A1(n1206), .A2(n1458), .ZN(n1457) );
  NAND2_X2 U427 ( .A1(n1206), .A2(n1459), .ZN(n1456) );
  MUX2_X1 U428 ( .A(n1460), .B(n1461), .S(n1188), .Z(n1454) );
  NAND2_X2 U429 ( .A1(n1462), .A2(n1194), .ZN(n1461) );
  NAND2_X2 U430 ( .A1(n1463), .A2(n1195), .ZN(n1460) );
  MUX2_X1 U431 ( .A(n1464), .B(n1465), .S(n1170), .Z(n1452) );
  NAND2_X2 U432 ( .A1(n1216), .A2(n1186), .ZN(n1465) );
  NAND2_X2 U433 ( .A1(n1466), .A2(n1467), .ZN(n1216) );
  NAND3_X1 U434 ( .A1(n1197), .A2(n1192), .A3(n1468), .ZN(n1467) );
  MUX2_X1 U435 ( .A(n1469), .B(n1470), .S(n1201), .Z(n1466) );
  NAND2_X2 U436 ( .A1(n1471), .A2(n1191), .ZN(n1470) );
  NAND2_X2 U437 ( .A1(n1187), .A2(n1472), .ZN(n1469) );
  NAND2_X2 U438 ( .A1(n1183), .A2(n1376), .ZN(n1464) );
  NAND2_X2 U439 ( .A1(n1473), .A2(n1474), .ZN(n1376) );
  MUX2_X1 U440 ( .A(n1475), .B(n1476), .S(n1188), .Z(n1474) );
  NAND2_X2 U441 ( .A1(n1205), .A2(n1436), .ZN(n1476) );
  NAND2_X2 U442 ( .A1(n1205), .A2(n1451), .ZN(n1475) );
  MUX2_X1 U443 ( .A(n1477), .B(n1478), .S(n1188), .Z(n1473) );
  NAND2_X2 U444 ( .A1(n1439), .A2(n1195), .ZN(n1478) );
  NAND2_X2 U445 ( .A1(n1479), .A2(n1195), .ZN(n1477) );
  NAND2_X2 U446 ( .A1(n1480), .A2(n1481), .ZN(B[12]) );
  NAND3_X1 U447 ( .A1(n1186), .A2(n1166), .A3(n1230), .ZN(n1481) );
  NAND2_X2 U448 ( .A1(n1482), .A2(n1483), .ZN(n1230) );
  MUX2_X1 U449 ( .A(n1484), .B(n1485), .S(n1188), .Z(n1483) );
  NAND2_X2 U450 ( .A1(n1205), .A2(n1462), .ZN(n1485) );
  NAND2_X2 U451 ( .A1(n1204), .A2(n1463), .ZN(n1484) );
  MUX2_X1 U452 ( .A(n1486), .B(n1487), .S(n1188), .Z(n1482) );
  NAND2_X2 U453 ( .A1(n1459), .A2(n1195), .ZN(n1487) );
  NAND2_X2 U454 ( .A1(n1263), .A2(n1195), .ZN(n1486) );
  MUX2_X1 U455 ( .A(n1488), .B(n1489), .S(n1171), .Z(n1480) );
  NAND2_X2 U456 ( .A1(n1226), .A2(n1186), .ZN(n1489) );
  NAND2_X2 U457 ( .A1(n1490), .A2(n1491), .ZN(n1226) );
  MUX2_X1 U458 ( .A(n1492), .B(n1493), .S(n1188), .Z(n1491) );
  NAND2_X2 U459 ( .A1(n1472), .A2(n1199), .ZN(n1493) );
  NAND2_X2 U460 ( .A1(n1468), .A2(n1200), .ZN(n1492) );
  MUX2_X1 U461 ( .A(n1494), .B(n1495), .S(n1188), .Z(n1490) );
  NAND2_X2 U462 ( .A1(n1471), .A2(n1195), .ZN(n1495) );
  NAND2_X2 U463 ( .A1(n1357), .A2(n1195), .ZN(n1494) );
  NAND2_X2 U464 ( .A1(n1183), .A2(n1426), .ZN(n1488) );
  NAND2_X2 U465 ( .A1(n1496), .A2(n1497), .ZN(B[11]) );
  MUX2_X1 U466 ( .A(n1498), .B(n1499), .S(n1183), .Z(n1497) );
  NAND2_X2 U467 ( .A1(n1309), .A2(n1167), .ZN(n1499) );
  INV_X2 U468 ( .A(n1500), .ZN(n1309) );
  NAND3_X1 U469 ( .A1(n1197), .A2(n1192), .A3(n1472), .ZN(n1500) );
  NAND2_X2 U470 ( .A1(n1170), .A2(n1236), .ZN(n1498) );
  NAND2_X2 U471 ( .A1(n1501), .A2(n1502), .ZN(n1236) );
  MUX2_X1 U472 ( .A(n1503), .B(n1504), .S(n1188), .Z(n1502) );
  NAND2_X2 U473 ( .A1(n1205), .A2(n1471), .ZN(n1504) );
  NAND2_X2 U474 ( .A1(n1357), .A2(n1200), .ZN(n1503) );
  MUX2_X1 U475 ( .A(n1505), .B(n1506), .S(n1188), .Z(n1501) );
  NAND2_X2 U476 ( .A1(n1468), .A2(n1195), .ZN(n1506) );
  NAND2_X2 U477 ( .A1(n1361), .A2(n1195), .ZN(n1505) );
  MUX2_X1 U478 ( .A(n1507), .B(n1508), .S(n1183), .Z(n1496) );
  NAND2_X2 U479 ( .A1(n1429), .A2(n1163), .ZN(n1508) );
  NAND2_X2 U480 ( .A1(n1509), .A2(n1510), .ZN(n1429) );
  MUX2_X1 U481 ( .A(n1511), .B(n1512), .S(n1188), .Z(n1510) );
  NAND2_X2 U482 ( .A1(n1204), .A2(n1451), .ZN(n1512) );
  NAND2_X2 U483 ( .A1(n1202), .A2(n1458), .ZN(n1511) );
  MUX2_X1 U484 ( .A(n1513), .B(n1514), .S(n1188), .Z(n1509) );
  NAND2_X2 U485 ( .A1(n1479), .A2(n1196), .ZN(n1514) );
  NAND2_X2 U486 ( .A1(n1462), .A2(n1195), .ZN(n1513) );
  NAND2_X2 U487 ( .A1(n1240), .A2(n1163), .ZN(n1507) );
  NAND2_X2 U488 ( .A1(n1515), .A2(n1516), .ZN(n1240) );
  MUX2_X1 U489 ( .A(n1517), .B(n1518), .S(n1187), .Z(n1516) );
  NAND2_X2 U490 ( .A1(n1204), .A2(n1459), .ZN(n1518) );
  NAND2_X2 U491 ( .A1(n1202), .A2(n1263), .ZN(n1517) );
  MUX2_X1 U492 ( .A(n1519), .B(n1520), .S(n1188), .Z(n1515) );
  NAND2_X2 U493 ( .A1(n1463), .A2(n1196), .ZN(n1520) );
  NAND2_X2 U494 ( .A1(n1267), .A2(n1195), .ZN(n1519) );
  NAND2_X2 U495 ( .A1(n1521), .A2(n1522), .ZN(B[10]) );
  MUX2_X1 U496 ( .A(n1523), .B(n1524), .S(n1183), .Z(n1522) );
  NAND2_X2 U497 ( .A1(n1170), .A2(n1310), .ZN(n1524) );
  MUX2_X1 U498 ( .A(n1525), .B(n1526), .S(n1202), .Z(n1310) );
  INV_X2 U499 ( .A(n1527), .ZN(n1526) );
  NAND2_X2 U500 ( .A1(n1472), .A2(n1191), .ZN(n1527) );
  INV_X2 U501 ( .A(n1528), .ZN(n1472) );
  INV_X2 U502 ( .A(n1529), .ZN(n1525) );
  NAND2_X2 U503 ( .A1(n1471), .A2(n1191), .ZN(n1529) );
  INV_X2 U504 ( .A(n1530), .ZN(n1471) );
  NAND2_X2 U505 ( .A1(n1169), .A2(n1246), .ZN(n1523) );
  NAND2_X2 U506 ( .A1(n1531), .A2(n1532), .ZN(n1246) );
  MUX2_X1 U507 ( .A(n1533), .B(n1534), .S(n1187), .Z(n1532) );
  NAND2_X2 U508 ( .A1(n1468), .A2(n1198), .ZN(n1534) );
  INV_X2 U509 ( .A(n1535), .ZN(n1468) );
  NAND2_X2 U510 ( .A1(n1361), .A2(n1199), .ZN(n1533) );
  INV_X2 U511 ( .A(n1536), .ZN(n1361) );
  MUX2_X1 U512 ( .A(n1537), .B(n1538), .S(n1187), .Z(n1531) );
  NAND2_X2 U513 ( .A1(n1357), .A2(n1196), .ZN(n1538) );
  INV_X2 U514 ( .A(n1539), .ZN(n1357) );
  NAND2_X2 U515 ( .A1(n1358), .A2(n1196), .ZN(n1537) );
  INV_X2 U516 ( .A(n1540), .ZN(n1358) );
  MUX2_X1 U517 ( .A(n1541), .B(n1542), .S(n1183), .Z(n1521) );
  NAND2_X2 U518 ( .A1(n1442), .A2(n1163), .ZN(n1542) );
  NAND2_X2 U519 ( .A1(n1543), .A2(n1544), .ZN(n1442) );
  MUX2_X1 U520 ( .A(n1545), .B(n1546), .S(n1187), .Z(n1544) );
  NAND2_X2 U521 ( .A1(n1204), .A2(n1479), .ZN(n1546) );
  NAND2_X2 U522 ( .A1(n1202), .A2(n1462), .ZN(n1545) );
  INV_X2 U523 ( .A(n1547), .ZN(n1462) );
  MUX2_X1 U524 ( .A(n1548), .B(n1549), .S(n1176), .Z(n1547) );
  MUX2_X1 U525 ( .A(n1550), .B(n1551), .S(n1187), .Z(n1543) );
  NAND2_X2 U526 ( .A1(n1458), .A2(n1196), .ZN(n1551) );
  NAND2_X2 U527 ( .A1(n1459), .A2(n1196), .ZN(n1550) );
  INV_X2 U528 ( .A(n1552), .ZN(n1459) );
  MUX2_X1 U529 ( .A(n1553), .B(n1554), .S(n1176), .Z(n1552) );
  NAND2_X2 U530 ( .A1(n1250), .A2(n1163), .ZN(n1541) );
  NAND2_X2 U531 ( .A1(n1555), .A2(n1556), .ZN(n1250) );
  MUX2_X1 U532 ( .A(n1557), .B(n1558), .S(n1187), .Z(n1556) );
  NAND2_X2 U533 ( .A1(n1203), .A2(n1463), .ZN(n1558) );
  INV_X2 U534 ( .A(n1559), .ZN(n1463) );
  MUX2_X1 U535 ( .A(n1560), .B(n1561), .S(n1176), .Z(n1559) );
  NAND2_X2 U536 ( .A1(n1202), .A2(n1267), .ZN(n1557) );
  INV_X2 U537 ( .A(n1562), .ZN(n1267) );
  MUX2_X1 U538 ( .A(n1563), .B(n1564), .S(n1176), .Z(n1562) );
  MUX2_X1 U539 ( .A(n1565), .B(n1566), .S(n1187), .Z(n1555) );
  NAND2_X2 U540 ( .A1(n1263), .A2(n1196), .ZN(n1566) );
  INV_X2 U541 ( .A(n1567), .ZN(n1263) );
  MUX2_X1 U542 ( .A(n1568), .B(n1569), .S(n1176), .Z(n1567) );
  NAND2_X2 U543 ( .A1(n1264), .A2(n1196), .ZN(n1565) );
  INV_X2 U544 ( .A(n1570), .ZN(n1264) );
  MUX2_X1 U545 ( .A(n1571), .B(n1572), .S(n1176), .Z(n1570) );
  NAND2_X2 U546 ( .A1(n1573), .A2(n1574), .ZN(B[0]) );
  MUX2_X1 U547 ( .A(n1575), .B(n1576), .S(n1183), .Z(n1574) );
  NAND2_X2 U548 ( .A1(n1169), .A2(n1274), .ZN(n1576) );
  NAND2_X2 U549 ( .A1(n1577), .A2(n1578), .ZN(n1274) );
  MUX2_X1 U550 ( .A(n1579), .B(n1580), .S(n1187), .Z(n1578) );
  NAND2_X2 U551 ( .A1(n1203), .A2(n1403), .ZN(n1580) );
  INV_X2 U552 ( .A(n1581), .ZN(n1403) );
  MUX2_X1 U553 ( .A(n1549), .B(n1582), .S(n1176), .Z(n1581) );
  NAND2_X2 U554 ( .A1(n1201), .A2(n1423), .ZN(n1579) );
  INV_X2 U555 ( .A(n1583), .ZN(n1423) );
  MUX2_X1 U556 ( .A(n1561), .B(n1584), .S(n1176), .Z(n1583) );
  MUX2_X1 U557 ( .A(n1585), .B(n1586), .S(n1187), .Z(n1577) );
  NAND2_X2 U558 ( .A1(n1413), .A2(n1196), .ZN(n1586) );
  INV_X2 U559 ( .A(n1587), .ZN(n1413) );
  MUX2_X1 U560 ( .A(n1554), .B(n1588), .S(n1176), .Z(n1587) );
  NAND2_X2 U561 ( .A1(n1436), .A2(n1196), .ZN(n1585) );
  INV_X2 U562 ( .A(n1589), .ZN(n1436) );
  MUX2_X1 U563 ( .A(n1569), .B(n1590), .S(n1176), .Z(n1589) );
  NAND2_X2 U564 ( .A1(n1171), .A2(n1426), .ZN(n1575) );
  NAND2_X2 U565 ( .A1(n1591), .A2(n1592), .ZN(n1426) );
  MUX2_X1 U566 ( .A(n1593), .B(n1594), .S(n1187), .Z(n1592) );
  NAND2_X2 U567 ( .A1(n1203), .A2(n1439), .ZN(n1594) );
  INV_X2 U568 ( .A(n1595), .ZN(n1439) );
  MUX2_X1 U569 ( .A(n1564), .B(n1596), .S(n1177), .Z(n1595) );
  NAND2_X2 U570 ( .A1(n1201), .A2(n1479), .ZN(n1593) );
  INV_X2 U571 ( .A(n1597), .ZN(n1479) );
  MUX2_X1 U572 ( .A(n1324), .B(n1598), .S(n1177), .Z(n1597) );
  MUX2_X1 U573 ( .A(n1599), .B(n1600), .S(n1187), .Z(n1591) );
  NAND2_X2 U574 ( .A1(n1451), .A2(n1197), .ZN(n1600) );
  INV_X2 U575 ( .A(n1601), .ZN(n1451) );
  MUX2_X1 U576 ( .A(n1572), .B(n1602), .S(n1177), .Z(n1601) );
  NAND2_X2 U577 ( .A1(n1458), .A2(n1196), .ZN(n1599) );
  INV_X2 U578 ( .A(n1603), .ZN(n1458) );
  MUX2_X1 U579 ( .A(n1385), .B(n1604), .S(n1177), .Z(n1603) );
  MUX2_X1 U580 ( .A(n1605), .B(n1606), .S(n1184), .Z(n1573) );
  NAND2_X2 U581 ( .A1(n1284), .A2(n1163), .ZN(n1606) );
  NAND2_X2 U582 ( .A1(n1607), .A2(n1608), .ZN(n1284) );
  MUX2_X1 U583 ( .A(n1609), .B(n1610), .S(n1187), .Z(n1608) );
  NAND2_X2 U584 ( .A1(n1203), .A2(n1298), .ZN(n1610) );
  INV_X2 U585 ( .A(n1611), .ZN(n1298) );
  MUX2_X1 U586 ( .A(n1612), .B(n1548), .S(n1177), .Z(n1611) );
  NAND2_X2 U587 ( .A1(n1201), .A2(n1303), .ZN(n1609) );
  INV_X2 U588 ( .A(n1613), .ZN(n1303) );
  MUX2_X1 U589 ( .A(n1614), .B(n1560), .S(n1177), .Z(n1613) );
  MUX2_X1 U590 ( .A(n1615), .B(n1616), .S(n1187), .Z(n1607) );
  NAND2_X2 U591 ( .A1(n1307), .A2(n1197), .ZN(n1616) );
  INV_X2 U592 ( .A(n1617), .ZN(n1307) );
  MUX2_X1 U593 ( .A(n1618), .B(n1553), .S(n1177), .Z(n1617) );
  NAND2_X2 U594 ( .A1(n1308), .A2(n1196), .ZN(n1615) );
  INV_X2 U595 ( .A(n1619), .ZN(n1308) );
  MUX2_X1 U596 ( .A(n1620), .B(n1568), .S(n1177), .Z(n1619) );
  OAI21_X2 U597 ( .B1(n1621), .B2(n1622), .A(n1164), .ZN(n1605) );
  MUX2_X1 U598 ( .A(n1623), .B(n1624), .S(n1187), .Z(n1622) );
  AND2_X2 U599 ( .A1(n1331), .A2(n1197), .ZN(n1624) );
  INV_X2 U600 ( .A(n1625), .ZN(n1331) );
  MUX2_X1 U601 ( .A(n1626), .B(n1571), .S(n1177), .Z(n1625) );
  AND2_X2 U602 ( .A1(n1627), .A2(n1197), .ZN(n1623) );
  MUX2_X1 U603 ( .A(A[0]), .B(A[8]), .S(n1177), .Z(n1627) );
  MUX2_X1 U604 ( .A(n1628), .B(n1629), .S(n1188), .Z(n1621) );
  AND2_X2 U605 ( .A1(n1211), .A2(n1304), .ZN(n1629) );
  INV_X2 U606 ( .A(n1630), .ZN(n1304) );
  MUX2_X1 U607 ( .A(n1631), .B(n1563), .S(n1177), .Z(n1630) );
  AND2_X2 U608 ( .A1(n1210), .A2(n1392), .ZN(n1628) );
  INV_X2 U609 ( .A(n1632), .ZN(n1392) );
  MUX2_X1 U610 ( .A(n1633), .B(n1323), .S(n1177), .Z(n1632) );
endmodule


module up_island_DW01_add_3 ( A, B, SUM, CI, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n107, n108, n109, n110, n111, n112,
         n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n360, n362, n364, n366, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414;

  XOR2_X2 U2 ( .A(B[63]), .B(A[63]), .Z(n1) );
  FA_X1 U3 ( .A(B[62]), .B(A[62]), .CI(n59), .CO(n58), .S(SUM[62]) );
  FA_X1 U4 ( .A(B[61]), .B(A[61]), .CI(n60), .CO(n59), .S(SUM[61]) );
  FA_X1 U5 ( .A(B[60]), .B(A[60]), .CI(n61), .CO(n60), .S(SUM[60]) );
  FA_X1 U6 ( .A(B[59]), .B(A[59]), .CI(n62), .CO(n61), .S(SUM[59]) );
  FA_X1 U7 ( .A(B[58]), .B(A[58]), .CI(n63), .CO(n62), .S(SUM[58]) );
  FA_X1 U8 ( .A(B[57]), .B(A[57]), .CI(n64), .CO(n63), .S(SUM[57]) );
  FA_X1 U9 ( .A(B[56]), .B(A[56]), .CI(n358), .CO(n64), .S(SUM[56]) );
  NAND2_X4 U15 ( .A1(n66), .A2(n69), .ZN(n2) );
  NOR2_X4 U17 ( .A1(B[55]), .A2(A[55]), .ZN(n68) );
  NAND2_X4 U18 ( .A1(B[55]), .A2(A[55]), .ZN(n69) );
  NAND2_X4 U21 ( .A1(n360), .A2(n72), .ZN(n3) );
  NOR2_X4 U23 ( .A1(B[54]), .A2(A[54]), .ZN(n71) );
  NAND2_X4 U24 ( .A1(B[54]), .A2(A[54]), .ZN(n72) );
  XNOR2_X2 U25 ( .A(n78), .B(n4), .ZN(SUM[53]) );
  AOI21_X4 U26 ( .B1(n78), .B2(n74), .A(n75), .ZN(n73) );
  NAND2_X4 U29 ( .A1(n74), .A2(n77), .ZN(n4) );
  NOR2_X4 U31 ( .A1(B[53]), .A2(A[53]), .ZN(n76) );
  NAND2_X4 U32 ( .A1(B[53]), .A2(A[53]), .ZN(n77) );
  XOR2_X2 U33 ( .A(n81), .B(n5), .Z(SUM[52]) );
  OAI21_X4 U34 ( .B1(n81), .B2(n79), .A(n80), .ZN(n78) );
  NAND2_X4 U35 ( .A1(n362), .A2(n80), .ZN(n5) );
  NOR2_X4 U37 ( .A1(B[52]), .A2(A[52]), .ZN(n79) );
  NAND2_X4 U38 ( .A1(B[52]), .A2(A[52]), .ZN(n80) );
  AOI21_X4 U40 ( .B1(n86), .B2(n82), .A(n83), .ZN(n81) );
  NAND2_X4 U43 ( .A1(n82), .A2(n85), .ZN(n6) );
  NOR2_X4 U45 ( .A1(B[51]), .A2(A[51]), .ZN(n84) );
  NAND2_X4 U46 ( .A1(B[51]), .A2(A[51]), .ZN(n85) );
  XOR2_X2 U47 ( .A(n89), .B(n7), .Z(SUM[50]) );
  NAND2_X4 U49 ( .A1(n364), .A2(n88), .ZN(n7) );
  NOR2_X4 U51 ( .A1(B[50]), .A2(A[50]), .ZN(n87) );
  NAND2_X4 U52 ( .A1(B[50]), .A2(A[50]), .ZN(n88) );
  AOI21_X4 U54 ( .B1(n94), .B2(n90), .A(n91), .ZN(n89) );
  NAND2_X4 U57 ( .A1(n90), .A2(n93), .ZN(n8) );
  NOR2_X4 U59 ( .A1(B[49]), .A2(A[49]), .ZN(n92) );
  NAND2_X4 U60 ( .A1(B[49]), .A2(A[49]), .ZN(n93) );
  XOR2_X2 U61 ( .A(n97), .B(n9), .Z(SUM[48]) );
  NAND2_X4 U63 ( .A1(n366), .A2(n96), .ZN(n9) );
  NOR2_X4 U65 ( .A1(B[48]), .A2(A[48]), .ZN(n95) );
  NAND2_X4 U66 ( .A1(B[48]), .A2(A[48]), .ZN(n96) );
  XNOR2_X2 U67 ( .A(n102), .B(n10), .ZN(SUM[47]) );
  AOI21_X4 U68 ( .B1(n102), .B2(n98), .A(n99), .ZN(n97) );
  NAND2_X4 U71 ( .A1(n98), .A2(n101), .ZN(n10) );
  NOR2_X4 U73 ( .A1(B[47]), .A2(A[47]), .ZN(n100) );
  NAND2_X4 U74 ( .A1(B[47]), .A2(A[47]), .ZN(n101) );
  NAND2_X4 U77 ( .A1(n368), .A2(n104), .ZN(n11) );
  NOR2_X4 U79 ( .A1(B[46]), .A2(A[46]), .ZN(n103) );
  NAND2_X4 U80 ( .A1(B[46]), .A2(A[46]), .ZN(n104) );
  XNOR2_X2 U81 ( .A(n110), .B(n12), .ZN(SUM[45]) );
  AOI21_X4 U82 ( .B1(n110), .B2(n369), .A(n107), .ZN(n105) );
  NAND2_X4 U85 ( .A1(n369), .A2(n109), .ZN(n12) );
  NOR2_X4 U87 ( .A1(B[45]), .A2(A[45]), .ZN(n108) );
  NAND2_X4 U88 ( .A1(B[45]), .A2(A[45]), .ZN(n109) );
  XOR2_X2 U89 ( .A(n113), .B(n13), .Z(SUM[44]) );
  OAI21_X4 U90 ( .B1(n113), .B2(n111), .A(n112), .ZN(n110) );
  NAND2_X4 U91 ( .A1(n370), .A2(n112), .ZN(n13) );
  NOR2_X4 U93 ( .A1(B[44]), .A2(A[44]), .ZN(n111) );
  NAND2_X4 U94 ( .A1(B[44]), .A2(A[44]), .ZN(n112) );
  AOI21_X4 U96 ( .B1(n118), .B2(n371), .A(n115), .ZN(n113) );
  NAND2_X4 U99 ( .A1(n371), .A2(n117), .ZN(n14) );
  NOR2_X4 U101 ( .A1(B[43]), .A2(A[43]), .ZN(n116) );
  NAND2_X4 U102 ( .A1(B[43]), .A2(A[43]), .ZN(n117) );
  NAND2_X4 U105 ( .A1(n372), .A2(n120), .ZN(n15) );
  NOR2_X4 U107 ( .A1(B[42]), .A2(A[42]), .ZN(n119) );
  NAND2_X4 U108 ( .A1(B[42]), .A2(A[42]), .ZN(n120) );
  XNOR2_X2 U109 ( .A(n126), .B(n16), .ZN(SUM[41]) );
  AOI21_X4 U110 ( .B1(n185), .B2(n122), .A(n123), .ZN(n121) );
  NOR2_X4 U111 ( .A1(n127), .A2(n124), .ZN(n122) );
  NAND2_X4 U113 ( .A1(n373), .A2(n125), .ZN(n16) );
  NOR2_X4 U115 ( .A1(B[41]), .A2(A[41]), .ZN(n124) );
  NAND2_X4 U116 ( .A1(B[41]), .A2(A[41]), .ZN(n125) );
  XNOR2_X2 U117 ( .A(n133), .B(n17), .ZN(SUM[40]) );
  NAND2_X4 U119 ( .A1(n136), .A2(n374), .ZN(n127) );
  AOI21_X4 U120 ( .B1(n137), .B2(n374), .A(n130), .ZN(n128) );
  NAND2_X4 U123 ( .A1(n374), .A2(n132), .ZN(n17) );
  NOR2_X4 U125 ( .A1(B[40]), .A2(A[40]), .ZN(n131) );
  NAND2_X4 U126 ( .A1(B[40]), .A2(A[40]), .ZN(n132) );
  XOR2_X2 U127 ( .A(n144), .B(n18), .Z(SUM[39]) );
  OAI21_X4 U128 ( .B1(n184), .B2(n134), .A(n135), .ZN(n133) );
  NOR2_X4 U131 ( .A1(n163), .A2(n138), .ZN(n136) );
  OAI21_X4 U132 ( .B1(n164), .B2(n138), .A(n139), .ZN(n137) );
  NAND2_X4 U133 ( .A1(n152), .A2(n140), .ZN(n138) );
  AOI21_X4 U134 ( .B1(n140), .B2(n153), .A(n141), .ZN(n139) );
  NOR2_X4 U135 ( .A1(n147), .A2(n142), .ZN(n140) );
  OAI21_X4 U136 ( .B1(n142), .B2(n148), .A(n143), .ZN(n141) );
  NAND2_X4 U137 ( .A1(n375), .A2(n143), .ZN(n18) );
  NOR2_X4 U139 ( .A1(B[39]), .A2(A[39]), .ZN(n142) );
  NAND2_X4 U140 ( .A1(B[39]), .A2(A[39]), .ZN(n143) );
  XNOR2_X2 U141 ( .A(n149), .B(n19), .ZN(SUM[38]) );
  AOI21_X4 U142 ( .B1(n149), .B2(n376), .A(n146), .ZN(n144) );
  NAND2_X4 U145 ( .A1(n376), .A2(n148), .ZN(n19) );
  NOR2_X4 U147 ( .A1(B[38]), .A2(A[38]), .ZN(n147) );
  NAND2_X4 U148 ( .A1(B[38]), .A2(A[38]), .ZN(n148) );
  XOR2_X2 U149 ( .A(n156), .B(n20), .Z(SUM[37]) );
  OAI21_X4 U150 ( .B1(n161), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X4 U153 ( .A1(n159), .A2(n154), .ZN(n152) );
  OAI21_X4 U154 ( .B1(n154), .B2(n160), .A(n155), .ZN(n153) );
  NAND2_X4 U155 ( .A1(n377), .A2(n155), .ZN(n20) );
  NOR2_X4 U157 ( .A1(B[37]), .A2(A[37]), .ZN(n154) );
  NAND2_X4 U158 ( .A1(B[37]), .A2(A[37]), .ZN(n155) );
  XOR2_X2 U159 ( .A(n161), .B(n21), .Z(SUM[36]) );
  AOI21_X4 U160 ( .B1(n162), .B2(n378), .A(n158), .ZN(n156) );
  NAND2_X4 U163 ( .A1(n378), .A2(n160), .ZN(n21) );
  NOR2_X4 U165 ( .A1(B[36]), .A2(A[36]), .ZN(n159) );
  NAND2_X4 U166 ( .A1(B[36]), .A2(A[36]), .ZN(n160) );
  XOR2_X2 U167 ( .A(n169), .B(n22), .Z(SUM[35]) );
  OAI21_X4 U169 ( .B1(n184), .B2(n163), .A(n164), .ZN(n162) );
  NAND2_X4 U170 ( .A1(n177), .A2(n165), .ZN(n163) );
  AOI21_X4 U171 ( .B1(n165), .B2(n178), .A(n166), .ZN(n164) );
  NOR2_X4 U172 ( .A1(n172), .A2(n167), .ZN(n165) );
  NAND2_X4 U174 ( .A1(n379), .A2(n168), .ZN(n22) );
  NOR2_X4 U176 ( .A1(B[35]), .A2(A[35]), .ZN(n167) );
  NAND2_X4 U177 ( .A1(B[35]), .A2(A[35]), .ZN(n168) );
  XNOR2_X2 U178 ( .A(n174), .B(n23), .ZN(SUM[34]) );
  AOI21_X4 U179 ( .B1(n174), .B2(n380), .A(n171), .ZN(n169) );
  NAND2_X4 U182 ( .A1(n380), .A2(n173), .ZN(n23) );
  NOR2_X4 U184 ( .A1(B[34]), .A2(A[34]), .ZN(n172) );
  NAND2_X4 U185 ( .A1(B[34]), .A2(A[34]), .ZN(n173) );
  XNOR2_X2 U186 ( .A(n181), .B(n24), .ZN(SUM[33]) );
  OAI21_X4 U187 ( .B1(n184), .B2(n175), .A(n176), .ZN(n174) );
  NOR2_X4 U190 ( .A1(n182), .A2(n179), .ZN(n177) );
  NAND2_X4 U192 ( .A1(n381), .A2(n180), .ZN(n24) );
  NOR2_X4 U194 ( .A1(B[33]), .A2(A[33]), .ZN(n179) );
  NAND2_X4 U195 ( .A1(B[33]), .A2(A[33]), .ZN(n180) );
  XOR2_X2 U196 ( .A(n184), .B(n25), .Z(SUM[32]) );
  OAI21_X4 U197 ( .B1(n184), .B2(n182), .A(n183), .ZN(n181) );
  NAND2_X4 U198 ( .A1(n382), .A2(n183), .ZN(n25) );
  NOR2_X4 U200 ( .A1(B[32]), .A2(A[32]), .ZN(n182) );
  NAND2_X4 U201 ( .A1(B[32]), .A2(A[32]), .ZN(n183) );
  XNOR2_X2 U202 ( .A(n196), .B(n26), .ZN(SUM[31]) );
  OAI21_X4 U204 ( .B1(n273), .B2(n186), .A(n187), .ZN(n185) );
  NAND2_X4 U205 ( .A1(n230), .A2(n188), .ZN(n186) );
  AOI21_X4 U206 ( .B1(n231), .B2(n188), .A(n189), .ZN(n187) );
  NOR2_X4 U207 ( .A1(n211), .A2(n190), .ZN(n188) );
  OAI21_X4 U208 ( .B1(n212), .B2(n190), .A(n191), .ZN(n189) );
  NAND2_X4 U209 ( .A1(n200), .A2(n192), .ZN(n190) );
  AOI21_X4 U210 ( .B1(n192), .B2(n201), .A(n193), .ZN(n191) );
  NOR2_X4 U211 ( .A1(n197), .A2(n194), .ZN(n192) );
  OAI21_X4 U212 ( .B1(n194), .B2(n198), .A(n195), .ZN(n193) );
  NAND2_X4 U213 ( .A1(n383), .A2(n195), .ZN(n26) );
  NOR2_X4 U215 ( .A1(B[31]), .A2(A[31]), .ZN(n194) );
  NAND2_X4 U216 ( .A1(B[31]), .A2(A[31]), .ZN(n195) );
  XOR2_X2 U217 ( .A(n199), .B(n27), .Z(SUM[30]) );
  OAI21_X4 U218 ( .B1(n199), .B2(n197), .A(n198), .ZN(n196) );
  NAND2_X4 U219 ( .A1(n384), .A2(n198), .ZN(n27) );
  NOR2_X4 U221 ( .A1(B[30]), .A2(A[30]), .ZN(n197) );
  NAND2_X4 U222 ( .A1(B[30]), .A2(A[30]), .ZN(n198) );
  XNOR2_X2 U223 ( .A(n204), .B(n28), .ZN(SUM[29]) );
  AOI21_X4 U224 ( .B1(n207), .B2(n200), .A(n201), .ZN(n199) );
  NOR2_X4 U225 ( .A1(n205), .A2(n202), .ZN(n200) );
  OAI21_X4 U226 ( .B1(n202), .B2(n206), .A(n203), .ZN(n201) );
  NAND2_X4 U227 ( .A1(n385), .A2(n203), .ZN(n28) );
  NOR2_X4 U229 ( .A1(B[29]), .A2(A[29]), .ZN(n202) );
  NAND2_X4 U230 ( .A1(B[29]), .A2(A[29]), .ZN(n203) );
  XNOR2_X2 U231 ( .A(n207), .B(n29), .ZN(SUM[28]) );
  OAI21_X4 U232 ( .B1(n208), .B2(n205), .A(n206), .ZN(n204) );
  NAND2_X4 U233 ( .A1(n386), .A2(n206), .ZN(n29) );
  NOR2_X4 U235 ( .A1(B[28]), .A2(A[28]), .ZN(n205) );
  NAND2_X4 U236 ( .A1(B[28]), .A2(A[28]), .ZN(n206) );
  XNOR2_X2 U237 ( .A(n217), .B(n30), .ZN(SUM[27]) );
  AOI21_X4 U239 ( .B1(n228), .B2(n209), .A(n210), .ZN(n208) );
  NAND2_X4 U242 ( .A1(n221), .A2(n213), .ZN(n211) );
  AOI21_X4 U243 ( .B1(n213), .B2(n222), .A(n214), .ZN(n212) );
  NOR2_X4 U244 ( .A1(n218), .A2(n215), .ZN(n213) );
  OAI21_X4 U245 ( .B1(n215), .B2(n219), .A(n216), .ZN(n214) );
  NAND2_X4 U246 ( .A1(n387), .A2(n216), .ZN(n30) );
  NOR2_X4 U248 ( .A1(B[27]), .A2(A[27]), .ZN(n215) );
  NAND2_X4 U249 ( .A1(B[27]), .A2(A[27]), .ZN(n216) );
  XOR2_X2 U250 ( .A(n220), .B(n31), .Z(SUM[26]) );
  OAI21_X4 U251 ( .B1(n220), .B2(n218), .A(n219), .ZN(n217) );
  NAND2_X4 U252 ( .A1(n388), .A2(n219), .ZN(n31) );
  NOR2_X4 U254 ( .A1(B[26]), .A2(A[26]), .ZN(n218) );
  NAND2_X4 U255 ( .A1(B[26]), .A2(A[26]), .ZN(n219) );
  XNOR2_X2 U256 ( .A(n225), .B(n32), .ZN(SUM[25]) );
  AOI21_X4 U257 ( .B1(n228), .B2(n221), .A(n222), .ZN(n220) );
  NOR2_X4 U258 ( .A1(n226), .A2(n223), .ZN(n221) );
  OAI21_X4 U259 ( .B1(n223), .B2(n227), .A(n224), .ZN(n222) );
  NAND2_X4 U260 ( .A1(n389), .A2(n224), .ZN(n32) );
  NOR2_X4 U262 ( .A1(B[25]), .A2(A[25]), .ZN(n223) );
  NAND2_X4 U263 ( .A1(B[25]), .A2(A[25]), .ZN(n224) );
  XNOR2_X2 U264 ( .A(n228), .B(n33), .ZN(SUM[24]) );
  OAI21_X4 U265 ( .B1(n229), .B2(n226), .A(n227), .ZN(n225) );
  NAND2_X4 U266 ( .A1(n390), .A2(n227), .ZN(n33) );
  NOR2_X4 U268 ( .A1(B[24]), .A2(A[24]), .ZN(n226) );
  NAND2_X4 U269 ( .A1(B[24]), .A2(A[24]), .ZN(n227) );
  XNOR2_X2 U270 ( .A(n238), .B(n34), .ZN(SUM[23]) );
  AOI21_X4 U272 ( .B1(n272), .B2(n230), .A(n231), .ZN(n229) );
  NOR2_X4 U273 ( .A1(n253), .A2(n232), .ZN(n230) );
  OAI21_X4 U274 ( .B1(n254), .B2(n232), .A(n233), .ZN(n231) );
  NAND2_X4 U275 ( .A1(n242), .A2(n234), .ZN(n232) );
  AOI21_X4 U276 ( .B1(n234), .B2(n243), .A(n235), .ZN(n233) );
  NOR2_X4 U277 ( .A1(n239), .A2(n236), .ZN(n234) );
  OAI21_X4 U278 ( .B1(n236), .B2(n240), .A(n237), .ZN(n235) );
  NAND2_X4 U279 ( .A1(n391), .A2(n237), .ZN(n34) );
  NOR2_X4 U281 ( .A1(B[23]), .A2(A[23]), .ZN(n236) );
  NAND2_X4 U282 ( .A1(B[23]), .A2(A[23]), .ZN(n237) );
  XOR2_X2 U283 ( .A(n241), .B(n35), .Z(SUM[22]) );
  OAI21_X4 U284 ( .B1(n241), .B2(n239), .A(n240), .ZN(n238) );
  NAND2_X4 U285 ( .A1(n392), .A2(n240), .ZN(n35) );
  NOR2_X4 U287 ( .A1(B[22]), .A2(A[22]), .ZN(n239) );
  NAND2_X4 U288 ( .A1(B[22]), .A2(A[22]), .ZN(n240) );
  XNOR2_X2 U289 ( .A(n246), .B(n36), .ZN(SUM[21]) );
  AOI21_X4 U290 ( .B1(n249), .B2(n242), .A(n243), .ZN(n241) );
  NOR2_X4 U291 ( .A1(n247), .A2(n244), .ZN(n242) );
  OAI21_X4 U292 ( .B1(n244), .B2(n248), .A(n245), .ZN(n243) );
  NAND2_X4 U293 ( .A1(n393), .A2(n245), .ZN(n36) );
  NOR2_X4 U295 ( .A1(B[21]), .A2(A[21]), .ZN(n244) );
  NAND2_X4 U296 ( .A1(B[21]), .A2(A[21]), .ZN(n245) );
  XNOR2_X2 U297 ( .A(n249), .B(n37), .ZN(SUM[20]) );
  OAI21_X4 U298 ( .B1(n250), .B2(n247), .A(n248), .ZN(n246) );
  NAND2_X4 U299 ( .A1(n394), .A2(n248), .ZN(n37) );
  NOR2_X4 U301 ( .A1(B[20]), .A2(A[20]), .ZN(n247) );
  NAND2_X4 U302 ( .A1(B[20]), .A2(A[20]), .ZN(n248) );
  XNOR2_X2 U303 ( .A(n259), .B(n38), .ZN(SUM[19]) );
  AOI21_X4 U305 ( .B1(n272), .B2(n251), .A(n252), .ZN(n250) );
  NAND2_X4 U308 ( .A1(n263), .A2(n255), .ZN(n253) );
  AOI21_X4 U309 ( .B1(n255), .B2(n264), .A(n256), .ZN(n254) );
  NOR2_X4 U310 ( .A1(n260), .A2(n257), .ZN(n255) );
  OAI21_X4 U311 ( .B1(n257), .B2(n261), .A(n258), .ZN(n256) );
  NAND2_X4 U312 ( .A1(n395), .A2(n258), .ZN(n38) );
  NOR2_X4 U314 ( .A1(B[19]), .A2(A[19]), .ZN(n257) );
  NAND2_X4 U315 ( .A1(B[19]), .A2(A[19]), .ZN(n258) );
  XOR2_X2 U316 ( .A(n262), .B(n39), .Z(SUM[18]) );
  OAI21_X4 U317 ( .B1(n262), .B2(n260), .A(n261), .ZN(n259) );
  NAND2_X4 U318 ( .A1(n396), .A2(n261), .ZN(n39) );
  NOR2_X4 U320 ( .A1(B[18]), .A2(A[18]), .ZN(n260) );
  NAND2_X4 U321 ( .A1(B[18]), .A2(A[18]), .ZN(n261) );
  XOR2_X2 U322 ( .A(n267), .B(n40), .Z(SUM[17]) );
  AOI21_X4 U323 ( .B1(n272), .B2(n263), .A(n264), .ZN(n262) );
  NOR2_X4 U324 ( .A1(n270), .A2(n265), .ZN(n263) );
  OAI21_X4 U325 ( .B1(n265), .B2(n271), .A(n266), .ZN(n264) );
  NAND2_X4 U326 ( .A1(n397), .A2(n266), .ZN(n40) );
  NOR2_X4 U328 ( .A1(B[17]), .A2(A[17]), .ZN(n265) );
  NAND2_X4 U329 ( .A1(B[17]), .A2(A[17]), .ZN(n266) );
  XNOR2_X2 U330 ( .A(n272), .B(n41), .ZN(SUM[16]) );
  AOI21_X4 U331 ( .B1(n272), .B2(n398), .A(n269), .ZN(n267) );
  NAND2_X4 U334 ( .A1(n398), .A2(n271), .ZN(n41) );
  NOR2_X4 U336 ( .A1(B[16]), .A2(A[16]), .ZN(n270) );
  NAND2_X4 U337 ( .A1(B[16]), .A2(A[16]), .ZN(n271) );
  XOR2_X2 U338 ( .A(n282), .B(n42), .Z(SUM[15]) );
  AOI21_X4 U340 ( .B1(n323), .B2(n274), .A(n275), .ZN(n273) );
  NOR2_X4 U341 ( .A1(n301), .A2(n276), .ZN(n274) );
  NAND2_X4 U343 ( .A1(n290), .A2(n278), .ZN(n276) );
  AOI21_X4 U344 ( .B1(n278), .B2(n291), .A(n279), .ZN(n277) );
  NOR2_X4 U345 ( .A1(n285), .A2(n280), .ZN(n278) );
  OAI21_X4 U346 ( .B1(n280), .B2(n286), .A(n281), .ZN(n279) );
  NAND2_X4 U347 ( .A1(n399), .A2(n281), .ZN(n42) );
  NOR2_X4 U349 ( .A1(B[15]), .A2(A[15]), .ZN(n280) );
  NAND2_X4 U350 ( .A1(B[15]), .A2(A[15]), .ZN(n281) );
  XNOR2_X2 U351 ( .A(n287), .B(n43), .ZN(SUM[14]) );
  AOI21_X4 U352 ( .B1(n287), .B2(n400), .A(n284), .ZN(n282) );
  NAND2_X4 U355 ( .A1(n400), .A2(n286), .ZN(n43) );
  NOR2_X4 U357 ( .A1(B[14]), .A2(A[14]), .ZN(n285) );
  NAND2_X4 U358 ( .A1(B[14]), .A2(A[14]), .ZN(n286) );
  XOR2_X2 U359 ( .A(n294), .B(n44), .Z(SUM[13]) );
  OAI21_X4 U360 ( .B1(n299), .B2(n288), .A(n289), .ZN(n287) );
  NOR2_X4 U363 ( .A1(n297), .A2(n292), .ZN(n290) );
  OAI21_X4 U364 ( .B1(n292), .B2(n298), .A(n293), .ZN(n291) );
  NAND2_X4 U365 ( .A1(n401), .A2(n293), .ZN(n44) );
  NOR2_X4 U367 ( .A1(B[13]), .A2(A[13]), .ZN(n292) );
  NAND2_X4 U368 ( .A1(B[13]), .A2(A[13]), .ZN(n293) );
  XOR2_X2 U369 ( .A(n299), .B(n45), .Z(SUM[12]) );
  AOI21_X4 U370 ( .B1(n300), .B2(n402), .A(n296), .ZN(n294) );
  NAND2_X4 U373 ( .A1(n402), .A2(n298), .ZN(n45) );
  NOR2_X4 U375 ( .A1(B[12]), .A2(A[12]), .ZN(n297) );
  NAND2_X4 U376 ( .A1(B[12]), .A2(A[12]), .ZN(n298) );
  XOR2_X2 U377 ( .A(n307), .B(n46), .Z(SUM[11]) );
  NAND2_X4 U380 ( .A1(n315), .A2(n303), .ZN(n301) );
  AOI21_X4 U381 ( .B1(n303), .B2(n316), .A(n304), .ZN(n302) );
  NOR2_X4 U382 ( .A1(n310), .A2(n305), .ZN(n303) );
  OAI21_X4 U383 ( .B1(n305), .B2(n311), .A(n306), .ZN(n304) );
  NAND2_X4 U384 ( .A1(n403), .A2(n306), .ZN(n46) );
  NOR2_X4 U386 ( .A1(B[11]), .A2(A[11]), .ZN(n305) );
  XNOR2_X2 U388 ( .A(n312), .B(n47), .ZN(SUM[10]) );
  AOI21_X4 U389 ( .B1(n312), .B2(n404), .A(n309), .ZN(n307) );
  NAND2_X4 U392 ( .A1(n404), .A2(n311), .ZN(n47) );
  NOR2_X4 U394 ( .A1(B[10]), .A2(A[10]), .ZN(n310) );
  NAND2_X4 U395 ( .A1(B[10]), .A2(A[10]), .ZN(n311) );
  XNOR2_X2 U396 ( .A(n319), .B(n48), .ZN(SUM[9]) );
  OAI21_X4 U397 ( .B1(n322), .B2(n313), .A(n314), .ZN(n312) );
  NOR2_X4 U400 ( .A1(n320), .A2(n317), .ZN(n315) );
  OAI21_X4 U401 ( .B1(n317), .B2(n321), .A(n318), .ZN(n316) );
  NAND2_X4 U402 ( .A1(n405), .A2(n318), .ZN(n48) );
  NOR2_X4 U404 ( .A1(B[9]), .A2(A[9]), .ZN(n317) );
  NAND2_X4 U405 ( .A1(B[9]), .A2(A[9]), .ZN(n318) );
  XOR2_X2 U406 ( .A(n322), .B(n49), .Z(SUM[8]) );
  OAI21_X4 U407 ( .B1(n322), .B2(n320), .A(n321), .ZN(n319) );
  NAND2_X4 U408 ( .A1(n406), .A2(n321), .ZN(n49) );
  NOR2_X4 U410 ( .A1(B[8]), .A2(A[8]), .ZN(n320) );
  NAND2_X4 U411 ( .A1(B[8]), .A2(A[8]), .ZN(n321) );
  XNOR2_X2 U412 ( .A(n330), .B(n50), .ZN(SUM[7]) );
  OAI21_X4 U414 ( .B1(n344), .B2(n324), .A(n325), .ZN(n323) );
  NAND2_X4 U415 ( .A1(n334), .A2(n326), .ZN(n324) );
  AOI21_X4 U416 ( .B1(n326), .B2(n335), .A(n327), .ZN(n325) );
  NOR2_X4 U417 ( .A1(n331), .A2(n328), .ZN(n326) );
  OAI21_X4 U418 ( .B1(n328), .B2(n332), .A(n329), .ZN(n327) );
  NAND2_X4 U419 ( .A1(n407), .A2(n329), .ZN(n50) );
  NOR2_X4 U421 ( .A1(B[7]), .A2(A[7]), .ZN(n328) );
  NAND2_X4 U422 ( .A1(B[7]), .A2(A[7]), .ZN(n329) );
  XOR2_X2 U423 ( .A(n333), .B(n51), .Z(SUM[6]) );
  OAI21_X4 U424 ( .B1(n333), .B2(n331), .A(n332), .ZN(n330) );
  NAND2_X4 U425 ( .A1(n408), .A2(n332), .ZN(n51) );
  NOR2_X4 U427 ( .A1(B[6]), .A2(A[6]), .ZN(n331) );
  NAND2_X4 U428 ( .A1(B[6]), .A2(A[6]), .ZN(n332) );
  XOR2_X2 U429 ( .A(n338), .B(n52), .Z(SUM[5]) );
  AOI21_X4 U430 ( .B1(n343), .B2(n334), .A(n335), .ZN(n333) );
  NOR2_X4 U431 ( .A1(n341), .A2(n336), .ZN(n334) );
  OAI21_X4 U432 ( .B1(n336), .B2(n342), .A(n337), .ZN(n335) );
  NAND2_X4 U433 ( .A1(n409), .A2(n337), .ZN(n52) );
  NOR2_X4 U435 ( .A1(B[5]), .A2(A[5]), .ZN(n336) );
  NAND2_X4 U436 ( .A1(B[5]), .A2(A[5]), .ZN(n337) );
  XNOR2_X2 U437 ( .A(n343), .B(n53), .ZN(SUM[4]) );
  AOI21_X4 U438 ( .B1(n343), .B2(n410), .A(n340), .ZN(n338) );
  NAND2_X4 U441 ( .A1(n410), .A2(n342), .ZN(n53) );
  NOR2_X4 U443 ( .A1(B[4]), .A2(A[4]), .ZN(n341) );
  NAND2_X4 U444 ( .A1(B[4]), .A2(A[4]), .ZN(n342) );
  XNOR2_X2 U445 ( .A(n349), .B(n54), .ZN(SUM[3]) );
  AOI21_X4 U447 ( .B1(n345), .B2(n353), .A(n346), .ZN(n344) );
  NOR2_X4 U448 ( .A1(n350), .A2(n347), .ZN(n345) );
  OAI21_X4 U449 ( .B1(n347), .B2(n351), .A(n348), .ZN(n346) );
  NAND2_X4 U450 ( .A1(n411), .A2(n348), .ZN(n54) );
  NOR2_X4 U452 ( .A1(B[3]), .A2(A[3]), .ZN(n347) );
  NAND2_X4 U453 ( .A1(B[3]), .A2(A[3]), .ZN(n348) );
  XOR2_X2 U454 ( .A(n352), .B(n55), .Z(SUM[2]) );
  OAI21_X4 U455 ( .B1(n352), .B2(n350), .A(n351), .ZN(n349) );
  NAND2_X4 U456 ( .A1(n412), .A2(n351), .ZN(n55) );
  NOR2_X4 U458 ( .A1(B[2]), .A2(A[2]), .ZN(n350) );
  NAND2_X4 U459 ( .A1(B[2]), .A2(A[2]), .ZN(n351) );
  XOR2_X2 U460 ( .A(n56), .B(n357), .Z(SUM[1]) );
  OAI21_X4 U462 ( .B1(n354), .B2(n357), .A(n355), .ZN(n353) );
  NAND2_X4 U463 ( .A1(n413), .A2(n355), .ZN(n56) );
  NOR2_X4 U465 ( .A1(B[1]), .A2(A[1]), .ZN(n354) );
  NAND2_X4 U466 ( .A1(B[1]), .A2(A[1]), .ZN(n355) );
  NAND2_X4 U468 ( .A1(n414), .A2(n357), .ZN(n57) );
  NOR2_X4 U470 ( .A1(B[0]), .A2(A[0]), .ZN(n356) );
  NAND2_X4 U471 ( .A1(B[0]), .A2(A[0]), .ZN(n357) );
  XNOR2_X1 U475 ( .A(n70), .B(n2), .ZN(SUM[55]) );
  XNOR2_X1 U476 ( .A(n118), .B(n14), .ZN(SUM[43]) );
  XOR2_X1 U477 ( .A(n105), .B(n11), .Z(SUM[46]) );
  INV_X1 U478 ( .A(n65), .ZN(n358) );
  AOI21_X2 U479 ( .B1(n70), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X2 U480 ( .B1(n105), .B2(n103), .A(n104), .ZN(n102) );
  XOR2_X1 U481 ( .A(n121), .B(n15), .Z(SUM[42]) );
  XOR2_X1 U482 ( .A(n73), .B(n3), .Z(SUM[54]) );
  OAI21_X1 U483 ( .B1(n184), .B2(n127), .A(n128), .ZN(n126) );
  OAI21_X2 U484 ( .B1(n73), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X2 U485 ( .B1(n121), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U486 ( .B1(n128), .B2(n124), .A(n125), .ZN(n123) );
  XNOR2_X1 U487 ( .A(n86), .B(n6), .ZN(SUM[51]) );
  XNOR2_X1 U488 ( .A(n94), .B(n8), .ZN(SUM[49]) );
  OAI21_X1 U489 ( .B1(n322), .B2(n301), .A(n302), .ZN(n300) );
  OAI21_X1 U490 ( .B1(n302), .B2(n276), .A(n277), .ZN(n275) );
  NAND2_X1 U491 ( .A1(B[11]), .A2(A[11]), .ZN(n306) );
  OAI21_X2 U492 ( .B1(n97), .B2(n95), .A(n96), .ZN(n94) );
  OAI21_X2 U493 ( .B1(n89), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X2 U494 ( .B1(n167), .B2(n173), .A(n168), .ZN(n166) );
  OAI21_X2 U495 ( .B1(n179), .B2(n183), .A(n180), .ZN(n178) );
  XOR2_X1 U496 ( .A(n58), .B(n1), .Z(SUM[63]) );
  INV_X2 U497 ( .A(n101), .ZN(n99) );
  INV_X2 U498 ( .A(n93), .ZN(n91) );
  INV_X2 U499 ( .A(n85), .ZN(n83) );
  INV_X2 U500 ( .A(n77), .ZN(n75) );
  INV_X2 U501 ( .A(n69), .ZN(n67) );
  INV_X2 U502 ( .A(n356), .ZN(n414) );
  INV_X2 U503 ( .A(n354), .ZN(n413) );
  INV_X2 U504 ( .A(n350), .ZN(n412) );
  INV_X2 U505 ( .A(n347), .ZN(n411) );
  INV_X2 U506 ( .A(n336), .ZN(n409) );
  INV_X2 U507 ( .A(n331), .ZN(n408) );
  INV_X2 U508 ( .A(n328), .ZN(n407) );
  INV_X2 U509 ( .A(n320), .ZN(n406) );
  INV_X2 U510 ( .A(n317), .ZN(n405) );
  INV_X2 U511 ( .A(n305), .ZN(n403) );
  INV_X2 U512 ( .A(n292), .ZN(n401) );
  INV_X2 U513 ( .A(n280), .ZN(n399) );
  INV_X2 U514 ( .A(n265), .ZN(n397) );
  INV_X2 U515 ( .A(n260), .ZN(n396) );
  INV_X2 U516 ( .A(n257), .ZN(n395) );
  INV_X2 U517 ( .A(n247), .ZN(n394) );
  INV_X2 U518 ( .A(n244), .ZN(n393) );
  INV_X2 U519 ( .A(n239), .ZN(n392) );
  INV_X2 U520 ( .A(n236), .ZN(n391) );
  INV_X2 U521 ( .A(n226), .ZN(n390) );
  INV_X2 U522 ( .A(n223), .ZN(n389) );
  INV_X2 U523 ( .A(n218), .ZN(n388) );
  INV_X2 U524 ( .A(n215), .ZN(n387) );
  INV_X2 U525 ( .A(n205), .ZN(n386) );
  INV_X2 U526 ( .A(n202), .ZN(n385) );
  INV_X2 U527 ( .A(n197), .ZN(n384) );
  INV_X2 U528 ( .A(n194), .ZN(n383) );
  INV_X2 U529 ( .A(n182), .ZN(n382) );
  INV_X2 U530 ( .A(n179), .ZN(n381) );
  INV_X2 U531 ( .A(n167), .ZN(n379) );
  INV_X2 U532 ( .A(n154), .ZN(n377) );
  INV_X2 U533 ( .A(n142), .ZN(n375) );
  INV_X2 U534 ( .A(n124), .ZN(n373) );
  INV_X2 U535 ( .A(n119), .ZN(n372) );
  INV_X2 U536 ( .A(n111), .ZN(n370) );
  INV_X2 U537 ( .A(n103), .ZN(n368) );
  INV_X2 U538 ( .A(n100), .ZN(n98) );
  INV_X2 U539 ( .A(n95), .ZN(n366) );
  INV_X2 U540 ( .A(n92), .ZN(n90) );
  INV_X2 U541 ( .A(n87), .ZN(n364) );
  INV_X2 U542 ( .A(n84), .ZN(n82) );
  INV_X2 U543 ( .A(n79), .ZN(n362) );
  INV_X2 U544 ( .A(n76), .ZN(n74) );
  INV_X2 U545 ( .A(n71), .ZN(n360) );
  INV_X2 U546 ( .A(n68), .ZN(n66) );
  INV_X2 U547 ( .A(n353), .ZN(n352) );
  INV_X2 U548 ( .A(n344), .ZN(n343) );
  INV_X2 U549 ( .A(n342), .ZN(n340) );
  INV_X2 U550 ( .A(n341), .ZN(n410) );
  INV_X2 U551 ( .A(n323), .ZN(n322) );
  INV_X2 U552 ( .A(n316), .ZN(n314) );
  INV_X2 U553 ( .A(n315), .ZN(n313) );
  INV_X2 U554 ( .A(n311), .ZN(n309) );
  INV_X2 U555 ( .A(n310), .ZN(n404) );
  INV_X2 U556 ( .A(n300), .ZN(n299) );
  INV_X2 U557 ( .A(n298), .ZN(n296) );
  INV_X2 U558 ( .A(n297), .ZN(n402) );
  INV_X2 U559 ( .A(n291), .ZN(n289) );
  INV_X2 U560 ( .A(n290), .ZN(n288) );
  INV_X2 U561 ( .A(n286), .ZN(n284) );
  INV_X2 U562 ( .A(n285), .ZN(n400) );
  INV_X2 U563 ( .A(n273), .ZN(n272) );
  INV_X2 U564 ( .A(n271), .ZN(n269) );
  INV_X2 U565 ( .A(n270), .ZN(n398) );
  INV_X2 U566 ( .A(n254), .ZN(n252) );
  INV_X2 U567 ( .A(n253), .ZN(n251) );
  INV_X2 U568 ( .A(n250), .ZN(n249) );
  INV_X2 U569 ( .A(n229), .ZN(n228) );
  INV_X2 U570 ( .A(n212), .ZN(n210) );
  INV_X2 U571 ( .A(n211), .ZN(n209) );
  INV_X2 U572 ( .A(n208), .ZN(n207) );
  INV_X2 U573 ( .A(n185), .ZN(n184) );
  INV_X2 U574 ( .A(n178), .ZN(n176) );
  INV_X2 U575 ( .A(n177), .ZN(n175) );
  INV_X2 U576 ( .A(n173), .ZN(n171) );
  INV_X2 U577 ( .A(n172), .ZN(n380) );
  INV_X2 U578 ( .A(n162), .ZN(n161) );
  INV_X2 U579 ( .A(n160), .ZN(n158) );
  INV_X2 U580 ( .A(n159), .ZN(n378) );
  INV_X2 U581 ( .A(n153), .ZN(n151) );
  INV_X2 U582 ( .A(n152), .ZN(n150) );
  INV_X2 U583 ( .A(n148), .ZN(n146) );
  INV_X2 U584 ( .A(n147), .ZN(n376) );
  INV_X2 U585 ( .A(n137), .ZN(n135) );
  INV_X2 U586 ( .A(n136), .ZN(n134) );
  INV_X2 U587 ( .A(n132), .ZN(n130) );
  INV_X2 U588 ( .A(n131), .ZN(n374) );
  INV_X2 U589 ( .A(n117), .ZN(n115) );
  INV_X2 U590 ( .A(n116), .ZN(n371) );
  INV_X2 U591 ( .A(n109), .ZN(n107) );
  INV_X2 U592 ( .A(n108), .ZN(n369) );
  INV_X2 U593 ( .A(n57), .ZN(SUM[0]) );
endmodule


module up_island_DW01_add_4 ( A, B, SUM, CI, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n42, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n56, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n105, n106, n107, n108, n110, n111, n112, n113,
         n114, n115, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n130, n131, n132, n133, n134, n135, n138, n139, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157,
         n158, n159, n160, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n191, n192, n193, n194, n195,
         n196, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n213, n214, n215, n216, n217, n218, n219, n220,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n235, n236, n237, n238, n239, n240, n242, n243, n244, n245, n246,
         n247, n248, n249, n252, n253, n254, n255, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n285, n286, n287, n288,
         n289, n290, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n329,
         n331, n332, n333, n334, n335, n336, n340, n341, n342, n343, n345,
         n347, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524;

  NAND2_X4 U6 ( .A1(n364), .A2(n38), .ZN(n5) );
  NAND2_X4 U20 ( .A1(n46), .A2(n49), .ZN(n6) );
  AOI21_X4 U35 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NAND2_X4 U38 ( .A1(n61), .A2(n64), .ZN(n7) );
  NAND2_X4 U44 ( .A1(n77), .A2(n70), .ZN(n66) );
  NAND2_X4 U50 ( .A1(n70), .A2(n73), .ZN(n8) );
  XNOR2_X2 U54 ( .A(n87), .B(n9), .ZN(SUM[27]) );
  NAND2_X4 U66 ( .A1(n83), .A2(n86), .ZN(n9) );
  XNOR2_X2 U70 ( .A(n96), .B(n10), .ZN(SUM[26]) );
  NAND2_X4 U78 ( .A1(n369), .A2(n95), .ZN(n10) );
  XNOR2_X2 U82 ( .A(n113), .B(n11), .ZN(SUM[25]) );
  NAND2_X4 U84 ( .A1(n391), .A2(n99), .ZN(n97) );
  AOI21_X4 U85 ( .B1(n347), .B2(n99), .A(n100), .ZN(n98) );
  NOR2_X4 U92 ( .A1(n107), .A2(n131), .ZN(n105) );
  AOI21_X4 U95 ( .B1(n370), .B2(n119), .A(n110), .ZN(n108) );
  NAND2_X4 U98 ( .A1(n370), .A2(n112), .ZN(n11) );
  XNOR2_X2 U102 ( .A(n122), .B(n12), .ZN(SUM[24]) );
  XNOR2_X2 U114 ( .A(n133), .B(n13), .ZN(SUM[23]) );
  NOR2_X4 U118 ( .A1(n4), .A2(n127), .ZN(n125) );
  OAI21_X4 U119 ( .B1(n345), .B2(n127), .A(n128), .ZN(n126) );
  XNOR2_X2 U128 ( .A(n146), .B(n14), .ZN(SUM[22]) );
  NAND2_X4 U140 ( .A1(n373), .A2(n145), .ZN(n14) );
  XNOR2_X2 U144 ( .A(n157), .B(n15), .ZN(SUM[21]) );
  NAND2_X4 U146 ( .A1(n391), .A2(n149), .ZN(n147) );
  AOI21_X4 U147 ( .B1(n347), .B2(n149), .A(n150), .ZN(n148) );
  NAND2_X4 U154 ( .A1(n374), .A2(n156), .ZN(n15) );
  NAND2_X4 U174 ( .A1(n375), .A2(n173), .ZN(n16) );
  XNOR2_X2 U178 ( .A(n181), .B(n17), .ZN(SUM[19]) );
  NAND2_X4 U180 ( .A1(n184), .A2(n376), .ZN(n175) );
  AOI21_X4 U181 ( .B1(n185), .B2(n376), .A(n178), .ZN(n176) );
  NAND2_X4 U184 ( .A1(n376), .A2(n180), .ZN(n17) );
  NOR2_X4 U192 ( .A1(n4), .A2(n186), .ZN(n184) );
  OAI21_X4 U193 ( .B1(n345), .B2(n186), .A(n187), .ZN(n185) );
  XNOR2_X2 U204 ( .A(n201), .B(n19), .ZN(SUM[17]) );
  NAND2_X4 U206 ( .A1(n204), .A2(n378), .ZN(n195) );
  AOI21_X4 U207 ( .B1(n205), .B2(n378), .A(n198), .ZN(n196) );
  NAND2_X4 U210 ( .A1(n378), .A2(n200), .ZN(n19) );
  XNOR2_X2 U214 ( .A(n218), .B(n20), .ZN(SUM[16]) );
  NOR2_X4 U218 ( .A1(n4), .A2(n206), .ZN(n204) );
  OAI21_X4 U219 ( .B1(n345), .B2(n206), .A(n207), .ZN(n205) );
  NAND2_X4 U230 ( .A1(n379), .A2(n217), .ZN(n20) );
  XNOR2_X2 U234 ( .A(n225), .B(n21), .ZN(SUM[15]) );
  NAND2_X4 U236 ( .A1(n228), .A2(n380), .ZN(n219) );
  AOI21_X4 U237 ( .B1(n229), .B2(n380), .A(n222), .ZN(n220) );
  NAND2_X4 U240 ( .A1(n380), .A2(n224), .ZN(n21) );
  XNOR2_X2 U244 ( .A(n238), .B(n22), .ZN(SUM[14]) );
  NOR2_X4 U248 ( .A1(n4), .A2(n230), .ZN(n228) );
  OAI21_X4 U249 ( .B1(n345), .B2(n230), .A(n231), .ZN(n229) );
  NAND2_X4 U256 ( .A1(n381), .A2(n237), .ZN(n22) );
  XNOR2_X2 U260 ( .A(n245), .B(n23), .ZN(SUM[13]) );
  NAND2_X4 U262 ( .A1(n248), .A2(n382), .ZN(n239) );
  AOI21_X4 U263 ( .B1(n249), .B2(n382), .A(n242), .ZN(n240) );
  XNOR2_X2 U270 ( .A(n268), .B(n24), .ZN(SUM[12]) );
  NAND2_X4 U292 ( .A1(n383), .A2(n267), .ZN(n24) );
  XNOR2_X2 U296 ( .A(n275), .B(n25), .ZN(SUM[11]) );
  NAND2_X4 U298 ( .A1(n278), .A2(n384), .ZN(n269) );
  AOI21_X4 U299 ( .B1(n279), .B2(n384), .A(n272), .ZN(n270) );
  XNOR2_X2 U306 ( .A(n288), .B(n26), .ZN(SUM[10]) );
  NAND2_X4 U318 ( .A1(n385), .A2(n287), .ZN(n26) );
  XNOR2_X2 U322 ( .A(n295), .B(n27), .ZN(SUM[9]) );
  NAND2_X4 U324 ( .A1(n298), .A2(n386), .ZN(n289) );
  AOI21_X4 U325 ( .B1(n299), .B2(n386), .A(n292), .ZN(n290) );
  XNOR2_X2 U332 ( .A(n314), .B(n28), .ZN(SUM[8]) );
  NAND2_X4 U350 ( .A1(n387), .A2(n313), .ZN(n28) );
  XNOR2_X2 U354 ( .A(n321), .B(n29), .ZN(SUM[7]) );
  NAND2_X4 U356 ( .A1(n324), .A2(n388), .ZN(n315) );
  AOI21_X4 U357 ( .B1(n325), .B2(n388), .A(n318), .ZN(n316) );
  XNOR2_X2 U364 ( .A(n334), .B(n30), .ZN(SUM[6]) );
  NOR2_X4 U368 ( .A1(n4), .A2(n326), .ZN(n324) );
  XNOR2_X2 U380 ( .A(n343), .B(n31), .ZN(SUM[5]) );
  NAND2_X4 U382 ( .A1(n391), .A2(n390), .ZN(n335) );
  AOI21_X4 U383 ( .B1(n347), .B2(n390), .A(n340), .ZN(n336) );
  NAND2_X4 U388 ( .A1(n390), .A2(n342), .ZN(n31) );
  NAND2_X4 U398 ( .A1(n391), .A2(n345), .ZN(n32) );
  NOR2_X4 U400 ( .A1(B[4]), .A2(A[4]), .ZN(n4) );
  NAND2_X4 U401 ( .A1(B[4]), .A2(A[4]), .ZN(n345) );
  XNOR2_X2 U402 ( .A(n355), .B(n33), .ZN(SUM[3]) );
  AOI21_X4 U403 ( .B1(n351), .B2(n359), .A(n352), .ZN(n2) );
  NOR2_X4 U404 ( .A1(n356), .A2(n353), .ZN(n351) );
  OAI21_X4 U405 ( .B1(n357), .B2(n353), .A(n354), .ZN(n352) );
  NAND2_X4 U406 ( .A1(n392), .A2(n354), .ZN(n33) );
  XOR2_X2 U410 ( .A(n34), .B(n358), .Z(SUM[2]) );
  OAI21_X4 U411 ( .B1(n358), .B2(n356), .A(n357), .ZN(n355) );
  NAND2_X4 U412 ( .A1(n393), .A2(n357), .ZN(n34) );
  XOR2_X2 U416 ( .A(n35), .B(n363), .Z(SUM[1]) );
  OAI21_X4 U418 ( .B1(n360), .B2(n363), .A(n361), .ZN(n359) );
  NAND2_X4 U419 ( .A1(n394), .A2(n361), .ZN(n35) );
  NAND2_X4 U424 ( .A1(n395), .A2(n363), .ZN(n36) );
  NAND2_X1 U431 ( .A1(A[29]), .A2(B[29]), .ZN(n64) );
  NOR2_X1 U432 ( .A1(B[8]), .A2(A[8]), .ZN(n312) );
  XNOR2_X1 U433 ( .A(n174), .B(n16), .ZN(SUM[20]) );
  NOR2_X1 U434 ( .A1(A[29]), .A2(B[29]), .ZN(n63) );
  INV_X1 U435 ( .A(n78), .ZN(n76) );
  AOI21_X1 U436 ( .B1(n78), .B2(n70), .A(n71), .ZN(n67) );
  AOI21_X1 U437 ( .B1(n285), .B2(n264), .A(n265), .ZN(n263) );
  AOI21_X2 U438 ( .B1(n214), .B2(n235), .A(n215), .ZN(n213) );
  AOI21_X1 U439 ( .B1(n170), .B2(n191), .A(n171), .ZN(n169) );
  NOR2_X1 U440 ( .A1(n179), .A2(n172), .ZN(n170) );
  CLKBUF_X1 U441 ( .A(n255), .Z(n498) );
  NOR2_X1 U442 ( .A1(n243), .A2(n236), .ZN(n232) );
  NOR2_X1 U443 ( .A1(n199), .A2(n192), .ZN(n188) );
  INV_X1 U444 ( .A(n253), .ZN(n499) );
  AOI21_X2 U445 ( .B1(n303), .B2(n260), .A(n261), .ZN(n255) );
  NOR2_X1 U446 ( .A1(B[0]), .A2(A[0]), .ZN(n362) );
  NAND2_X1 U447 ( .A1(B[0]), .A2(A[0]), .ZN(n363) );
  NOR2_X1 U448 ( .A1(B[2]), .A2(A[2]), .ZN(n356) );
  NAND2_X1 U449 ( .A1(B[2]), .A2(A[2]), .ZN(n357) );
  INV_X1 U450 ( .A(n302), .ZN(n300) );
  NOR2_X1 U451 ( .A1(n4), .A2(n300), .ZN(n298) );
  OAI21_X1 U452 ( .B1(n345), .B2(n300), .A(n301), .ZN(n299) );
  NOR2_X1 U453 ( .A1(n4), .A2(n280), .ZN(n278) );
  OAI21_X1 U454 ( .B1(n345), .B2(n280), .A(n281), .ZN(n279) );
  NOR2_X4 U455 ( .A1(A[10]), .A2(B[10]), .ZN(n286) );
  NOR2_X2 U456 ( .A1(n308), .A2(n326), .ZN(n302) );
  BUF_X2 U457 ( .A(n216), .Z(n500) );
  CLKBUF_X1 U458 ( .A(n320), .Z(n501) );
  INV_X1 U459 ( .A(n310), .ZN(n308) );
  OAI21_X1 U460 ( .B1(n499), .B2(n164), .A(n165), .ZN(n502) );
  XNOR2_X1 U461 ( .A(n74), .B(n8), .ZN(SUM[28]) );
  CLKBUF_X1 U462 ( .A(n319), .Z(n503) );
  CLKBUF_X1 U463 ( .A(n232), .Z(n504) );
  CLKBUF_X1 U464 ( .A(n236), .Z(n505) );
  NOR2_X2 U465 ( .A1(A[12]), .A2(B[12]), .ZN(n266) );
  AOI21_X2 U466 ( .B1(n389), .B2(n340), .A(n331), .ZN(n329) );
  INV_X1 U467 ( .A(n274), .ZN(n272) );
  NAND2_X1 U468 ( .A1(n384), .A2(n274), .ZN(n25) );
  NOR2_X1 U469 ( .A1(n168), .A2(n210), .ZN(n166) );
  NAND2_X1 U470 ( .A1(n232), .A2(n214), .ZN(n210) );
  INV_X1 U471 ( .A(n244), .ZN(n242) );
  NAND2_X1 U472 ( .A1(n382), .A2(n244), .ZN(n23) );
  XNOR2_X1 U473 ( .A(n65), .B(n7), .ZN(SUM[29]) );
  OAI21_X1 U474 ( .B1(n213), .B2(n168), .A(n169), .ZN(n167) );
  OAI21_X1 U475 ( .B1(n236), .B2(n244), .A(n237), .ZN(n235) );
  OAI21_X2 U476 ( .B1(n308), .B2(n329), .A(n309), .ZN(n303) );
  INV_X1 U477 ( .A(n311), .ZN(n309) );
  NOR2_X2 U478 ( .A1(n164), .A2(n254), .ZN(n160) );
  CLKBUF_X1 U479 ( .A(n502), .Z(n506) );
  NAND2_X1 U480 ( .A1(n377), .A2(n193), .ZN(n18) );
  XNOR2_X1 U481 ( .A(n194), .B(n18), .ZN(SUM[18]) );
  NAND2_X1 U482 ( .A1(n208), .A2(n188), .ZN(n186) );
  NAND2_X1 U483 ( .A1(n188), .A2(n170), .ZN(n168) );
  NAND2_X1 U484 ( .A1(n388), .A2(n501), .ZN(n29) );
  INV_X1 U485 ( .A(n501), .ZN(n318) );
  OAI21_X1 U486 ( .B1(n312), .B2(n320), .A(n313), .ZN(n311) );
  INV_X1 U487 ( .A(n166), .ZN(n164) );
  CLKBUF_X1 U488 ( .A(n93), .Z(n507) );
  CLKBUF_X1 U489 ( .A(n152), .Z(n508) );
  AND2_X2 U490 ( .A1(n509), .A2(n160), .ZN(n138) );
  NOR2_X1 U491 ( .A1(n144), .A2(n155), .ZN(n509) );
  BUF_X2 U492 ( .A(n160), .Z(n510) );
  NOR2_X1 U493 ( .A1(n293), .A2(n286), .ZN(n282) );
  INV_X1 U494 ( .A(n151), .ZN(n149) );
  NAND2_X2 U495 ( .A1(n302), .A2(n260), .ZN(n254) );
  OAI21_X2 U496 ( .B1(n255), .B2(n164), .A(n165), .ZN(n163) );
  AOI21_X2 U497 ( .B1(n163), .B2(n374), .A(n154), .ZN(n152) );
  NAND2_X1 U498 ( .A1(n389), .A2(n333), .ZN(n30) );
  NAND2_X2 U499 ( .A1(n390), .A2(n389), .ZN(n326) );
  AND2_X1 U500 ( .A1(n45), .A2(n516), .ZN(n511) );
  CLKBUF_X1 U501 ( .A(n329), .Z(n513) );
  CLKBUF_X1 U502 ( .A(n303), .Z(n512) );
  NOR2_X1 U503 ( .A1(n273), .A2(n266), .ZN(n264) );
  NAND2_X1 U504 ( .A1(n514), .A2(n515), .ZN(n516) );
  INV_X1 U505 ( .A(n345), .ZN(n514) );
  INV_X1 U506 ( .A(n44), .ZN(n515) );
  AOI21_X1 U507 ( .B1(n56), .B2(n46), .A(n47), .ZN(n45) );
  CLKBUF_X1 U508 ( .A(n102), .Z(n517) );
  CLKBUF_X1 U509 ( .A(n139), .Z(n518) );
  INV_X1 U510 ( .A(n512), .ZN(n301) );
  NOR2_X2 U511 ( .A1(n223), .A2(n500), .ZN(n214) );
  OAI21_X1 U512 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  AOI21_X1 U513 ( .B1(n209), .B2(n188), .A(n191), .ZN(n187) );
  NAND2_X2 U514 ( .A1(B[5]), .A2(A[5]), .ZN(n342) );
  AOI21_X1 U515 ( .B1(n93), .B2(n83), .A(n84), .ZN(n82) );
  NOR2_X2 U516 ( .A1(A[18]), .A2(B[18]), .ZN(n192) );
  AOI21_X1 U517 ( .B1(n253), .B2(n504), .A(n235), .ZN(n231) );
  NAND2_X1 U518 ( .A1(n252), .A2(n504), .ZN(n230) );
  OAI21_X1 U519 ( .B1(n345), .B2(n326), .A(n513), .ZN(n325) );
  NAND2_X1 U520 ( .A1(A[30]), .A2(B[30]), .ZN(n49) );
  NOR2_X1 U521 ( .A1(A[30]), .A2(B[30]), .ZN(n48) );
  AND2_X1 U522 ( .A1(n46), .A2(n520), .ZN(n521) );
  INV_X4 U523 ( .A(n79), .ZN(n519) );
  INV_X1 U524 ( .A(n59), .ZN(n520) );
  AND2_X2 U525 ( .A1(n519), .A2(n520), .ZN(n53) );
  AND2_X1 U526 ( .A1(n83), .A2(n523), .ZN(n524) );
  INV_X4 U527 ( .A(n101), .ZN(n522) );
  INV_X1 U528 ( .A(n94), .ZN(n523) );
  AND2_X2 U529 ( .A1(n522), .A2(n523), .ZN(n90) );
  NAND2_X1 U530 ( .A1(n61), .A2(n70), .ZN(n59) );
  NAND2_X1 U531 ( .A1(B[1]), .A2(A[1]), .ZN(n361) );
  NOR2_X1 U532 ( .A1(B[1]), .A2(A[1]), .ZN(n360) );
  NAND2_X1 U533 ( .A1(n302), .A2(n282), .ZN(n280) );
  AOI21_X1 U534 ( .B1(n303), .B2(n282), .A(n285), .ZN(n281) );
  INV_X1 U535 ( .A(n101), .ZN(n99) );
  NAND2_X1 U536 ( .A1(n282), .A2(n264), .ZN(n262) );
  OAI21_X1 U537 ( .B1(n216), .B2(n224), .A(n217), .ZN(n215) );
  OAI21_X2 U538 ( .B1(n102), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X2 U539 ( .B1(n139), .B2(n105), .A(n106), .ZN(n102) );
  OAI21_X2 U540 ( .B1(n152), .B2(n144), .A(n145), .ZN(n139) );
  INV_X1 U541 ( .A(n263), .ZN(n261) );
  OAI21_X1 U542 ( .B1(n82), .B2(n59), .A(n60), .ZN(n56) );
  OAI21_X1 U543 ( .B1(n286), .B2(n294), .A(n287), .ZN(n285) );
  INV_X1 U544 ( .A(n508), .ZN(n150) );
  INV_X1 U545 ( .A(n517), .ZN(n100) );
  NOR2_X1 U546 ( .A1(n4), .A2(n254), .ZN(n248) );
  INV_X1 U547 ( .A(n254), .ZN(n252) );
  NOR2_X1 U548 ( .A1(n254), .A2(n210), .ZN(n208) );
  NAND2_X1 U549 ( .A1(A[28]), .A2(B[28]), .ZN(n73) );
  NOR2_X1 U550 ( .A1(A[28]), .A2(B[28]), .ZN(n72) );
  NOR2_X2 U551 ( .A1(n4), .A2(n79), .ZN(n77) );
  XOR2_X1 U552 ( .A(n2), .B(n32), .Z(SUM[4]) );
  OAI21_X1 U553 ( .B1(n2), .B2(n4), .A(n345), .ZN(n343) );
  OAI21_X1 U554 ( .B1(n2), .B2(n335), .A(n336), .ZN(n334) );
  OAI21_X1 U555 ( .B1(n2), .B2(n219), .A(n220), .ZN(n218) );
  OAI21_X1 U556 ( .B1(n2), .B2(n276), .A(n277), .ZN(n275) );
  OAI21_X1 U557 ( .B1(n2), .B2(n239), .A(n240), .ZN(n238) );
  OAI21_X1 U558 ( .B1(n2), .B2(n226), .A(n227), .ZN(n225) );
  OAI21_X1 U559 ( .B1(n2), .B2(n246), .A(n247), .ZN(n245) );
  OAI21_X1 U560 ( .B1(n2), .B2(n269), .A(n270), .ZN(n268) );
  OAI21_X1 U561 ( .B1(n2), .B2(n175), .A(n176), .ZN(n174) );
  OAI21_X1 U562 ( .B1(n2), .B2(n182), .A(n183), .ZN(n181) );
  OAI21_X1 U563 ( .B1(n2), .B2(n289), .A(n290), .ZN(n288) );
  OAI21_X1 U564 ( .B1(n2), .B2(n315), .A(n316), .ZN(n314) );
  OAI21_X1 U565 ( .B1(n2), .B2(n123), .A(n124), .ZN(n122) );
  OAI21_X1 U566 ( .B1(n2), .B2(n322), .A(n323), .ZN(n321) );
  OAI21_X1 U567 ( .B1(n2), .B2(n195), .A(n196), .ZN(n194) );
  OAI21_X1 U568 ( .B1(n2), .B2(n202), .A(n203), .ZN(n201) );
  OAI21_X1 U569 ( .B1(n2), .B2(n296), .A(n297), .ZN(n295) );
  OAI21_X1 U570 ( .B1(n2), .B2(n134), .A(n135), .ZN(n133) );
  OAI21_X1 U571 ( .B1(n2), .B2(n88), .A(n89), .ZN(n87) );
  OAI21_X1 U572 ( .B1(n2), .B2(n75), .A(n76), .ZN(n74) );
  OAI21_X1 U573 ( .B1(n2), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U574 ( .B1(n2), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U575 ( .B1(n2), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X1 U576 ( .B1(n2), .B2(n40), .A(n511), .ZN(n39) );
  OAI21_X1 U577 ( .B1(n2), .B2(n97), .A(n98), .ZN(n96) );
  OAI21_X1 U578 ( .B1(n2), .B2(n114), .A(n115), .ZN(n113) );
  NAND2_X1 U579 ( .A1(B[3]), .A2(A[3]), .ZN(n354) );
  NOR2_X1 U580 ( .A1(B[3]), .A2(A[3]), .ZN(n353) );
  NAND2_X1 U581 ( .A1(A[26]), .A2(B[26]), .ZN(n95) );
  NOR2_X1 U582 ( .A1(A[26]), .A2(B[26]), .ZN(n94) );
  NAND2_X1 U583 ( .A1(n386), .A2(n294), .ZN(n27) );
  INV_X1 U584 ( .A(n294), .ZN(n292) );
  NAND2_X1 U585 ( .A1(A[27]), .A2(B[27]), .ZN(n86) );
  NOR2_X1 U586 ( .A1(A[27]), .A2(B[27]), .ZN(n85) );
  NAND2_X1 U587 ( .A1(n391), .A2(n510), .ZN(n158) );
  AOI21_X1 U588 ( .B1(n347), .B2(n510), .A(n506), .ZN(n159) );
  NAND2_X2 U589 ( .A1(n510), .A2(n374), .ZN(n151) );
  OAI21_X1 U590 ( .B1(n345), .B2(n254), .A(n499), .ZN(n249) );
  INV_X1 U591 ( .A(n498), .ZN(n253) );
  AOI21_X1 U592 ( .B1(n518), .B2(n372), .A(n130), .ZN(n128) );
  OAI21_X1 U593 ( .B1(n498), .B2(n210), .A(n213), .ZN(n209) );
  OAI21_X1 U594 ( .B1(n345), .B2(n79), .A(n82), .ZN(n78) );
  OAI21_X1 U595 ( .B1(n266), .B2(n274), .A(n267), .ZN(n265) );
  NAND2_X1 U596 ( .A1(n372), .A2(n132), .ZN(n13) );
  INV_X1 U597 ( .A(n132), .ZN(n130) );
  OAI21_X2 U598 ( .B1(n107), .B2(n132), .A(n108), .ZN(n106) );
  NOR2_X1 U599 ( .A1(A[23]), .A2(B[23]), .ZN(n131) );
  NAND2_X1 U600 ( .A1(A[23]), .A2(B[23]), .ZN(n132) );
  XNOR2_X1 U601 ( .A(n50), .B(n6), .ZN(SUM[30]) );
  OAI21_X1 U602 ( .B1(n2), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U603 ( .A(n144), .ZN(n373) );
  NAND2_X1 U604 ( .A1(A[22]), .A2(B[22]), .ZN(n145) );
  NOR2_X1 U605 ( .A1(A[22]), .A2(B[22]), .ZN(n144) );
  NAND2_X1 U606 ( .A1(A[24]), .A2(B[24]), .ZN(n121) );
  NOR2_X1 U607 ( .A1(A[24]), .A2(B[24]), .ZN(n120) );
  NAND2_X1 U608 ( .A1(A[25]), .A2(B[25]), .ZN(n112) );
  NOR2_X1 U609 ( .A1(A[25]), .A2(B[25]), .ZN(n111) );
  NAND2_X1 U610 ( .A1(A[31]), .A2(B[31]), .ZN(n38) );
  NOR2_X1 U611 ( .A1(A[31]), .A2(B[31]), .ZN(n37) );
  NAND2_X1 U612 ( .A1(n371), .A2(n121), .ZN(n12) );
  NAND2_X1 U613 ( .A1(n125), .A2(n371), .ZN(n114) );
  AOI21_X1 U614 ( .B1(n126), .B2(n371), .A(n119), .ZN(n115) );
  NAND2_X2 U615 ( .A1(n370), .A2(n371), .ZN(n107) );
  INV_X1 U616 ( .A(n179), .ZN(n376) );
  NAND2_X1 U617 ( .A1(A[21]), .A2(B[21]), .ZN(n156) );
  NOR2_X1 U618 ( .A1(A[21]), .A2(B[21]), .ZN(n155) );
  NOR2_X1 U619 ( .A1(A[15]), .A2(B[15]), .ZN(n223) );
  INV_X1 U620 ( .A(n192), .ZN(n377) );
  NAND2_X1 U621 ( .A1(A[18]), .A2(B[18]), .ZN(n193) );
  OAI21_X2 U622 ( .B1(n192), .B2(n200), .A(n193), .ZN(n191) );
  NAND2_X1 U623 ( .A1(n521), .A2(n519), .ZN(n44) );
  NAND2_X1 U624 ( .A1(n391), .A2(n53), .ZN(n51) );
  AOI21_X1 U625 ( .B1(n347), .B2(n53), .A(n56), .ZN(n52) );
  NOR2_X1 U626 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U627 ( .A1(A[19]), .A2(B[19]), .ZN(n180) );
  NOR2_X1 U628 ( .A1(A[19]), .A2(B[19]), .ZN(n179) );
  NAND2_X1 U629 ( .A1(n138), .A2(n372), .ZN(n127) );
  NAND2_X1 U630 ( .A1(n391), .A2(n138), .ZN(n134) );
  NAND2_X2 U631 ( .A1(n138), .A2(n105), .ZN(n101) );
  AOI21_X1 U632 ( .B1(n347), .B2(n138), .A(n518), .ZN(n135) );
  NAND2_X2 U633 ( .A1(n524), .A2(n522), .ZN(n79) );
  NAND2_X1 U634 ( .A1(n391), .A2(n90), .ZN(n88) );
  AOI21_X1 U635 ( .B1(n347), .B2(n90), .A(n507), .ZN(n89) );
  NAND2_X1 U636 ( .A1(A[15]), .A2(B[15]), .ZN(n224) );
  INV_X1 U637 ( .A(n42), .ZN(n40) );
  INV_X1 U638 ( .A(n199), .ZN(n378) );
  NAND2_X1 U639 ( .A1(A[17]), .A2(B[17]), .ZN(n200) );
  NOR2_X1 U640 ( .A1(A[17]), .A2(B[17]), .ZN(n199) );
  INV_X1 U641 ( .A(n243), .ZN(n382) );
  NAND2_X1 U642 ( .A1(A[13]), .A2(B[13]), .ZN(n244) );
  NOR2_X1 U643 ( .A1(A[13]), .A2(B[13]), .ZN(n243) );
  INV_X1 U644 ( .A(n503), .ZN(n388) );
  NAND2_X1 U645 ( .A1(B[7]), .A2(A[7]), .ZN(n320) );
  NOR2_X1 U646 ( .A1(A[7]), .A2(B[7]), .ZN(n319) );
  INV_X1 U647 ( .A(n273), .ZN(n384) );
  NOR2_X1 U648 ( .A1(A[11]), .A2(B[11]), .ZN(n273) );
  NAND2_X1 U649 ( .A1(A[11]), .A2(B[11]), .ZN(n274) );
  INV_X1 U650 ( .A(n172), .ZN(n375) );
  NAND2_X1 U651 ( .A1(A[20]), .A2(B[20]), .ZN(n173) );
  NOR2_X1 U652 ( .A1(A[20]), .A2(B[20]), .ZN(n172) );
  INV_X1 U653 ( .A(n500), .ZN(n379) );
  NAND2_X1 U654 ( .A1(A[16]), .A2(B[16]), .ZN(n217) );
  NOR2_X1 U655 ( .A1(A[16]), .A2(B[16]), .ZN(n216) );
  INV_X1 U656 ( .A(n293), .ZN(n386) );
  NOR2_X1 U657 ( .A1(A[9]), .A2(B[9]), .ZN(n293) );
  NAND2_X1 U658 ( .A1(A[9]), .A2(B[9]), .ZN(n294) );
  INV_X1 U659 ( .A(n266), .ZN(n383) );
  NAND2_X1 U660 ( .A1(A[12]), .A2(B[12]), .ZN(n267) );
  NAND2_X1 U661 ( .A1(A[6]), .A2(B[6]), .ZN(n333) );
  NOR2_X1 U662 ( .A1(A[6]), .A2(B[6]), .ZN(n332) );
  INV_X1 U663 ( .A(n505), .ZN(n381) );
  NAND2_X1 U664 ( .A1(A[14]), .A2(B[14]), .ZN(n237) );
  NOR2_X1 U665 ( .A1(A[14]), .A2(B[14]), .ZN(n236) );
  INV_X1 U666 ( .A(n312), .ZN(n387) );
  NOR2_X2 U667 ( .A1(n319), .A2(n312), .ZN(n310) );
  NAND2_X1 U668 ( .A1(A[8]), .A2(B[8]), .ZN(n313) );
  INV_X1 U669 ( .A(n286), .ZN(n385) );
  NAND2_X1 U670 ( .A1(A[10]), .A2(B[10]), .ZN(n287) );
  NOR2_X1 U671 ( .A1(A[5]), .A2(B[5]), .ZN(n341) );
  INV_X4 U672 ( .A(n341), .ZN(n390) );
  XNOR2_X1 U673 ( .A(n39), .B(n5), .ZN(SUM[31]) );
  INV_X2 U674 ( .A(n86), .ZN(n84) );
  INV_X2 U675 ( .A(n77), .ZN(n75) );
  INV_X2 U676 ( .A(n73), .ZN(n71) );
  INV_X2 U677 ( .A(n64), .ZN(n62) );
  INV_X2 U678 ( .A(n49), .ZN(n47) );
  INV_X2 U679 ( .A(n362), .ZN(n395) );
  INV_X2 U680 ( .A(n360), .ZN(n394) );
  INV_X2 U681 ( .A(n356), .ZN(n393) );
  INV_X2 U682 ( .A(n353), .ZN(n392) );
  INV_X2 U683 ( .A(n94), .ZN(n369) );
  INV_X2 U684 ( .A(n85), .ZN(n83) );
  INV_X2 U685 ( .A(n72), .ZN(n70) );
  INV_X2 U686 ( .A(n63), .ZN(n61) );
  INV_X2 U687 ( .A(n48), .ZN(n46) );
  INV_X2 U688 ( .A(n37), .ZN(n364) );
  INV_X2 U689 ( .A(n359), .ZN(n358) );
  INV_X2 U690 ( .A(n345), .ZN(n347) );
  INV_X2 U691 ( .A(n4), .ZN(n391) );
  INV_X2 U692 ( .A(n342), .ZN(n340) );
  INV_X2 U693 ( .A(n333), .ZN(n331) );
  INV_X2 U694 ( .A(n332), .ZN(n389) );
  INV_X2 U695 ( .A(n325), .ZN(n323) );
  INV_X2 U696 ( .A(n324), .ZN(n322) );
  INV_X2 U697 ( .A(n299), .ZN(n297) );
  INV_X2 U698 ( .A(n298), .ZN(n296) );
  INV_X2 U699 ( .A(n279), .ZN(n277) );
  INV_X2 U700 ( .A(n278), .ZN(n276) );
  INV_X2 U701 ( .A(n262), .ZN(n260) );
  INV_X2 U702 ( .A(n249), .ZN(n247) );
  INV_X2 U703 ( .A(n248), .ZN(n246) );
  INV_X2 U704 ( .A(n229), .ZN(n227) );
  INV_X2 U705 ( .A(n228), .ZN(n226) );
  INV_X2 U706 ( .A(n224), .ZN(n222) );
  INV_X2 U707 ( .A(n223), .ZN(n380) );
  INV_X2 U708 ( .A(n209), .ZN(n207) );
  INV_X2 U709 ( .A(n208), .ZN(n206) );
  INV_X2 U710 ( .A(n205), .ZN(n203) );
  INV_X2 U711 ( .A(n204), .ZN(n202) );
  INV_X2 U712 ( .A(n200), .ZN(n198) );
  INV_X2 U713 ( .A(n185), .ZN(n183) );
  INV_X2 U714 ( .A(n184), .ZN(n182) );
  INV_X2 U715 ( .A(n180), .ZN(n178) );
  INV_X2 U716 ( .A(n167), .ZN(n165) );
  INV_X2 U717 ( .A(n156), .ZN(n154) );
  INV_X2 U718 ( .A(n155), .ZN(n374) );
  INV_X2 U719 ( .A(n131), .ZN(n372) );
  INV_X2 U720 ( .A(n126), .ZN(n124) );
  INV_X2 U721 ( .A(n125), .ZN(n123) );
  INV_X2 U722 ( .A(n121), .ZN(n119) );
  INV_X2 U723 ( .A(n120), .ZN(n371) );
  INV_X2 U724 ( .A(n112), .ZN(n110) );
  INV_X2 U725 ( .A(n111), .ZN(n370) );
  INV_X2 U726 ( .A(n36), .ZN(SUM[0]) );
endmodule


module up_island_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n299, n302, n305, n308, n311, n314, n317, n320, n323, n326, n329,
         n332, n335, n338, n341, n342, n347, n350, n353, n356, n359, n362,
         n365, n368, n371, n374, n377, n380, n383, n386, n389, n392, n395,
         n398, n401, n404, n407, n410, n413, n416, n419, n422, n425, n428,
         n431, n434, n437, n440, n441, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n574, n575, n576, n577, n578, n579, n581, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n594, n595, n596, n597, n598, n599,
         n601, n604, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n622, n623, n624, n625, n626,
         n627, n629, n632, n633, n634, n635, n636, n638, n639, n640, n641,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n657, n658, n659, n660, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n733, n734, n735, n736,
         n737, n738, n742, n743, n744, n745, n746, n747, n748, n749, n753,
         n754, n755, n756, n757, n758, n760, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n794, n795, n796, n797, n798, n799, n801, n804, n805,
         n806, n807, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n836, n837, n838, n839, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n859, n860, n861, n862, n863, n864, n865,
         n867, n868, n869, n870, n871, n872, n873, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297;
  assign n299 = b[1];
  assign n302 = b[3];
  assign n305 = b[5];
  assign n308 = b[7];
  assign n311 = b[9];
  assign n314 = b[11];
  assign n317 = b[13];
  assign n320 = b[15];
  assign n323 = b[17];
  assign n326 = b[19];
  assign n329 = b[21];
  assign n332 = b[23];
  assign n335 = b[25];
  assign n338 = b[27];
  assign n341 = b[29];
  assign n342 = b[31];
  assign n441 = a[0];
  assign n2929 = a[31];
  assign n2930 = a[30];
  assign n2931 = a[29];
  assign n2932 = a[28];
  assign n2933 = a[27];
  assign n2934 = a[26];
  assign n2935 = a[25];
  assign n2936 = a[24];
  assign n2937 = a[23];
  assign n2938 = a[22];
  assign n2939 = a[21];
  assign n2940 = a[20];
  assign n2941 = a[19];
  assign n2942 = a[18];
  assign n2943 = a[17];
  assign n2944 = a[16];
  assign n2945 = a[15];
  assign n2946 = a[14];
  assign n2947 = a[13];
  assign n2948 = a[12];
  assign n2949 = a[11];
  assign n2950 = a[10];
  assign n2951 = a[9];
  assign n2952 = a[8];
  assign n2953 = a[7];
  assign n2954 = a[6];
  assign n2955 = a[5];
  assign n2956 = a[4];
  assign n2957 = a[3];
  assign n2958 = a[2];
  assign n2959 = a[1];

  FA_X1 U239 ( .A(n1889), .B(n943), .CI(n505), .CO(n504), .S(product[62]) );
  FA_X1 U240 ( .A(n945), .B(n944), .CI(n506), .CO(n505), .S(product[61]) );
  XOR2_X2 U241 ( .A(n513), .B(n444), .Z(product[60]) );
  NAND2_X4 U243 ( .A1(n514), .A2(n883), .ZN(n507) );
  NAND2_X4 U247 ( .A1(n883), .A2(n512), .ZN(n444) );
  NOR2_X4 U249 ( .A1(n947), .A2(n946), .ZN(n511) );
  NAND2_X4 U250 ( .A1(n947), .A2(n946), .ZN(n512) );
  XOR2_X2 U251 ( .A(n518), .B(n445), .Z(product[59]) );
  NOR2_X4 U253 ( .A1(n521), .A2(n516), .ZN(n514) );
  NAND2_X4 U255 ( .A1(n884), .A2(n517), .ZN(n445) );
  NOR2_X4 U257 ( .A1(n948), .A2(n951), .ZN(n516) );
  NAND2_X4 U258 ( .A1(n948), .A2(n951), .ZN(n517) );
  NAND2_X4 U263 ( .A1(n612), .A2(n523), .ZN(n521) );
  NOR2_X4 U265 ( .A1(n544), .A2(n525), .ZN(n523) );
  NAND2_X4 U267 ( .A1(n534), .A2(n885), .ZN(n525) );
  AOI21_X4 U268 ( .B1(n535), .B2(n885), .A(n528), .ZN(n526) );
  NAND2_X4 U271 ( .A1(n885), .A2(n530), .ZN(n446) );
  NOR2_X4 U273 ( .A1(n952), .A2(n955), .ZN(n529) );
  NAND2_X4 U274 ( .A1(n952), .A2(n955), .ZN(n530) );
  XNOR2_X2 U275 ( .A(n538), .B(n447), .ZN(product[57]) );
  NOR2_X4 U279 ( .A1(n539), .A2(n536), .ZN(n534) );
  OAI21_X4 U280 ( .B1(n540), .B2(n536), .A(n537), .ZN(n535) );
  NAND2_X4 U281 ( .A1(n886), .A2(n537), .ZN(n447) );
  NOR2_X4 U283 ( .A1(n956), .A2(n961), .ZN(n536) );
  NAND2_X4 U284 ( .A1(n956), .A2(n961), .ZN(n537) );
  NAND2_X4 U287 ( .A1(n887), .A2(n540), .ZN(n448) );
  NOR2_X4 U289 ( .A1(n962), .A2(n967), .ZN(n539) );
  NAND2_X4 U290 ( .A1(n962), .A2(n967), .ZN(n540) );
  XNOR2_X2 U291 ( .A(n554), .B(n449), .ZN(product[55]) );
  NAND2_X4 U295 ( .A1(n589), .A2(n546), .ZN(n544) );
  AOI21_X4 U296 ( .B1(n590), .B2(n546), .A(n547), .ZN(n545) );
  NOR2_X4 U297 ( .A1(n548), .A2(n571), .ZN(n546) );
  OAI21_X4 U298 ( .B1(n548), .B2(n572), .A(n549), .ZN(n547) );
  NAND2_X4 U299 ( .A1(n558), .A2(n550), .ZN(n548) );
  AOI21_X4 U300 ( .B1(n559), .B2(n550), .A(n551), .ZN(n549) );
  NOR2_X4 U301 ( .A1(n555), .A2(n552), .ZN(n550) );
  OAI21_X4 U302 ( .B1(n552), .B2(n556), .A(n553), .ZN(n551) );
  NAND2_X4 U303 ( .A1(n888), .A2(n553), .ZN(n449) );
  NOR2_X4 U305 ( .A1(n968), .A2(n975), .ZN(n552) );
  NAND2_X4 U306 ( .A1(n968), .A2(n975), .ZN(n553) );
  XOR2_X2 U307 ( .A(n557), .B(n450), .Z(product[54]) );
  OAI21_X4 U308 ( .B1(n557), .B2(n555), .A(n556), .ZN(n554) );
  NAND2_X4 U309 ( .A1(n889), .A2(n556), .ZN(n450) );
  NOR2_X4 U317 ( .A1(n976), .A2(n983), .ZN(n555) );
  NAND2_X4 U318 ( .A1(n976), .A2(n983), .ZN(n556) );
  XNOR2_X2 U319 ( .A(n562), .B(n451), .ZN(product[53]) );
  AOI21_X4 U320 ( .B1(n566), .B2(n558), .A(n559), .ZN(n557) );
  NOR2_X4 U321 ( .A1(n563), .A2(n560), .ZN(n558) );
  OAI21_X4 U322 ( .B1(n560), .B2(n564), .A(n561), .ZN(n559) );
  NAND2_X4 U323 ( .A1(n890), .A2(n561), .ZN(n451) );
  NOR2_X4 U325 ( .A1(n984), .A2(n993), .ZN(n560) );
  NAND2_X4 U326 ( .A1(n984), .A2(n993), .ZN(n561) );
  XOR2_X2 U327 ( .A(n565), .B(n452), .Z(product[52]) );
  OAI21_X4 U328 ( .B1(n565), .B2(n563), .A(n564), .ZN(n562) );
  NAND2_X4 U329 ( .A1(n891), .A2(n564), .ZN(n452) );
  NOR2_X4 U331 ( .A1(n994), .A2(n1003), .ZN(n563) );
  NAND2_X4 U332 ( .A1(n994), .A2(n1003), .ZN(n564) );
  XNOR2_X2 U333 ( .A(n577), .B(n453), .ZN(product[51]) );
  NAND2_X4 U336 ( .A1(n585), .A2(n569), .ZN(n567) );
  AOI21_X4 U337 ( .B1(n586), .B2(n569), .A(n570), .ZN(n568) );
  NAND2_X4 U340 ( .A1(n893), .A2(n892), .ZN(n571) );
  AOI21_X4 U341 ( .B1(n892), .B2(n581), .A(n574), .ZN(n572) );
  NAND2_X4 U344 ( .A1(n892), .A2(n576), .ZN(n453) );
  NOR2_X4 U346 ( .A1(n1004), .A2(n1015), .ZN(n575) );
  NAND2_X4 U347 ( .A1(n1004), .A2(n1015), .ZN(n576) );
  XOR2_X2 U348 ( .A(n584), .B(n454), .Z(product[50]) );
  OAI21_X4 U349 ( .B1(n584), .B2(n578), .A(n579), .ZN(n577) );
  NAND2_X4 U354 ( .A1(n893), .A2(n579), .ZN(n454) );
  NOR2_X4 U356 ( .A1(n1016), .A2(n1027), .ZN(n578) );
  NAND2_X4 U357 ( .A1(n1016), .A2(n1027), .ZN(n579) );
  XNOR2_X2 U358 ( .A(n597), .B(n455), .ZN(product[49]) );
  NOR2_X4 U360 ( .A1(n610), .A2(n587), .ZN(n585) );
  OAI21_X4 U361 ( .B1(n611), .B2(n587), .A(n588), .ZN(n586) );
  NOR2_X4 U364 ( .A1(n607), .A2(n591), .ZN(n589) );
  OAI21_X4 U365 ( .B1(n591), .B2(n608), .A(n592), .ZN(n590) );
  NAND2_X4 U366 ( .A1(n894), .A2(n895), .ZN(n591) );
  AOI21_X4 U367 ( .B1(n894), .B2(n601), .A(n594), .ZN(n592) );
  NAND2_X4 U370 ( .A1(n894), .A2(n596), .ZN(n455) );
  NOR2_X4 U372 ( .A1(n1028), .A2(n1041), .ZN(n595) );
  NAND2_X4 U373 ( .A1(n1028), .A2(n1041), .ZN(n596) );
  XOR2_X2 U374 ( .A(n604), .B(n456), .Z(product[48]) );
  NAND2_X4 U380 ( .A1(n895), .A2(n599), .ZN(n456) );
  NAND2_X4 U388 ( .A1(n896), .A2(n608), .ZN(n457) );
  NOR2_X4 U390 ( .A1(n1056), .A2(n1071), .ZN(n607) );
  NAND2_X4 U391 ( .A1(n1056), .A2(n1071), .ZN(n608) );
  XOR2_X2 U392 ( .A(n620), .B(n458), .Z(product[46]) );
  NOR2_X4 U396 ( .A1(n614), .A2(n635), .ZN(n612) );
  OAI21_X4 U397 ( .B1(n614), .B2(n636), .A(n615), .ZN(n613) );
  NAND2_X4 U398 ( .A1(n616), .A2(n899), .ZN(n614) );
  AOI21_X4 U399 ( .B1(n616), .B2(n629), .A(n617), .ZN(n615) );
  NOR2_X4 U400 ( .A1(n623), .A2(n618), .ZN(n616) );
  OAI21_X4 U401 ( .B1(n618), .B2(n624), .A(n619), .ZN(n617) );
  NAND2_X4 U402 ( .A1(n897), .A2(n619), .ZN(n458) );
  NOR2_X4 U404 ( .A1(n1072), .A2(n1087), .ZN(n618) );
  NAND2_X4 U410 ( .A1(n898), .A2(n624), .ZN(n459) );
  NOR2_X4 U412 ( .A1(n1088), .A2(n1105), .ZN(n623) );
  NAND2_X4 U413 ( .A1(n1088), .A2(n1105), .ZN(n624) );
  NAND2_X4 U420 ( .A1(n899), .A2(n627), .ZN(n460) );
  NOR2_X4 U422 ( .A1(n1106), .A2(n1123), .ZN(n626) );
  NAND2_X4 U423 ( .A1(n1106), .A2(n1123), .ZN(n627) );
  XOR2_X2 U424 ( .A(n641), .B(n461), .Z(product[43]) );
  NAND2_X4 U428 ( .A1(n901), .A2(n900), .ZN(n635) );
  AOI21_X4 U429 ( .B1(n900), .B2(n643), .A(n638), .ZN(n636) );
  NAND2_X4 U432 ( .A1(n900), .A2(n640), .ZN(n461) );
  NOR2_X4 U434 ( .A1(n1124), .A2(n1143), .ZN(n639) );
  NAND2_X4 U435 ( .A1(n1124), .A2(n1143), .ZN(n640) );
  NAND2_X4 U440 ( .A1(n901), .A2(n645), .ZN(n462) );
  NOR2_X4 U442 ( .A1(n1144), .A2(n1163), .ZN(n644) );
  NAND2_X4 U443 ( .A1(n1144), .A2(n1163), .ZN(n645) );
  AOI21_X4 U446 ( .B1(n648), .B2(n700), .A(n649), .ZN(n647) );
  NOR2_X4 U447 ( .A1(n678), .A2(n650), .ZN(n648) );
  NAND2_X4 U457 ( .A1(n902), .A2(n659), .ZN(n463) );
  XNOR2_X2 U461 ( .A(n665), .B(n464), .ZN(product[40]) );
  NAND2_X4 U471 ( .A1(n904), .A2(n667), .ZN(n465) );
  XNOR2_X2 U475 ( .A(n673), .B(n466), .ZN(product[38]) );
  NAND2_X4 U479 ( .A1(n905), .A2(n672), .ZN(n466) );
  XOR2_X2 U483 ( .A(n676), .B(n467), .Z(product[37]) );
  OAI21_X4 U484 ( .B1(n676), .B2(n674), .A(n675), .ZN(n673) );
  NAND2_X4 U485 ( .A1(n906), .A2(n675), .ZN(n467) );
  NOR2_X4 U487 ( .A1(n1256), .A2(n1281), .ZN(n674) );
  XOR2_X2 U489 ( .A(n684), .B(n468), .Z(product[36]) );
  NAND2_X4 U496 ( .A1(n907), .A2(n683), .ZN(n468) );
  XNOR2_X2 U500 ( .A(n689), .B(n469), .ZN(product[35]) );
  AOI21_X4 U501 ( .B1(n689), .B2(n908), .A(n686), .ZN(n684) );
  NAND2_X4 U504 ( .A1(n908), .A2(n688), .ZN(n469) );
  XNOR2_X2 U508 ( .A(n696), .B(n470), .ZN(product[34]) );
  OAI21_X4 U509 ( .B1(n699), .B2(n690), .A(n691), .ZN(n689) );
  XOR2_X2 U518 ( .A(n699), .B(n471), .Z(product[33]) );
  XOR2_X2 U524 ( .A(n707), .B(n472), .Z(product[32]) );
  NAND2_X4 U527 ( .A1(n703), .A2(n717), .ZN(n701) );
  NOR2_X4 U529 ( .A1(n705), .A2(n714), .ZN(n703) );
  NAND2_X4 U531 ( .A1(n911), .A2(n706), .ZN(n472) );
  NAND2_X4 U539 ( .A1(n717), .A2(n912), .ZN(n710) );
  AOI21_X4 U540 ( .B1(n718), .B2(n912), .A(n713), .ZN(n711) );
  NAND2_X4 U543 ( .A1(n912), .A2(n715), .ZN(n473) );
  NOR2_X4 U545 ( .A1(n1424), .A2(n1453), .ZN(n714) );
  NAND2_X4 U546 ( .A1(n1424), .A2(n1453), .ZN(n715) );
  NOR2_X4 U549 ( .A1(n719), .A2(n724), .ZN(n717) );
  NAND2_X4 U551 ( .A1(n913), .A2(n720), .ZN(n474) );
  NAND2_X4 U559 ( .A1(n914), .A2(n725), .ZN(n475) );
  NAND2_X4 U562 ( .A1(n1482), .A2(n1509), .ZN(n725) );
  XNOR2_X2 U563 ( .A(n736), .B(n476), .ZN(product[28]) );
  OAI21_X4 U577 ( .B1(n763), .B2(n737), .A(n738), .ZN(n736) );
  XNOR2_X2 U612 ( .A(n771), .B(n480), .ZN(product[24]) );
  NAND2_X4 U619 ( .A1(n919), .A2(n770), .ZN(n480) );
  XOR2_X2 U623 ( .A(n774), .B(n481), .Z(product[23]) );
  OAI21_X4 U624 ( .B1(n774), .B2(n772), .A(n773), .ZN(n771) );
  NAND2_X4 U625 ( .A1(n920), .A2(n773), .ZN(n481) );
  NOR2_X4 U627 ( .A1(n1632), .A2(n1653), .ZN(n772) );
  XOR2_X2 U629 ( .A(n779), .B(n482), .Z(product[22]) );
  AOI21_X4 U630 ( .B1(n784), .B2(n775), .A(n776), .ZN(n774) );
  NOR2_X4 U631 ( .A1(n782), .A2(n777), .ZN(n775) );
  OAI21_X4 U632 ( .B1(n777), .B2(n783), .A(n778), .ZN(n776) );
  NAND2_X4 U633 ( .A1(n921), .A2(n778), .ZN(n482) );
  NOR2_X4 U635 ( .A1(n1654), .A2(n1673), .ZN(n777) );
  NAND2_X4 U636 ( .A1(n1654), .A2(n1673), .ZN(n778) );
  NAND2_X4 U641 ( .A1(n922), .A2(n783), .ZN(n483) );
  NOR2_X4 U643 ( .A1(n1674), .A2(n1693), .ZN(n782) );
  NAND2_X4 U644 ( .A1(n1674), .A2(n1693), .ZN(n783) );
  XNOR2_X2 U645 ( .A(n790), .B(n484), .ZN(product[20]) );
  NOR2_X4 U648 ( .A1(n791), .A2(n788), .ZN(n786) );
  NAND2_X4 U650 ( .A1(n923), .A2(n789), .ZN(n484) );
  NOR2_X4 U652 ( .A1(n1694), .A2(n1711), .ZN(n788) );
  NAND2_X4 U653 ( .A1(n1694), .A2(n1711), .ZN(n789) );
  XNOR2_X2 U654 ( .A(n797), .B(n485), .ZN(product[19]) );
  NAND2_X4 U656 ( .A1(n924), .A2(n925), .ZN(n791) );
  XOR2_X2 U664 ( .A(n804), .B(n486), .Z(product[18]) );
  OAI21_X4 U665 ( .B1(n804), .B2(n798), .A(n799), .ZN(n797) );
  NAND2_X4 U670 ( .A1(n925), .A2(n799), .ZN(n486) );
  NOR2_X4 U672 ( .A1(n1730), .A2(n1745), .ZN(n798) );
  NAND2_X4 U673 ( .A1(n1730), .A2(n1745), .ZN(n799) );
  XOR2_X2 U674 ( .A(n812), .B(n487), .Z(product[17]) );
  NAND2_X4 U677 ( .A1(n813), .A2(n926), .ZN(n806) );
  AOI21_X4 U678 ( .B1(n814), .B2(n926), .A(n809), .ZN(n807) );
  NAND2_X4 U681 ( .A1(n926), .A2(n811), .ZN(n487) );
  XOR2_X2 U685 ( .A(n817), .B(n488), .Z(product[16]) );
  AOI21_X4 U686 ( .B1(n822), .B2(n813), .A(n814), .ZN(n812) );
  NOR2_X4 U687 ( .A1(n815), .A2(n820), .ZN(n813) );
  OAI21_X4 U688 ( .B1(n815), .B2(n821), .A(n816), .ZN(n814) );
  NAND2_X4 U689 ( .A1(n927), .A2(n816), .ZN(n488) );
  NOR2_X4 U691 ( .A1(n1762), .A2(n1775), .ZN(n815) );
  XNOR2_X2 U693 ( .A(n822), .B(n489), .ZN(product[15]) );
  AOI21_X4 U694 ( .B1(n822), .B2(n928), .A(n819), .ZN(n817) );
  NAND2_X4 U697 ( .A1(n928), .A2(n821), .ZN(n489) );
  NOR2_X4 U699 ( .A1(n1776), .A2(n1789), .ZN(n820) );
  NAND2_X4 U700 ( .A1(n1776), .A2(n1789), .ZN(n821) );
  XNOR2_X2 U701 ( .A(n828), .B(n490), .ZN(product[14]) );
  AOI21_X4 U703 ( .B1(n832), .B2(n824), .A(n825), .ZN(n823) );
  NOR2_X4 U704 ( .A1(n826), .A2(n829), .ZN(n824) );
  OAI21_X4 U705 ( .B1(n826), .B2(n830), .A(n827), .ZN(n825) );
  NAND2_X4 U706 ( .A1(n929), .A2(n827), .ZN(n490) );
  NOR2_X4 U708 ( .A1(n1790), .A2(n1801), .ZN(n826) );
  NAND2_X4 U709 ( .A1(n1790), .A2(n1801), .ZN(n827) );
  XOR2_X2 U710 ( .A(n831), .B(n491), .Z(product[13]) );
  OAI21_X4 U711 ( .B1(n831), .B2(n829), .A(n830), .ZN(n828) );
  NAND2_X4 U712 ( .A1(n930), .A2(n830), .ZN(n491) );
  NOR2_X4 U714 ( .A1(n1802), .A2(n1813), .ZN(n829) );
  NAND2_X4 U715 ( .A1(n1802), .A2(n1813), .ZN(n830) );
  XOR2_X2 U716 ( .A(n839), .B(n492), .Z(product[12]) );
  OAI21_X4 U718 ( .B1(n845), .B2(n833), .A(n834), .ZN(n832) );
  NAND2_X4 U719 ( .A1(n932), .A2(n931), .ZN(n833) );
  AOI21_X4 U720 ( .B1(n931), .B2(n841), .A(n836), .ZN(n834) );
  NAND2_X4 U723 ( .A1(n931), .A2(n838), .ZN(n492) );
  XNOR2_X2 U727 ( .A(n844), .B(n493), .ZN(product[11]) );
  AOI21_X4 U728 ( .B1(n844), .B2(n932), .A(n841), .ZN(n839) );
  NAND2_X4 U731 ( .A1(n932), .A2(n843), .ZN(n493) );
  NOR2_X4 U733 ( .A1(n1824), .A2(n1833), .ZN(n842) );
  NAND2_X4 U734 ( .A1(n1824), .A2(n1833), .ZN(n843) );
  XNOR2_X2 U735 ( .A(n850), .B(n494), .ZN(product[10]) );
  AOI21_X4 U737 ( .B1(n846), .B2(n854), .A(n847), .ZN(n845) );
  NOR2_X4 U738 ( .A1(n848), .A2(n851), .ZN(n846) );
  OAI21_X4 U739 ( .B1(n848), .B2(n852), .A(n849), .ZN(n847) );
  NAND2_X4 U740 ( .A1(n933), .A2(n849), .ZN(n494) );
  NOR2_X4 U742 ( .A1(n1834), .A2(n1841), .ZN(n848) );
  NAND2_X4 U743 ( .A1(n1834), .A2(n1841), .ZN(n849) );
  XOR2_X2 U744 ( .A(n853), .B(n495), .Z(product[9]) );
  OAI21_X4 U745 ( .B1(n853), .B2(n851), .A(n852), .ZN(n850) );
  NAND2_X4 U746 ( .A1(n934), .A2(n852), .ZN(n495) );
  NOR2_X4 U748 ( .A1(n1842), .A2(n1849), .ZN(n851) );
  NAND2_X4 U749 ( .A1(n1842), .A2(n1849), .ZN(n852) );
  XOR2_X2 U750 ( .A(n857), .B(n496), .Z(product[8]) );
  OAI21_X4 U752 ( .B1(n857), .B2(n855), .A(n856), .ZN(n854) );
  NAND2_X4 U753 ( .A1(n935), .A2(n856), .ZN(n496) );
  NOR2_X4 U755 ( .A1(n1850), .A2(n1855), .ZN(n855) );
  NAND2_X4 U756 ( .A1(n1850), .A2(n1855), .ZN(n856) );
  XNOR2_X2 U757 ( .A(n497), .B(n862), .ZN(product[7]) );
  AOI21_X4 U758 ( .B1(n862), .B2(n936), .A(n859), .ZN(n857) );
  NAND2_X4 U761 ( .A1(n936), .A2(n861), .ZN(n497) );
  NOR2_X4 U763 ( .A1(n1856), .A2(n1861), .ZN(n860) );
  NAND2_X4 U764 ( .A1(n1856), .A2(n1861), .ZN(n861) );
  XOR2_X2 U765 ( .A(n498), .B(n865), .Z(product[6]) );
  OAI21_X4 U766 ( .B1(n863), .B2(n865), .A(n864), .ZN(n862) );
  NAND2_X4 U767 ( .A1(n937), .A2(n864), .ZN(n498) );
  NOR2_X4 U769 ( .A1(n1862), .A2(n1865), .ZN(n863) );
  NAND2_X4 U770 ( .A1(n1862), .A2(n1865), .ZN(n864) );
  XNOR2_X2 U771 ( .A(n499), .B(n870), .ZN(product[5]) );
  AOI21_X4 U772 ( .B1(n938), .B2(n870), .A(n867), .ZN(n865) );
  NAND2_X4 U775 ( .A1(n938), .A2(n869), .ZN(n499) );
  NOR2_X4 U777 ( .A1(n1866), .A2(n1869), .ZN(n868) );
  NAND2_X4 U778 ( .A1(n1866), .A2(n1869), .ZN(n869) );
  XOR2_X2 U779 ( .A(n500), .B(n873), .Z(product[4]) );
  OAI21_X4 U780 ( .B1(n873), .B2(n871), .A(n872), .ZN(n870) );
  NAND2_X4 U781 ( .A1(n939), .A2(n872), .ZN(n500) );
  NOR2_X4 U783 ( .A1(n1870), .A2(n2366), .ZN(n871) );
  NAND2_X4 U784 ( .A1(n1870), .A2(n2366), .ZN(n872) );
  XNOR2_X2 U785 ( .A(n878), .B(n501), .ZN(product[3]) );
  AOI21_X4 U786 ( .B1(n878), .B2(n940), .A(n875), .ZN(n873) );
  NAND2_X4 U789 ( .A1(n940), .A2(n877), .ZN(n501) );
  NOR2_X4 U791 ( .A1(n2398), .A2(n1872), .ZN(n876) );
  NAND2_X4 U792 ( .A1(n2398), .A2(n1872), .ZN(n877) );
  XOR2_X2 U793 ( .A(n502), .B(n882), .Z(product[2]) );
  OAI21_X4 U794 ( .B1(n879), .B2(n882), .A(n880), .ZN(n878) );
  NAND2_X4 U795 ( .A1(n941), .A2(n880), .ZN(n502) );
  NOR2_X4 U797 ( .A1(n2399), .A2(n2368), .ZN(n879) );
  NAND2_X4 U798 ( .A1(n2399), .A2(n2368), .ZN(n880) );
  NAND2_X4 U800 ( .A1(n942), .A2(n882), .ZN(n503) );
  NOR2_X4 U802 ( .A1(n2400), .A2(n1888), .ZN(n881) );
  NAND2_X4 U803 ( .A1(n2400), .A2(n1888), .ZN(n882) );
  FA_X1 U805 ( .A(n1890), .B(n949), .CI(n1921), .CO(n945), .S(n946) );
  FA_X1 U806 ( .A(n1891), .B(n950), .CI(n953), .CO(n947), .S(n948) );
  FA_X1 U808 ( .A(n957), .B(n1948), .CI(n954), .CO(n951), .S(n952) );
  FA_X1 U809 ( .A(n1922), .B(n959), .CI(n1892), .CO(n953), .S(n954) );
  FA_X1 U810 ( .A(n958), .B(n965), .CI(n963), .CO(n955), .S(n956) );
  FA_X1 U811 ( .A(n1949), .B(n960), .CI(n1893), .CO(n957), .S(n958) );
  FA_X1 U813 ( .A(n969), .B(n966), .CI(n964), .CO(n961), .S(n962) );
  FA_X1 U814 ( .A(n1979), .B(n1894), .CI(n971), .CO(n963), .S(n964) );
  FA_X1 U815 ( .A(n973), .B(n1923), .CI(n1950), .CO(n965), .S(n966) );
  FA_X1 U816 ( .A(n977), .B(n972), .CI(n970), .CO(n967), .S(n968) );
  FA_X1 U817 ( .A(n981), .B(n1895), .CI(n979), .CO(n969), .S(n970) );
  FA_X1 U818 ( .A(n974), .B(n1924), .CI(n1980), .CO(n971), .S(n972) );
  FA_X1 U820 ( .A(n985), .B(n980), .CI(n978), .CO(n975), .S(n976) );
  FA_X1 U821 ( .A(n982), .B(n989), .CI(n987), .CO(n977), .S(n978) );
  FA_X1 U822 ( .A(n1896), .B(n1925), .CI(n2010), .CO(n979), .S(n980) );
  FA_X1 U823 ( .A(n1951), .B(n991), .CI(n1981), .CO(n981), .S(n982) );
  FA_X1 U824 ( .A(n995), .B(n988), .CI(n986), .CO(n983), .S(n984) );
  FA_X1 U825 ( .A(n999), .B(n990), .CI(n997), .CO(n985), .S(n986) );
  FA_X1 U826 ( .A(n1897), .B(n2011), .CI(n1001), .CO(n987), .S(n988) );
  FA_X1 U827 ( .A(n1982), .B(n992), .CI(n1952), .CO(n989), .S(n990) );
  FA_X1 U829 ( .A(n1005), .B(n998), .CI(n996), .CO(n993), .S(n994) );
  FA_X1 U830 ( .A(n1000), .B(n1009), .CI(n1007), .CO(n995), .S(n996) );
  FA_X1 U831 ( .A(n1011), .B(n2043), .CI(n1002), .CO(n997), .S(n998) );
  FA_X1 U832 ( .A(n2012), .B(n1926), .CI(n1898), .CO(n999), .S(n1000) );
  FA_X1 U833 ( .A(n1983), .B(n1013), .CI(n1953), .CO(n1001), .S(n1002) );
  FA_X1 U834 ( .A(n1017), .B(n1008), .CI(n1006), .CO(n1003), .S(n1004) );
  FA_X1 U835 ( .A(n1010), .B(n1021), .CI(n1019), .CO(n1005), .S(n1006) );
  FA_X1 U836 ( .A(n1023), .B(n1899), .CI(n1012), .CO(n1007), .S(n1008) );
  FA_X1 U837 ( .A(n1025), .B(n2013), .CI(n2044), .CO(n1009), .S(n1010) );
  FA_X1 U838 ( .A(n1984), .B(n1014), .CI(n1927), .CO(n1011), .S(n1012) );
  FA_X1 U840 ( .A(n1029), .B(n1020), .CI(n1018), .CO(n1015), .S(n1016) );
  FA_X1 U841 ( .A(n1022), .B(n1033), .CI(n1031), .CO(n1017), .S(n1018) );
  FA_X1 U842 ( .A(n1035), .B(n1037), .CI(n1024), .CO(n1019), .S(n1020) );
  FA_X1 U843 ( .A(n2073), .B(n1900), .CI(n1026), .CO(n1021), .S(n1022) );
  FA_X1 U844 ( .A(n2045), .B(n1954), .CI(n1985), .CO(n1023), .S(n1024) );
  FA_X1 U845 ( .A(n1039), .B(n1928), .CI(n2014), .CO(n1025), .S(n1026) );
  FA_X1 U846 ( .A(n1043), .B(n1032), .CI(n1030), .CO(n1027), .S(n1028) );
  FA_X1 U847 ( .A(n1034), .B(n1047), .CI(n1045), .CO(n1029), .S(n1030) );
  FA_X1 U848 ( .A(n1049), .B(n1038), .CI(n1036), .CO(n1031), .S(n1032) );
  FA_X1 U849 ( .A(n1901), .B(n2074), .CI(n1051), .CO(n1033), .S(n1034) );
  FA_X1 U850 ( .A(n1929), .B(n2046), .CI(n1053), .CO(n1035), .S(n1036) );
  FA_X1 U851 ( .A(n2015), .B(n1040), .CI(n1955), .CO(n1037), .S(n1038) );
  FA_X1 U853 ( .A(n1057), .B(n1046), .CI(n1044), .CO(n1041), .S(n1042) );
  FA_X1 U854 ( .A(n1048), .B(n1061), .CI(n1059), .CO(n1043), .S(n1044) );
  FA_X1 U855 ( .A(n1052), .B(n1063), .CI(n1050), .CO(n1045), .S(n1046) );
  FA_X1 U856 ( .A(n1067), .B(n1054), .CI(n1065), .CO(n1047), .S(n1048) );
  FA_X1 U857 ( .A(n1902), .B(n2075), .CI(n2106), .CO(n1049), .S(n1050) );
  FA_X1 U858 ( .A(n2016), .B(n1986), .CI(n1930), .CO(n1051), .S(n1052) );
  FA_X1 U859 ( .A(n1956), .B(n2047), .CI(n1069), .CO(n1053), .S(n1054) );
  FA_X1 U860 ( .A(n1073), .B(n1060), .CI(n1058), .CO(n1055), .S(n1056) );
  FA_X1 U861 ( .A(n1062), .B(n1077), .CI(n1075), .CO(n1057), .S(n1058) );
  FA_X1 U862 ( .A(n1079), .B(n1066), .CI(n1064), .CO(n1059), .S(n1060) );
  FA_X1 U863 ( .A(n1068), .B(n1083), .CI(n1081), .CO(n1061), .S(n1062) );
  FA_X1 U864 ( .A(n2107), .B(n1085), .CI(n1903), .CO(n1063), .S(n1064) );
  FA_X1 U865 ( .A(n2048), .B(n1957), .CI(n2076), .CO(n1065), .S(n1066) );
  FA_X1 U866 ( .A(n1070), .B(n2017), .CI(n1987), .CO(n1067), .S(n1068) );
  FA_X1 U868 ( .A(n1089), .B(n1076), .CI(n1074), .CO(n1071), .S(n1072) );
  FA_X1 U869 ( .A(n1078), .B(n1093), .CI(n1091), .CO(n1073), .S(n1074) );
  FA_X1 U870 ( .A(n1095), .B(n1082), .CI(n1080), .CO(n1075), .S(n1076) );
  FA_X1 U871 ( .A(n1097), .B(n1099), .CI(n1084), .CO(n1077), .S(n1078) );
  FA_X1 U872 ( .A(n1086), .B(n2139), .CI(n1101), .CO(n1079), .S(n1080) );
  FA_X1 U873 ( .A(n2018), .B(n2108), .CI(n1904), .CO(n1081), .S(n1082) );
  FA_X1 U874 ( .A(n1931), .B(n1958), .CI(n2049), .CO(n1083), .S(n1084) );
  FA_X1 U875 ( .A(n1988), .B(n1103), .CI(n2077), .CO(n1085), .S(n1086) );
  FA_X1 U876 ( .A(n1107), .B(n1092), .CI(n1090), .CO(n1087), .S(n1088) );
  FA_X1 U877 ( .A(n1094), .B(n1111), .CI(n1109), .CO(n1089), .S(n1090) );
  FA_X1 U878 ( .A(n1113), .B(n1098), .CI(n1096), .CO(n1091), .S(n1092) );
  FA_X1 U879 ( .A(n1100), .B(n1102), .CI(n1115), .CO(n1093), .S(n1094) );
  FA_X1 U880 ( .A(n1119), .B(n1905), .CI(n1117), .CO(n1095), .S(n1096) );
  FA_X1 U881 ( .A(n1121), .B(n2109), .CI(n2140), .CO(n1097), .S(n1098) );
  FA_X1 U882 ( .A(n2078), .B(n1989), .CI(n1932), .CO(n1099), .S(n1100) );
  FA_X1 U883 ( .A(n1104), .B(n1959), .CI(n2019), .CO(n1101), .S(n1102) );
  FA_X1 U885 ( .A(n1125), .B(n1110), .CI(n1108), .CO(n1105), .S(n1106) );
  FA_X1 U886 ( .A(n1112), .B(n1129), .CI(n1127), .CO(n1107), .S(n1108) );
  FA_X1 U887 ( .A(n1131), .B(n1116), .CI(n1114), .CO(n1109), .S(n1110) );
  FA_X1 U888 ( .A(n1118), .B(n1120), .CI(n1133), .CO(n1111), .S(n1112) );
  FA_X1 U889 ( .A(n1137), .B(n1139), .CI(n1135), .CO(n1113), .S(n1114) );
  FA_X1 U890 ( .A(n2172), .B(n1906), .CI(n1122), .CO(n1115), .S(n1116) );
  FA_X1 U891 ( .A(n2050), .B(n2141), .CI(n2079), .CO(n1117), .S(n1118) );
  FA_X1 U892 ( .A(n1990), .B(n2110), .CI(n1960), .CO(n1119), .S(n1120) );
  FA_X1 U893 ( .A(n1141), .B(n1933), .CI(n2020), .CO(n1121), .S(n1122) );
  FA_X1 U894 ( .A(n1145), .B(n1128), .CI(n1126), .CO(n1123), .S(n1124) );
  FA_X1 U895 ( .A(n1130), .B(n1149), .CI(n1147), .CO(n1125), .S(n1126) );
  FA_X1 U896 ( .A(n1151), .B(n1134), .CI(n1132), .CO(n1127), .S(n1128) );
  FA_X1 U897 ( .A(n1136), .B(n1138), .CI(n1153), .CO(n1129), .S(n1130) );
  FA_X1 U898 ( .A(n1140), .B(n1157), .CI(n1155), .CO(n1131), .S(n1132) );
  FA_X1 U899 ( .A(n1907), .B(n2173), .CI(n1159), .CO(n1133), .S(n1134) );
  FA_X1 U900 ( .A(n2111), .B(n2142), .CI(n1161), .CO(n1135), .S(n1136) );
  FA_X1 U901 ( .A(n1934), .B(n1961), .CI(n2051), .CO(n1137), .S(n1138) );
  FA_X1 U902 ( .A(n1142), .B(n2080), .CI(n2021), .CO(n1139), .S(n1140) );
  FA_X1 U904 ( .A(n1165), .B(n1148), .CI(n1146), .CO(n1143), .S(n1144) );
  FA_X1 U905 ( .A(n1150), .B(n1169), .CI(n1167), .CO(n1145), .S(n1146) );
  FA_X1 U906 ( .A(n1171), .B(n1154), .CI(n1152), .CO(n1147), .S(n1148) );
  FA_X1 U907 ( .A(n1156), .B(n1158), .CI(n1173), .CO(n1149), .S(n1150) );
  FA_X1 U908 ( .A(n1160), .B(n1177), .CI(n1175), .CO(n1151), .S(n1152) );
  FA_X1 U909 ( .A(n1162), .B(n2204), .CI(n1179), .CO(n1153), .S(n1154) );
  FA_X1 U910 ( .A(n1181), .B(n2174), .CI(n1908), .CO(n1155), .S(n1156) );
  FA_X1 U911 ( .A(n1935), .B(n2112), .CI(n2081), .CO(n1157), .S(n1158) );
  FA_X1 U912 ( .A(n2022), .B(n1183), .CI(n1991), .CO(n1159), .S(n1160) );
  FA_X1 U913 ( .A(n1962), .B(n2052), .CI(n2143), .CO(n1161), .S(n1162) );
  FA_X1 U914 ( .A(n1187), .B(n1168), .CI(n1166), .CO(n1163), .S(n1164) );
  FA_X1 U915 ( .A(n1170), .B(n1191), .CI(n1189), .CO(n1165), .S(n1166) );
  FA_X1 U916 ( .A(n1193), .B(n1174), .CI(n1172), .CO(n1167), .S(n1168) );
  FA_X1 U917 ( .A(n1176), .B(n1197), .CI(n1195), .CO(n1169), .S(n1170) );
  FA_X1 U918 ( .A(n1178), .B(n1199), .CI(n1180), .CO(n1171), .S(n1172) );
  FA_X1 U919 ( .A(n1203), .B(n1182), .CI(n1201), .CO(n1173), .S(n1174) );
  FA_X1 U920 ( .A(n2205), .B(n1205), .CI(n1909), .CO(n1175), .S(n1176) );
  FA_X1 U921 ( .A(n2053), .B(n2144), .CI(n2175), .CO(n1177), .S(n1178) );
  FA_X1 U922 ( .A(n1963), .B(n1992), .CI(n2082), .CO(n1179), .S(n1180) );
  FA_X1 U923 ( .A(n2023), .B(n2113), .CI(n1184), .CO(n1181), .S(n1182) );
  FA_X1 U925 ( .A(n1209), .B(n1190), .CI(n1188), .CO(n1185), .S(n1186) );
  FA_X1 U926 ( .A(n1192), .B(n1213), .CI(n1211), .CO(n1187), .S(n1188) );
  FA_X1 U927 ( .A(n1196), .B(n1215), .CI(n1194), .CO(n1189), .S(n1190) );
  FA_X1 U928 ( .A(n1198), .B(n1219), .CI(n1217), .CO(n1191), .S(n1192) );
  FA_X1 U929 ( .A(n1202), .B(n1204), .CI(n1200), .CO(n1193), .S(n1194) );
  FA_X1 U930 ( .A(n1223), .B(n1225), .CI(n1221), .CO(n1195), .S(n1196) );
  FA_X1 U931 ( .A(n2237), .B(n1910), .CI(n1206), .CO(n1197), .S(n1198) );
  FA_X1 U932 ( .A(n2145), .B(n2206), .CI(n1227), .CO(n1199), .S(n1200) );
  FA_X1 U933 ( .A(n2114), .B(n1936), .CI(n1964), .CO(n1201), .S(n1202) );
  FA_X1 U934 ( .A(n2024), .B(n1229), .CI(n2054), .CO(n1203), .S(n1204) );
  FA_X1 U935 ( .A(n1993), .B(n2176), .CI(n2083), .CO(n1205), .S(n1206) );
  FA_X1 U936 ( .A(n1233), .B(n1212), .CI(n1210), .CO(n1207), .S(n1208) );
  FA_X1 U937 ( .A(n1214), .B(n1237), .CI(n1235), .CO(n1209), .S(n1210) );
  FA_X1 U938 ( .A(n1239), .B(n1218), .CI(n1216), .CO(n1211), .S(n1212) );
  FA_X1 U939 ( .A(n1220), .B(n1243), .CI(n1241), .CO(n1213), .S(n1214) );
  FA_X1 U940 ( .A(n1245), .B(n1226), .CI(n1222), .CO(n1215), .S(n1216) );
  FA_X1 U941 ( .A(n1247), .B(n1249), .CI(n1224), .CO(n1217), .S(n1218) );
  FA_X1 U942 ( .A(n1228), .B(n1911), .CI(n1251), .CO(n1219), .S(n1220) );
  FA_X1 U943 ( .A(n1253), .B(n2115), .CI(n2238), .CO(n1221), .S(n1222) );
  FA_X1 U944 ( .A(n2084), .B(n2177), .CI(n2207), .CO(n1223), .S(n1224) );
  FA_X1 U945 ( .A(n1937), .B(n2025), .CI(n1994), .CO(n1225), .S(n1226) );
  FA_X1 U946 ( .A(n2146), .B(n1965), .CI(n1230), .CO(n1227), .S(n1228) );
  FA_X1 U948 ( .A(n1257), .B(n1236), .CI(n1234), .CO(n1231), .S(n1232) );
  FA_X1 U949 ( .A(n1238), .B(n1261), .CI(n1259), .CO(n1233), .S(n1234) );
  FA_X1 U950 ( .A(n1263), .B(n1242), .CI(n1240), .CO(n1235), .S(n1236) );
  FA_X1 U951 ( .A(n1244), .B(n1267), .CI(n1265), .CO(n1237), .S(n1238) );
  FA_X1 U952 ( .A(n1269), .B(n1250), .CI(n1246), .CO(n1239), .S(n1240) );
  FA_X1 U953 ( .A(n1252), .B(n1271), .CI(n1248), .CO(n1241), .S(n1242) );
  FA_X1 U954 ( .A(n1275), .B(n1254), .CI(n1273), .CO(n1243), .S(n1244) );
  FA_X1 U955 ( .A(n1912), .B(n1277), .CI(n2270), .CO(n1245), .S(n1246) );
  FA_X1 U956 ( .A(n1966), .B(n2178), .CI(n2239), .CO(n1247), .S(n1248) );
  FA_X1 U957 ( .A(n2085), .B(n1995), .CI(n2147), .CO(n1249), .S(n1250) );
  FA_X1 U958 ( .A(n2116), .B(n1938), .CI(n2055), .CO(n1251), .S(n1252) );
  FA_X1 U959 ( .A(n2208), .B(n1279), .CI(n2026), .CO(n1253), .S(n1254) );
  FA_X1 U960 ( .A(n1283), .B(n1260), .CI(n1258), .CO(n1255), .S(n1256) );
  FA_X1 U962 ( .A(n1289), .B(n1266), .CI(n1264), .CO(n1259), .S(n1260) );
  FA_X1 U963 ( .A(n1268), .B(n1293), .CI(n1291), .CO(n1261), .S(n1262) );
  FA_X1 U964 ( .A(n1295), .B(n1272), .CI(n1270), .CO(n1263), .S(n1264) );
  FA_X1 U965 ( .A(n1274), .B(n1297), .CI(n1276), .CO(n1265), .S(n1266) );
  FA_X1 U966 ( .A(n1301), .B(n1303), .CI(n1299), .CO(n1267), .S(n1268) );
  FA_X1 U967 ( .A(n1913), .B(n2271), .CI(n1278), .CO(n1269), .S(n1270) );
  FA_X1 U968 ( .A(n2240), .B(n2209), .CI(n1305), .CO(n1271), .S(n1272) );
  FA_X1 U969 ( .A(n2148), .B(n2027), .CI(n2117), .CO(n1273), .S(n1274) );
  FA_X1 U970 ( .A(n1967), .B(n2056), .CI(n1939), .CO(n1275), .S(n1276) );
  FA_X1 U971 ( .A(n2086), .B(n1996), .CI(n1280), .CO(n1277), .S(n1278) );
  FA_X1 U973 ( .A(n1309), .B(n1286), .CI(n1284), .CO(n1281), .S(n1282) );
  FA_X1 U974 ( .A(n1288), .B(n1313), .CI(n1311), .CO(n1283), .S(n1284) );
  FA_X1 U975 ( .A(n1315), .B(n1292), .CI(n1290), .CO(n1285), .S(n1286) );
  FA_X1 U976 ( .A(n1317), .B(n1296), .CI(n1294), .CO(n1287), .S(n1288) );
  FA_X1 U977 ( .A(n1321), .B(n1298), .CI(n1319), .CO(n1289), .S(n1290) );
  FA_X1 U978 ( .A(n1300), .B(n1323), .CI(n1302), .CO(n1291), .S(n1292) );
  FA_X1 U979 ( .A(n1325), .B(n1327), .CI(n1304), .CO(n1293), .S(n1294) );
  FA_X1 U980 ( .A(n1306), .B(n2303), .CI(n1329), .CO(n1295), .S(n1296) );
  FA_X1 U981 ( .A(n1331), .B(n2179), .CI(n1914), .CO(n1297), .S(n1298) );
  FA_X1 U982 ( .A(n1997), .B(n2210), .CI(n2272), .CO(n1299), .S(n1300) );
  FA_X1 U983 ( .A(n1940), .B(n2028), .CI(n2118), .CO(n1301), .S(n1302) );
  FA_X1 U984 ( .A(n1333), .B(n1968), .CI(n2087), .CO(n1303), .S(n1304) );
  FA_X1 U985 ( .A(n2149), .B(n2057), .CI(n2241), .CO(n1305), .S(n1306) );
  FA_X1 U986 ( .A(n1337), .B(n1312), .CI(n1310), .CO(n1307), .S(n1308) );
  FA_X1 U987 ( .A(n1314), .B(n1316), .CI(n1339), .CO(n1309), .S(n1310) );
  FA_X1 U988 ( .A(n1343), .B(n1318), .CI(n1341), .CO(n1311), .S(n1312) );
  FA_X1 U989 ( .A(n1345), .B(n1322), .CI(n1320), .CO(n1313), .S(n1314) );
  FA_X1 U990 ( .A(n1349), .B(n1324), .CI(n1347), .CO(n1315), .S(n1316) );
  FA_X1 U991 ( .A(n1328), .B(n1326), .CI(n1351), .CO(n1317), .S(n1318) );
  FA_X1 U992 ( .A(n1353), .B(n1355), .CI(n1330), .CO(n1319), .S(n1320) );
  FA_X1 U993 ( .A(n1359), .B(n1332), .CI(n1357), .CO(n1321), .S(n1322) );
  FA_X1 U994 ( .A(n2304), .B(n1361), .CI(n1915), .CO(n1323), .S(n1324) );
  FA_X1 U995 ( .A(n2273), .B(n2242), .CI(n1969), .CO(n1325), .S(n1326) );
  FA_X1 U996 ( .A(n2150), .B(n1998), .CI(n2180), .CO(n1327), .S(n1328) );
  FA_X1 U997 ( .A(n2088), .B(n2211), .CI(n2058), .CO(n1329), .S(n1330) );
  FA_X1 U998 ( .A(n2029), .B(n2119), .CI(n1334), .CO(n1331), .S(n1332) );
  FA_X1 U1000 ( .A(n1365), .B(n1340), .CI(n1338), .CO(n1335), .S(n1336) );
  FA_X1 U1001 ( .A(n1342), .B(n1369), .CI(n1367), .CO(n1337), .S(n1338) );
  FA_X1 U1002 ( .A(n1371), .B(n1346), .CI(n1344), .CO(n1339), .S(n1340) );
  FA_X1 U1003 ( .A(n1373), .B(n1375), .CI(n1348), .CO(n1341), .S(n1342) );
  FA_X1 U1004 ( .A(n1352), .B(n1377), .CI(n1350), .CO(n1343), .S(n1344) );
  FA_X1 U1005 ( .A(n1379), .B(n1356), .CI(n1354), .CO(n1345), .S(n1346) );
  FA_X1 U1006 ( .A(n1360), .B(n1381), .CI(n1358), .CO(n1347), .S(n1348) );
  FA_X1 U1007 ( .A(n1385), .B(n1387), .CI(n1383), .CO(n1349), .S(n1350) );
  FA_X1 U1008 ( .A(n2336), .B(n1916), .CI(n1362), .CO(n1351), .S(n1352) );
  FA_X1 U1009 ( .A(n2305), .B(n2212), .CI(n1389), .CO(n1353), .S(n1354) );
  FA_X1 U1010 ( .A(n2151), .B(n2243), .CI(n2030), .CO(n1355), .S(n1356) );
  FA_X1 U1011 ( .A(n1970), .B(n2120), .CI(n1941), .CO(n1357), .S(n1358) );
  FA_X1 U1012 ( .A(n2274), .B(n1391), .CI(n2059), .CO(n1359), .S(n1360) );
  FA_X1 U1013 ( .A(n1999), .B(n2181), .CI(n2089), .CO(n1361), .S(n1362) );
  FA_X1 U1014 ( .A(n1395), .B(n1368), .CI(n1366), .CO(n1363), .S(n1364) );
  FA_X1 U1015 ( .A(n1370), .B(n1372), .CI(n1397), .CO(n1365), .S(n1366) );
  FA_X1 U1016 ( .A(n1401), .B(n1374), .CI(n1399), .CO(n1367), .S(n1368) );
  FA_X1 U1017 ( .A(n1403), .B(n1378), .CI(n1376), .CO(n1369), .S(n1370) );
  FA_X1 U1018 ( .A(n1380), .B(n1407), .CI(n1405), .CO(n1371), .S(n1372) );
  FA_X1 U1019 ( .A(n1382), .B(n1384), .CI(n1409), .CO(n1373), .S(n1374) );
  FA_X1 U1020 ( .A(n1411), .B(n1388), .CI(n1386), .CO(n1375), .S(n1376) );
  FA_X1 U1021 ( .A(n1415), .B(n1417), .CI(n1413), .CO(n1377), .S(n1378) );
  FA_X1 U1022 ( .A(n1917), .B(n2337), .CI(n1390), .CO(n1379), .S(n1380) );
  FA_X1 U1023 ( .A(n2306), .B(n2213), .CI(n1419), .CO(n1381), .S(n1382) );
  FA_X1 U1024 ( .A(n2182), .B(n2275), .CI(n1942), .CO(n1383), .S(n1384) );
  FA_X1 U1025 ( .A(n2000), .B(n2121), .CI(n2031), .CO(n1385), .S(n1386) );
  FA_X1 U1026 ( .A(n1421), .B(n2152), .CI(n2090), .CO(n1387), .S(n1388) );
  FA_X1 U1027 ( .A(n2244), .B(n1971), .CI(n1392), .CO(n1389), .S(n1390) );
  FA_X1 U1029 ( .A(n1425), .B(n1398), .CI(n1396), .CO(n1393), .S(n1394) );
  FA_X1 U1030 ( .A(n1400), .B(n1402), .CI(n1427), .CO(n1395), .S(n1396) );
  FA_X1 U1031 ( .A(n1404), .B(n1431), .CI(n1429), .CO(n1397), .S(n1398) );
  FA_X1 U1032 ( .A(n1433), .B(n1408), .CI(n1406), .CO(n1399), .S(n1400) );
  FA_X1 U1033 ( .A(n1410), .B(n1437), .CI(n1435), .CO(n1401), .S(n1402) );
  FA_X1 U1034 ( .A(n1439), .B(n1414), .CI(n1412), .CO(n1403), .S(n1404) );
  FA_X1 U1035 ( .A(n1418), .B(n1441), .CI(n1416), .CO(n1405), .S(n1406) );
  FA_X1 U1036 ( .A(n1443), .B(n1447), .CI(n1445), .CO(n1407), .S(n1408) );
  FA_X1 U1037 ( .A(n1420), .B(n2369), .CI(n1449), .CO(n1409), .S(n1410) );
  FA_X1 U1038 ( .A(n2338), .B(n2245), .CI(n1918), .CO(n1411), .S(n1412) );
  FA_X1 U1039 ( .A(n2183), .B(n2276), .CI(n2060), .CO(n1413), .S(n1414) );
  FA_X1 U1040 ( .A(n2001), .B(n2153), .CI(n1972), .CO(n1415), .S(n1416) );
  FA_X1 U1041 ( .A(n2091), .B(n1451), .CI(n1422), .CO(n1417), .S(n1418) );
  FA_X1 U1042 ( .A(n2214), .B(n2307), .CI(n2032), .CO(n1419), .S(n1420) );
  FA_X1 U1045 ( .A(n1455), .B(n1428), .CI(n1426), .CO(n1423), .S(n1424) );
  FA_X1 U1046 ( .A(n1430), .B(n1459), .CI(n1457), .CO(n1425), .S(n1426) );
  FA_X1 U1047 ( .A(n1434), .B(n1461), .CI(n1432), .CO(n1427), .S(n1428) );
  FA_X1 U1048 ( .A(n1438), .B(n1463), .CI(n1436), .CO(n1429), .S(n1430) );
  FA_X1 U1049 ( .A(n1440), .B(n1467), .CI(n1465), .CO(n1431), .S(n1432) );
  FA_X1 U1050 ( .A(n1448), .B(n1444), .CI(n1442), .CO(n1433), .S(n1434) );
  FA_X1 U1051 ( .A(n1450), .B(n1469), .CI(n1446), .CO(n1435), .S(n1436) );
  FA_X1 U1052 ( .A(n1473), .B(n1475), .CI(n1471), .CO(n1437), .S(n1438) );
  FA_X1 U1053 ( .A(n1919), .B(n2370), .CI(n1873), .CO(n1439), .S(n1440) );
  FA_X1 U1054 ( .A(n1479), .B(n1944), .CI(n1477), .CO(n1441), .S(n1442) );
  FA_X1 U1055 ( .A(n2339), .B(n2308), .CI(n1973), .CO(n1443), .S(n1444) );
  FA_X1 U1056 ( .A(n2215), .B(n2154), .CI(n2246), .CO(n1445), .S(n1446) );
  FA_X1 U1057 ( .A(n2033), .B(n2061), .CI(n1452), .CO(n1447), .S(n1448) );
  FA_X1 U1058 ( .A(n2092), .B(n2002), .CI(n2123), .CO(n1449), .S(n1450) );
  HA_X1 U1059 ( .A(n2184), .B(n2277), .CO(n1451), .S(n1452) );
  FA_X1 U1060 ( .A(n1483), .B(n1458), .CI(n1456), .CO(n1453), .S(n1454) );
  FA_X1 U1061 ( .A(n1460), .B(n1462), .CI(n1485), .CO(n1455), .S(n1456) );
  FA_X1 U1062 ( .A(n1489), .B(n1464), .CI(n1487), .CO(n1457), .S(n1458) );
  FA_X1 U1063 ( .A(n1491), .B(n1468), .CI(n1466), .CO(n1459), .S(n1460) );
  FA_X1 U1064 ( .A(n1470), .B(n1495), .CI(n1493), .CO(n1461), .S(n1462) );
  FA_X1 U1065 ( .A(n1474), .B(n1476), .CI(n1472), .CO(n1463), .S(n1464) );
  FA_X1 U1066 ( .A(n1499), .B(n1501), .CI(n1497), .CO(n1465), .S(n1466) );
  FA_X1 U1067 ( .A(n1478), .B(n1480), .CI(n1503), .CO(n1467), .S(n1468) );
  FA_X1 U1068 ( .A(n1945), .B(n2278), .CI(n1505), .CO(n1469), .S(n1470) );
  FA_X1 U1069 ( .A(n2185), .B(n2309), .CI(n2216), .CO(n1471), .S(n1472) );
  FA_X1 U1070 ( .A(n2371), .B(n2003), .CI(n2034), .CO(n1473), .S(n1474) );
  FA_X1 U1071 ( .A(n2093), .B(n1507), .CI(n2124), .CO(n1475), .S(n1476) );
  FA_X1 U1072 ( .A(n2247), .B(n2062), .CI(n1974), .CO(n1477), .S(n1478) );
  FA_X1 U1073 ( .A(n1920), .B(n2340), .CI(n2155), .CO(n1479), .S(n1480) );
  FA_X1 U1074 ( .A(n1511), .B(n1486), .CI(n1484), .CO(n1481), .S(n1482) );
  FA_X1 U1075 ( .A(n1488), .B(n1490), .CI(n1513), .CO(n1483), .S(n1484) );
  FA_X1 U1076 ( .A(n1492), .B(n1517), .CI(n1515), .CO(n1485), .S(n1486) );
  FA_X1 U1077 ( .A(n1519), .B(n1496), .CI(n1494), .CO(n1487), .S(n1488) );
  FA_X1 U1078 ( .A(n1523), .B(n1500), .CI(n1521), .CO(n1489), .S(n1490) );
  FA_X1 U1079 ( .A(n1502), .B(n1504), .CI(n1498), .CO(n1491), .S(n1492) );
  FA_X1 U1080 ( .A(n1525), .B(n1529), .CI(n1527), .CO(n1493), .S(n1494) );
  FA_X1 U1081 ( .A(n1531), .B(n1533), .CI(n1506), .CO(n1495), .S(n1496) );
  FA_X1 U1082 ( .A(n2248), .B(n2279), .CI(n1975), .CO(n1497), .S(n1498) );
  FA_X1 U1083 ( .A(n2004), .B(n2341), .CI(n2186), .CO(n1499), .S(n1500) );
  FA_X1 U1084 ( .A(n2372), .B(n2156), .CI(n1508), .CO(n1501), .S(n1502) );
  FA_X1 U1085 ( .A(n2094), .B(n2310), .CI(n2063), .CO(n1503), .S(n1504) );
  FA_X1 U1086 ( .A(n2217), .B(n1946), .CI(n2035), .CO(n1505), .S(n1506) );
  HA_X1 U1087 ( .A(n1874), .B(n2125), .CO(n1507), .S(n1508) );
  FA_X1 U1088 ( .A(n1537), .B(n1514), .CI(n1512), .CO(n1509), .S(n1510) );
  FA_X1 U1089 ( .A(n1516), .B(n1518), .CI(n1539), .CO(n1511), .S(n1512) );
  FA_X1 U1090 ( .A(n1520), .B(n1543), .CI(n1541), .CO(n1513), .S(n1514) );
  FA_X1 U1091 ( .A(n1545), .B(n1524), .CI(n1522), .CO(n1515), .S(n1516) );
  FA_X1 U1092 ( .A(n1526), .B(n1528), .CI(n1547), .CO(n1517), .S(n1518) );
  FA_X1 U1093 ( .A(n1549), .B(n1551), .CI(n1530), .CO(n1519), .S(n1520) );
  FA_X1 U1094 ( .A(n1555), .B(n1532), .CI(n1553), .CO(n1521), .S(n1522) );
  FA_X1 U1095 ( .A(n1557), .B(n1976), .CI(n1534), .CO(n1523), .S(n1524) );
  FA_X1 U1096 ( .A(n2249), .B(n2342), .CI(n2311), .CO(n1525), .S(n1526) );
  FA_X1 U1097 ( .A(n2157), .B(n2036), .CI(n2218), .CO(n1527), .S(n1528) );
  FA_X1 U1098 ( .A(n2126), .B(n1559), .CI(n2064), .CO(n1529), .S(n1530) );
  FA_X1 U1099 ( .A(n1947), .B(n2005), .CI(n2095), .CO(n1531), .S(n1532) );
  FA_X1 U1100 ( .A(n2187), .B(n2373), .CI(n2280), .CO(n1533), .S(n1534) );
  FA_X1 U1102 ( .A(n1542), .B(n1567), .CI(n1565), .CO(n1537), .S(n1538) );
  FA_X1 U1103 ( .A(n1546), .B(n1569), .CI(n1544), .CO(n1539), .S(n1540) );
  FA_X1 U1104 ( .A(n1571), .B(n1573), .CI(n1548), .CO(n1541), .S(n1542) );
  FA_X1 U1105 ( .A(n1552), .B(n1554), .CI(n1550), .CO(n1543), .S(n1544) );
  FA_X1 U1106 ( .A(n1575), .B(n1577), .CI(n1556), .CO(n1545), .S(n1546) );
  FA_X1 U1107 ( .A(n1558), .B(n1581), .CI(n1579), .CO(n1547), .S(n1548) );
  FA_X1 U1108 ( .A(n2006), .B(n2312), .CI(n1583), .CO(n1549), .S(n1550) );
  FA_X1 U1109 ( .A(n2219), .B(n2374), .CI(n2281), .CO(n1551), .S(n1552) );
  FA_X1 U1110 ( .A(n2188), .B(n2037), .CI(n1560), .CO(n1553), .S(n1554) );
  FA_X1 U1111 ( .A(n2127), .B(n1977), .CI(n2096), .CO(n1555), .S(n1556) );
  FA_X1 U1112 ( .A(n2250), .B(n1875), .CI(n2158), .CO(n1557), .S(n1558) );
  HA_X1 U1113 ( .A(n2343), .B(n2065), .CO(n1559), .S(n1560) );
  FA_X1 U1116 ( .A(n1572), .B(n1593), .CI(n1591), .CO(n1565), .S(n1566) );
  FA_X1 U1117 ( .A(n1595), .B(n1578), .CI(n1574), .CO(n1567), .S(n1568) );
  FA_X1 U1118 ( .A(n1597), .B(n1580), .CI(n1576), .CO(n1569), .S(n1570) );
  FA_X1 U1119 ( .A(n1599), .B(n1603), .CI(n1601), .CO(n1571), .S(n1572) );
  FA_X1 U1120 ( .A(n1584), .B(n1605), .CI(n1582), .CO(n1573), .S(n1574) );
  FA_X1 U1121 ( .A(n2251), .B(n2282), .CI(n2007), .CO(n1575), .S(n1576) );
  FA_X1 U1122 ( .A(n2097), .B(n2344), .CI(n2189), .CO(n1577), .S(n1578) );
  FA_X1 U1123 ( .A(n2066), .B(n2159), .CI(n2375), .CO(n1579), .S(n1580) );
  FA_X1 U1124 ( .A(n1978), .B(n2128), .CI(n1607), .CO(n1581), .S(n1582) );
  FA_X1 U1125 ( .A(n2220), .B(n2313), .CI(n2038), .CO(n1583), .S(n1584) );
  FA_X1 U1126 ( .A(n1611), .B(n1590), .CI(n1588), .CO(n1585), .S(n1586) );
  FA_X1 U1127 ( .A(n1592), .B(n1594), .CI(n1613), .CO(n1587), .S(n1588) );
  FA_X1 U1128 ( .A(n1596), .B(n1617), .CI(n1615), .CO(n1589), .S(n1590) );
  FA_X1 U1129 ( .A(n1598), .B(n1602), .CI(n1619), .CO(n1591), .S(n1592) );
  FA_X1 U1130 ( .A(n1604), .B(n1621), .CI(n1600), .CO(n1593), .S(n1594) );
  FA_X1 U1131 ( .A(n1625), .B(n1606), .CI(n1623), .CO(n1595), .S(n1596) );
  FA_X1 U1132 ( .A(n1629), .B(n2039), .CI(n1627), .CO(n1597), .S(n1598) );
  FA_X1 U1133 ( .A(n2160), .B(n2252), .CI(n2221), .CO(n1599), .S(n1600) );
  FA_X1 U1134 ( .A(n2314), .B(n2345), .CI(n1608), .CO(n1601), .S(n1602) );
  FA_X1 U1135 ( .A(n2129), .B(n1876), .CI(n2067), .CO(n1603), .S(n1604) );
  FA_X1 U1136 ( .A(n2008), .B(n2283), .CI(n2098), .CO(n1605), .S(n1606) );
  HA_X1 U1137 ( .A(n2376), .B(n2190), .CO(n1607), .S(n1608) );
  FA_X1 U1138 ( .A(n1633), .B(n1614), .CI(n1612), .CO(n1609), .S(n1610) );
  FA_X1 U1139 ( .A(n1616), .B(n1618), .CI(n1635), .CO(n1611), .S(n1612) );
  FA_X1 U1140 ( .A(n1620), .B(n1639), .CI(n1637), .CO(n1613), .S(n1614) );
  FA_X1 U1141 ( .A(n1641), .B(n1626), .CI(n1622), .CO(n1615), .S(n1616) );
  FA_X1 U1142 ( .A(n1643), .B(n1628), .CI(n1624), .CO(n1617), .S(n1618) );
  FA_X1 U1143 ( .A(n1647), .B(n1630), .CI(n1645), .CO(n1619), .S(n1620) );
  FA_X1 U1144 ( .A(n2040), .B(n2222), .CI(n1649), .CO(n1621), .S(n1622) );
  FA_X1 U1145 ( .A(n2099), .B(n2284), .CI(n2130), .CO(n1623), .S(n1624) );
  FA_X1 U1146 ( .A(n2377), .B(n2191), .CI(n2315), .CO(n1625), .S(n1626) );
  FA_X1 U1147 ( .A(n2253), .B(n2161), .CI(n1651), .CO(n1627), .S(n1628) );
  FA_X1 U1148 ( .A(n2068), .B(n2346), .CI(n2009), .CO(n1629), .S(n1630) );
  FA_X1 U1149 ( .A(n1655), .B(n1636), .CI(n1634), .CO(n1631), .S(n1632) );
  FA_X1 U1150 ( .A(n1638), .B(n1640), .CI(n1657), .CO(n1633), .S(n1634) );
  FA_X1 U1151 ( .A(n1642), .B(n1661), .CI(n1659), .CO(n1635), .S(n1636) );
  FA_X1 U1152 ( .A(n1644), .B(n1648), .CI(n1663), .CO(n1637), .S(n1638) );
  FA_X1 U1153 ( .A(n1665), .B(n1667), .CI(n1646), .CO(n1639), .S(n1640) );
  FA_X1 U1154 ( .A(n1669), .B(n1671), .CI(n1650), .CO(n1641), .S(n1642) );
  FA_X1 U1155 ( .A(n2254), .B(n2285), .CI(n2069), .CO(n1643), .S(n1644) );
  FA_X1 U1156 ( .A(n2347), .B(n2100), .CI(n2192), .CO(n1645), .S(n1646) );
  FA_X1 U1157 ( .A(n2378), .B(n2162), .CI(n1652), .CO(n1647), .S(n1648) );
  FA_X1 U1158 ( .A(n2041), .B(n2223), .CI(n1877), .CO(n1649), .S(n1650) );
  HA_X1 U1159 ( .A(n2131), .B(n2316), .CO(n1651), .S(n1652) );
  FA_X1 U1160 ( .A(n1675), .B(n1658), .CI(n1656), .CO(n1653), .S(n1654) );
  FA_X1 U1161 ( .A(n1660), .B(n1662), .CI(n1677), .CO(n1655), .S(n1656) );
  FA_X1 U1162 ( .A(n1664), .B(n1681), .CI(n1679), .CO(n1657), .S(n1658) );
  FA_X1 U1163 ( .A(n1666), .B(n1683), .CI(n1668), .CO(n1659), .S(n1660) );
  FA_X1 U1164 ( .A(n1685), .B(n1687), .CI(n1670), .CO(n1661), .S(n1662) );
  FA_X1 U1165 ( .A(n1689), .B(n2070), .CI(n1672), .CO(n1663), .S(n1664) );
  FA_X1 U1166 ( .A(n2224), .B(n2317), .CI(n2255), .CO(n1665), .S(n1666) );
  FA_X1 U1167 ( .A(n2348), .B(n2163), .CI(n2132), .CO(n1667), .S(n1668) );
  FA_X1 U1168 ( .A(n2101), .B(n2042), .CI(n1691), .CO(n1669), .S(n1670) );
  FA_X1 U1169 ( .A(n2193), .B(n2379), .CI(n2286), .CO(n1671), .S(n1672) );
  FA_X1 U1170 ( .A(n1695), .B(n1678), .CI(n1676), .CO(n1673), .S(n1674) );
  FA_X1 U1171 ( .A(n1680), .B(n1682), .CI(n1697), .CO(n1675), .S(n1676) );
  FA_X1 U1172 ( .A(n1701), .B(n1684), .CI(n1699), .CO(n1677), .S(n1678) );
  FA_X1 U1173 ( .A(n1686), .B(n1703), .CI(n1688), .CO(n1679), .S(n1680) );
  FA_X1 U1174 ( .A(n1707), .B(n1690), .CI(n1705), .CO(n1681), .S(n1682) );
  FA_X1 U1175 ( .A(n2102), .B(n2225), .CI(n1709), .CO(n1683), .S(n1684) );
  FA_X1 U1176 ( .A(n2287), .B(n2318), .CI(n2194), .CO(n1685), .S(n1686) );
  FA_X1 U1177 ( .A(n2380), .B(n2133), .CI(n1692), .CO(n1687), .S(n1688) );
  FA_X1 U1178 ( .A(n2256), .B(n2071), .CI(n2164), .CO(n1689), .S(n1690) );
  HA_X1 U1179 ( .A(n1878), .B(n2349), .CO(n1691), .S(n1692) );
  FA_X1 U1180 ( .A(n1713), .B(n1698), .CI(n1696), .CO(n1693), .S(n1694) );
  FA_X1 U1181 ( .A(n1700), .B(n1702), .CI(n1715), .CO(n1695), .S(n1696) );
  FA_X1 U1182 ( .A(n1719), .B(n1704), .CI(n1717), .CO(n1697), .S(n1698) );
  FA_X1 U1183 ( .A(n1708), .B(n1721), .CI(n1706), .CO(n1699), .S(n1700) );
  FA_X1 U1184 ( .A(n1710), .B(n1725), .CI(n1723), .CO(n1701), .S(n1702) );
  FA_X1 U1185 ( .A(n2288), .B(n2350), .CI(n2103), .CO(n1703), .S(n1704) );
  FA_X1 U1186 ( .A(n2381), .B(n2257), .CI(n2165), .CO(n1705), .S(n1706) );
  FA_X1 U1187 ( .A(n1727), .B(n2134), .CI(n2195), .CO(n1707), .S(n1708) );
  FA_X1 U1188 ( .A(n2072), .B(n2319), .CI(n2226), .CO(n1709), .S(n1710) );
  FA_X1 U1189 ( .A(n1731), .B(n1716), .CI(n1714), .CO(n1711), .S(n1712) );
  FA_X1 U1190 ( .A(n1718), .B(n1720), .CI(n1733), .CO(n1713), .S(n1714) );
  FA_X1 U1191 ( .A(n1737), .B(n1724), .CI(n1735), .CO(n1715), .S(n1716) );
  FA_X1 U1192 ( .A(n1739), .B(n1741), .CI(n1722), .CO(n1717), .S(n1718) );
  FA_X1 U1193 ( .A(n1743), .B(n2135), .CI(n1726), .CO(n1719), .S(n1720) );
  FA_X1 U1194 ( .A(n2227), .B(n2320), .CI(n2258), .CO(n1721), .S(n1722) );
  FA_X1 U1195 ( .A(n2351), .B(n2166), .CI(n1728), .CO(n1723), .S(n1724) );
  FA_X1 U1196 ( .A(n1879), .B(n2289), .CI(n2104), .CO(n1725), .S(n1726) );
  HA_X1 U1197 ( .A(n2382), .B(n2196), .CO(n1727), .S(n1728) );
  FA_X1 U1198 ( .A(n1734), .B(n1747), .CI(n1732), .CO(n1729), .S(n1730) );
  FA_X1 U1199 ( .A(n1736), .B(n1738), .CI(n1749), .CO(n1731), .S(n1732) );
  FA_X1 U1200 ( .A(n1740), .B(n1742), .CI(n1751), .CO(n1733), .S(n1734) );
  FA_X1 U1201 ( .A(n1755), .B(n1757), .CI(n1753), .CO(n1735), .S(n1736) );
  FA_X1 U1202 ( .A(n2136), .B(n2383), .CI(n1744), .CO(n1737), .S(n1738) );
  FA_X1 U1203 ( .A(n2290), .B(n2197), .CI(n2321), .CO(n1739), .S(n1740) );
  FA_X1 U1204 ( .A(n1759), .B(n2259), .CI(n2228), .CO(n1741), .S(n1742) );
  FA_X1 U1205 ( .A(n2167), .B(n2352), .CI(n2105), .CO(n1743), .S(n1744) );
  FA_X1 U1206 ( .A(n1763), .B(n1750), .CI(n1748), .CO(n1745), .S(n1746) );
  FA_X1 U1207 ( .A(n1765), .B(n1767), .CI(n1752), .CO(n1747), .S(n1748) );
  FA_X1 U1208 ( .A(n1756), .B(n1758), .CI(n1754), .CO(n1749), .S(n1750) );
  FA_X1 U1209 ( .A(n1771), .B(n1773), .CI(n1769), .CO(n1751), .S(n1752) );
  FA_X1 U1210 ( .A(n2353), .B(n2384), .CI(n2168), .CO(n1753), .S(n1754) );
  FA_X1 U1211 ( .A(n2291), .B(n2198), .CI(n1760), .CO(n1755), .S(n1756) );
  FA_X1 U1212 ( .A(n2229), .B(n2137), .CI(n2260), .CO(n1757), .S(n1758) );
  HA_X1 U1213 ( .A(n1880), .B(n2322), .CO(n1759), .S(n1760) );
  FA_X1 U1214 ( .A(n1777), .B(n1766), .CI(n1764), .CO(n1761), .S(n1762) );
  FA_X1 U1215 ( .A(n1779), .B(n1770), .CI(n1768), .CO(n1763), .S(n1764) );
  FA_X1 U1216 ( .A(n1781), .B(n1783), .CI(n1772), .CO(n1765), .S(n1766) );
  FA_X1 U1217 ( .A(n1774), .B(n2169), .CI(n1785), .CO(n1767), .S(n1768) );
  FA_X1 U1218 ( .A(n2323), .B(n2354), .CI(n2261), .CO(n1769), .S(n1770) );
  FA_X1 U1219 ( .A(n1787), .B(n2138), .CI(n2230), .CO(n1771), .S(n1772) );
  FA_X1 U1220 ( .A(n2199), .B(n2385), .CI(n2292), .CO(n1773), .S(n1774) );
  FA_X1 U1221 ( .A(n1791), .B(n1780), .CI(n1778), .CO(n1775), .S(n1776) );
  FA_X1 U1222 ( .A(n1782), .B(n1784), .CI(n1793), .CO(n1777), .S(n1778) );
  FA_X1 U1223 ( .A(n1795), .B(n1797), .CI(n1786), .CO(n1779), .S(n1780) );
  FA_X1 U1224 ( .A(n2200), .B(n2324), .CI(n1799), .CO(n1781), .S(n1782) );
  FA_X1 U1225 ( .A(n2293), .B(n2386), .CI(n1788), .CO(n1783), .S(n1784) );
  FA_X1 U1226 ( .A(n2170), .B(n2262), .CI(n2231), .CO(n1785), .S(n1786) );
  HA_X1 U1227 ( .A(n2355), .B(n1881), .CO(n1787), .S(n1788) );
  FA_X1 U1228 ( .A(n1803), .B(n1794), .CI(n1792), .CO(n1789), .S(n1790) );
  FA_X1 U1229 ( .A(n1796), .B(n1798), .CI(n1805), .CO(n1791), .S(n1792) );
  FA_X1 U1230 ( .A(n1809), .B(n1800), .CI(n1807), .CO(n1793), .S(n1794) );
  FA_X1 U1231 ( .A(n2356), .B(n2387), .CI(n2201), .CO(n1795), .S(n1796) );
  FA_X1 U1232 ( .A(n2294), .B(n1811), .CI(n2263), .CO(n1797), .S(n1798) );
  FA_X1 U1233 ( .A(n2171), .B(n2325), .CI(n2232), .CO(n1799), .S(n1800) );
  FA_X1 U1234 ( .A(n1806), .B(n1815), .CI(n1804), .CO(n1801), .S(n1802) );
  FA_X1 U1235 ( .A(n1808), .B(n1810), .CI(n1817), .CO(n1803), .S(n1804) );
  FA_X1 U1236 ( .A(n1821), .B(n2233), .CI(n1819), .CO(n1805), .S(n1806) );
  FA_X1 U1237 ( .A(n2326), .B(n2357), .CI(n1812), .CO(n1807), .S(n1808) );
  FA_X1 U1238 ( .A(n2295), .B(n2202), .CI(n2264), .CO(n1809), .S(n1810) );
  HA_X1 U1239 ( .A(n2388), .B(n1882), .CO(n1811), .S(n1812) );
  FA_X1 U1240 ( .A(n1825), .B(n1818), .CI(n1816), .CO(n1813), .S(n1814) );
  FA_X1 U1241 ( .A(n1827), .B(n1829), .CI(n1820), .CO(n1815), .S(n1816) );
  FA_X1 U1242 ( .A(n2234), .B(n2327), .CI(n1822), .CO(n1817), .S(n1818) );
  FA_X1 U1243 ( .A(n2296), .B(n1831), .CI(n2389), .CO(n1819), .S(n1820) );
  FA_X1 U1244 ( .A(n2203), .B(n2358), .CI(n2265), .CO(n1821), .S(n1822) );
  FA_X1 U1245 ( .A(n1835), .B(n1828), .CI(n1826), .CO(n1823), .S(n1824) );
  FA_X1 U1246 ( .A(n1837), .B(n1839), .CI(n1830), .CO(n1825), .S(n1826) );
  FA_X1 U1247 ( .A(n1832), .B(n2359), .CI(n2266), .CO(n1827), .S(n1828) );
  FA_X1 U1248 ( .A(n2297), .B(n2235), .CI(n2390), .CO(n1829), .S(n1830) );
  HA_X1 U1249 ( .A(n2328), .B(n1883), .CO(n1831), .S(n1832) );
  FA_X1 U1250 ( .A(n1843), .B(n1838), .CI(n1836), .CO(n1833), .S(n1834) );
  FA_X1 U1251 ( .A(n1840), .B(n2267), .CI(n1845), .CO(n1835), .S(n1836) );
  FA_X1 U1252 ( .A(n2360), .B(n1847), .CI(n2329), .CO(n1837), .S(n1838) );
  FA_X1 U1253 ( .A(n2298), .B(n2391), .CI(n2236), .CO(n1839), .S(n1840) );
  FA_X1 U1254 ( .A(n1846), .B(n1851), .CI(n1844), .CO(n1841), .S(n1842) );
  FA_X1 U1255 ( .A(n2299), .B(n1848), .CI(n1853), .CO(n1843), .S(n1844) );
  FA_X1 U1256 ( .A(n2392), .B(n2268), .CI(n2330), .CO(n1845), .S(n1846) );
  HA_X1 U1257 ( .A(n2361), .B(n1884), .CO(n1847), .S(n1848) );
  FA_X1 U1258 ( .A(n1854), .B(n1857), .CI(n1852), .CO(n1849), .S(n1850) );
  FA_X1 U1259 ( .A(n2362), .B(n2393), .CI(n2300), .CO(n1851), .S(n1852) );
  FA_X1 U1260 ( .A(n2269), .B(n2331), .CI(n1859), .CO(n1853), .S(n1854) );
  FA_X1 U1261 ( .A(n1863), .B(n2332), .CI(n1858), .CO(n1855), .S(n1856) );
  FA_X1 U1262 ( .A(n2363), .B(n2301), .CI(n1860), .CO(n1857), .S(n1858) );
  HA_X1 U1263 ( .A(n2394), .B(n1885), .CO(n1859), .S(n1860) );
  FA_X1 U1264 ( .A(n2333), .B(n2395), .CI(n1864), .CO(n1861), .S(n1862) );
  FA_X1 U1265 ( .A(n2302), .B(n2364), .CI(n1867), .CO(n1863), .S(n1864) );
  FA_X1 U1266 ( .A(n1868), .B(n2396), .CI(n2365), .CO(n1865), .S(n1866) );
  HA_X1 U1267 ( .A(n1886), .B(n2334), .CO(n1867), .S(n1868) );
  FA_X1 U1268 ( .A(n2335), .B(n2397), .CI(n1871), .CO(n1869), .S(n1870) );
  HA_X1 U1269 ( .A(n1887), .B(n2367), .CO(n1871), .S(n1872) );
  OAI22_X2 U1270 ( .A1(n3188), .A2(n3009), .B1(n2433), .B2(n3186), .ZN(n1873)
         );
  OAI22_X2 U1271 ( .A1(n3190), .A2(n2402), .B1(n2401), .B2(n3186), .ZN(n943)
         );
  OAI22_X2 U1272 ( .A1(n3189), .A2(n2403), .B1(n2402), .B2(n3186), .ZN(n1890)
         );
  OAI22_X2 U1273 ( .A1(n3190), .A2(n2404), .B1(n2403), .B2(n3186), .ZN(n1891)
         );
  OAI22_X2 U1274 ( .A1(n3189), .A2(n2405), .B1(n2404), .B2(n3186), .ZN(n1892)
         );
  OAI22_X2 U1275 ( .A1(n3189), .A2(n2406), .B1(n2405), .B2(n3186), .ZN(n1893)
         );
  OAI22_X2 U1276 ( .A1(n3190), .A2(n2407), .B1(n2406), .B2(n3186), .ZN(n1894)
         );
  OAI22_X2 U1277 ( .A1(n3190), .A2(n2408), .B1(n2407), .B2(n3186), .ZN(n1895)
         );
  OAI22_X2 U1278 ( .A1(n3189), .A2(n2409), .B1(n2408), .B2(n3186), .ZN(n1896)
         );
  OAI22_X2 U1279 ( .A1(n3190), .A2(n2410), .B1(n2409), .B2(n3186), .ZN(n1897)
         );
  OAI22_X2 U1280 ( .A1(n3190), .A2(n2411), .B1(n2410), .B2(n3186), .ZN(n1898)
         );
  OAI22_X2 U1281 ( .A1(n3189), .A2(n2412), .B1(n2411), .B2(n3186), .ZN(n1899)
         );
  OAI22_X2 U1282 ( .A1(n3189), .A2(n2413), .B1(n2412), .B2(n3186), .ZN(n1900)
         );
  OAI22_X2 U1283 ( .A1(n3190), .A2(n2414), .B1(n2413), .B2(n3186), .ZN(n1901)
         );
  OAI22_X2 U1284 ( .A1(n3190), .A2(n2415), .B1(n2414), .B2(n3186), .ZN(n1902)
         );
  OAI22_X2 U1285 ( .A1(n3190), .A2(n2416), .B1(n2415), .B2(n3186), .ZN(n1903)
         );
  OAI22_X2 U1286 ( .A1(n3190), .A2(n2417), .B1(n2416), .B2(n3186), .ZN(n1904)
         );
  OAI22_X2 U1287 ( .A1(n3189), .A2(n2418), .B1(n2417), .B2(n3186), .ZN(n1905)
         );
  OAI22_X2 U1288 ( .A1(n3189), .A2(n2419), .B1(n2418), .B2(n3186), .ZN(n1906)
         );
  OAI22_X2 U1289 ( .A1(n3190), .A2(n2420), .B1(n2419), .B2(n3186), .ZN(n1907)
         );
  OAI22_X2 U1290 ( .A1(n3189), .A2(n2421), .B1(n2420), .B2(n3186), .ZN(n1908)
         );
  OAI22_X2 U1291 ( .A1(n3190), .A2(n2422), .B1(n2421), .B2(n3186), .ZN(n1909)
         );
  OAI22_X2 U1292 ( .A1(n3189), .A2(n2423), .B1(n2422), .B2(n3186), .ZN(n1910)
         );
  OAI22_X2 U1293 ( .A1(n3189), .A2(n2424), .B1(n2423), .B2(n3186), .ZN(n1911)
         );
  OAI22_X2 U1294 ( .A1(n3190), .A2(n2425), .B1(n2424), .B2(n3186), .ZN(n1912)
         );
  OAI22_X2 U1295 ( .A1(n3189), .A2(n2426), .B1(n2425), .B2(n3186), .ZN(n1913)
         );
  OAI22_X2 U1296 ( .A1(n3190), .A2(n2427), .B1(n2426), .B2(n3186), .ZN(n1914)
         );
  OAI22_X2 U1297 ( .A1(n3189), .A2(n2428), .B1(n2427), .B2(n3186), .ZN(n1915)
         );
  OAI22_X2 U1298 ( .A1(n3190), .A2(n2429), .B1(n2428), .B2(n3186), .ZN(n1916)
         );
  OAI22_X2 U1299 ( .A1(n3189), .A2(n2430), .B1(n2429), .B2(n3186), .ZN(n1917)
         );
  OAI22_X2 U1301 ( .A1(n3188), .A2(n2432), .B1(n2431), .B2(n3186), .ZN(n1919)
         );
  OAI22_X2 U1334 ( .A1(n3204), .A2(n3010), .B1(n389), .B2(n2466), .ZN(n1874)
         );
  OAI22_X2 U1336 ( .A1(n2436), .A2(n3204), .B1(n389), .B2(n2435), .ZN(n1922)
         );
  OAI22_X2 U1337 ( .A1(n2436), .A2(n389), .B1(n3204), .B2(n2437), .ZN(n959) );
  OAI22_X2 U1340 ( .A1(n2439), .A2(n389), .B1(n3204), .B2(n2440), .ZN(n1925)
         );
  OAI22_X2 U1343 ( .A1(n2442), .A2(n389), .B1(n3204), .B2(n2443), .ZN(n1927)
         );
  OAI22_X2 U1348 ( .A1(n2448), .A2(n3204), .B1(n389), .B2(n2447), .ZN(n1931)
         );
  OAI22_X2 U1349 ( .A1(n2448), .A2(n389), .B1(n3204), .B2(n2449), .ZN(n1932)
         );
  OAI22_X2 U1350 ( .A1(n3204), .A2(n2450), .B1(n389), .B2(n2449), .ZN(n1933)
         );
  OAI22_X2 U1352 ( .A1(n2451), .A2(n389), .B1(n3204), .B2(n2452), .ZN(n1935)
         );
  OAI22_X2 U1353 ( .A1(n3203), .A2(n2453), .B1(n389), .B2(n2452), .ZN(n1183)
         );
  OAI22_X2 U1356 ( .A1(n3204), .A2(n2456), .B1(n389), .B2(n2455), .ZN(n1938)
         );
  OAI22_X2 U1357 ( .A1(n2457), .A2(n3204), .B1(n389), .B2(n2456), .ZN(n1939)
         );
  OAI22_X2 U1358 ( .A1(n2457), .A2(n389), .B1(n3204), .B2(n2458), .ZN(n1940)
         );
  OAI22_X2 U1359 ( .A1(n3204), .A2(n2459), .B1(n389), .B2(n2458), .ZN(n1333)
         );
  OAI22_X2 U1363 ( .A1(n2463), .A2(n3204), .B1(n389), .B2(n2462), .ZN(n1944)
         );
  OAI22_X2 U1364 ( .A1(n2463), .A2(n389), .B1(n3204), .B2(n2464), .ZN(n1945)
         );
  OAI22_X2 U1399 ( .A1(n2467), .A2(n386), .B1(n434), .B2(n2468), .ZN(n1949) );
  OAI22_X2 U1400 ( .A1(n2469), .A2(n434), .B1(n386), .B2(n2468), .ZN(n1950) );
  OAI22_X2 U1401 ( .A1(n2469), .A2(n386), .B1(n434), .B2(n2470), .ZN(n973) );
  OAI22_X2 U1402 ( .A1(n434), .A2(n2471), .B1(n386), .B2(n2470), .ZN(n1951) );
  OAI22_X2 U1403 ( .A1(n2472), .A2(n434), .B1(n386), .B2(n2471), .ZN(n1952) );
  OAI22_X2 U1404 ( .A1(n2472), .A2(n386), .B1(n434), .B2(n2473), .ZN(n1953) );
  OAI22_X2 U1405 ( .A1(n434), .A2(n2474), .B1(n386), .B2(n2473), .ZN(n1013) );
  OAI22_X2 U1406 ( .A1(n2475), .A2(n434), .B1(n386), .B2(n2474), .ZN(n1954) );
  OAI22_X2 U1407 ( .A1(n2475), .A2(n386), .B1(n434), .B2(n2476), .ZN(n1955) );
  OAI22_X2 U1408 ( .A1(n434), .A2(n2477), .B1(n386), .B2(n2476), .ZN(n1956) );
  OAI22_X2 U1409 ( .A1(n2478), .A2(n434), .B1(n386), .B2(n2477), .ZN(n1957) );
  OAI22_X2 U1410 ( .A1(n2478), .A2(n386), .B1(n434), .B2(n2479), .ZN(n1958) );
  OAI22_X2 U1411 ( .A1(n434), .A2(n2480), .B1(n386), .B2(n2479), .ZN(n1959) );
  OAI22_X2 U1412 ( .A1(n2481), .A2(n434), .B1(n386), .B2(n2480), .ZN(n1960) );
  OAI22_X2 U1413 ( .A1(n2481), .A2(n386), .B1(n434), .B2(n2482), .ZN(n1961) );
  OAI22_X2 U1414 ( .A1(n434), .A2(n2483), .B1(n386), .B2(n2482), .ZN(n1962) );
  OAI22_X2 U1415 ( .A1(n2484), .A2(n434), .B1(n386), .B2(n2483), .ZN(n1963) );
  OAI22_X2 U1416 ( .A1(n2484), .A2(n386), .B1(n434), .B2(n2485), .ZN(n1964) );
  OAI22_X2 U1417 ( .A1(n434), .A2(n2486), .B1(n386), .B2(n2485), .ZN(n1965) );
  OAI22_X2 U1418 ( .A1(n2487), .A2(n434), .B1(n386), .B2(n2486), .ZN(n1966) );
  OAI22_X2 U1419 ( .A1(n2487), .A2(n386), .B1(n434), .B2(n2488), .ZN(n1967) );
  OAI22_X2 U1420 ( .A1(n434), .A2(n2489), .B1(n386), .B2(n2488), .ZN(n1968) );
  OAI22_X2 U1421 ( .A1(n2490), .A2(n434), .B1(n386), .B2(n2489), .ZN(n1969) );
  OAI22_X2 U1422 ( .A1(n2490), .A2(n386), .B1(n434), .B2(n2491), .ZN(n1970) );
  OAI22_X2 U1423 ( .A1(n434), .A2(n2492), .B1(n386), .B2(n2491), .ZN(n1971) );
  OAI22_X2 U1424 ( .A1(n2493), .A2(n434), .B1(n386), .B2(n2492), .ZN(n1972) );
  OAI22_X2 U1425 ( .A1(n2493), .A2(n386), .B1(n434), .B2(n2494), .ZN(n1973) );
  OAI22_X2 U1427 ( .A1(n2496), .A2(n434), .B1(n386), .B2(n2495), .ZN(n1975) );
  OAI22_X2 U1428 ( .A1(n2496), .A2(n386), .B1(n434), .B2(n2497), .ZN(n1976) );
  OAI22_X2 U1429 ( .A1(n434), .A2(n2498), .B1(n386), .B2(n2497), .ZN(n1977) );
  OAI22_X2 U1462 ( .A1(n431), .A2(n3012), .B1(n3212), .B2(n2532), .ZN(n1876)
         );
  OAI22_X2 U1463 ( .A1(n2500), .A2(n3212), .B1(n431), .B2(n2501), .ZN(n1980)
         );
  OAI22_X2 U1464 ( .A1(n2502), .A2(n431), .B1(n3213), .B2(n2501), .ZN(n1981)
         );
  OAI22_X2 U1465 ( .A1(n2502), .A2(n3212), .B1(n431), .B2(n2503), .ZN(n1982)
         );
  OAI22_X2 U1466 ( .A1(n431), .A2(n2504), .B1(n3213), .B2(n2503), .ZN(n1983)
         );
  OAI22_X2 U1467 ( .A1(n2505), .A2(n431), .B1(n3212), .B2(n2504), .ZN(n1984)
         );
  OAI22_X2 U1468 ( .A1(n2505), .A2(n3213), .B1(n431), .B2(n2506), .ZN(n1985)
         );
  OAI22_X2 U1469 ( .A1(n431), .A2(n2507), .B1(n3213), .B2(n2506), .ZN(n1039)
         );
  OAI22_X2 U1470 ( .A1(n2508), .A2(n431), .B1(n3213), .B2(n2507), .ZN(n1986)
         );
  OAI22_X2 U1471 ( .A1(n2508), .A2(n3213), .B1(n431), .B2(n2509), .ZN(n1987)
         );
  OAI22_X2 U1472 ( .A1(n431), .A2(n2510), .B1(n3212), .B2(n2509), .ZN(n1988)
         );
  OAI22_X2 U1473 ( .A1(n2511), .A2(n431), .B1(n3213), .B2(n2510), .ZN(n1989)
         );
  OAI22_X2 U1474 ( .A1(n2511), .A2(n3213), .B1(n431), .B2(n2512), .ZN(n1990)
         );
  OAI22_X2 U1475 ( .A1(n431), .A2(n2513), .B1(n3212), .B2(n2512), .ZN(n1141)
         );
  OAI22_X2 U1476 ( .A1(n2514), .A2(n431), .B1(n3212), .B2(n2513), .ZN(n1991)
         );
  OAI22_X2 U1477 ( .A1(n2514), .A2(n3212), .B1(n431), .B2(n2515), .ZN(n1992)
         );
  OAI22_X2 U1478 ( .A1(n431), .A2(n2516), .B1(n3213), .B2(n2515), .ZN(n1993)
         );
  OAI22_X2 U1479 ( .A1(n2517), .A2(n431), .B1(n3212), .B2(n2516), .ZN(n1994)
         );
  OAI22_X2 U1480 ( .A1(n2517), .A2(n3213), .B1(n431), .B2(n2518), .ZN(n1995)
         );
  OAI22_X2 U1481 ( .A1(n431), .A2(n2519), .B1(n3212), .B2(n2518), .ZN(n1996)
         );
  OAI22_X2 U1482 ( .A1(n2520), .A2(n431), .B1(n3212), .B2(n2519), .ZN(n1997)
         );
  OAI22_X2 U1483 ( .A1(n2520), .A2(n3213), .B1(n431), .B2(n2521), .ZN(n1998)
         );
  OAI22_X2 U1484 ( .A1(n431), .A2(n2522), .B1(n3212), .B2(n2521), .ZN(n1999)
         );
  OAI22_X2 U1485 ( .A1(n2523), .A2(n431), .B1(n3213), .B2(n2522), .ZN(n2000)
         );
  OAI22_X2 U1486 ( .A1(n2523), .A2(n3212), .B1(n431), .B2(n2524), .ZN(n2001)
         );
  OAI22_X2 U1487 ( .A1(n431), .A2(n2525), .B1(n3213), .B2(n2524), .ZN(n2002)
         );
  OAI22_X2 U1488 ( .A1(n2526), .A2(n431), .B1(n3212), .B2(n2525), .ZN(n2003)
         );
  OAI22_X2 U1489 ( .A1(n2526), .A2(n3213), .B1(n431), .B2(n2527), .ZN(n2004)
         );
  OAI22_X2 U1490 ( .A1(n431), .A2(n2528), .B1(n3212), .B2(n2527), .ZN(n2005)
         );
  OAI22_X2 U1491 ( .A1(n2529), .A2(n431), .B1(n3212), .B2(n2528), .ZN(n2006)
         );
  OAI22_X2 U1492 ( .A1(n2529), .A2(n3213), .B1(n431), .B2(n2530), .ZN(n2007)
         );
  OAI22_X2 U1493 ( .A1(n431), .A2(n2531), .B1(n3213), .B2(n2530), .ZN(n2008)
         );
  OAI22_X2 U1526 ( .A1(n428), .A2(n3013), .B1(n380), .B2(n2565), .ZN(n1877) );
  OAI22_X2 U1527 ( .A1(n2533), .A2(n380), .B1(n428), .B2(n2534), .ZN(n2011) );
  OAI22_X2 U1528 ( .A1(n2535), .A2(n428), .B1(n380), .B2(n2534), .ZN(n2012) );
  OAI22_X2 U1529 ( .A1(n2535), .A2(n380), .B1(n428), .B2(n2536), .ZN(n2013) );
  OAI22_X2 U1530 ( .A1(n428), .A2(n2537), .B1(n380), .B2(n2536), .ZN(n2014) );
  OAI22_X2 U1531 ( .A1(n2538), .A2(n428), .B1(n380), .B2(n2537), .ZN(n2015) );
  OAI22_X2 U1532 ( .A1(n2538), .A2(n380), .B1(n428), .B2(n2539), .ZN(n2016) );
  OAI22_X2 U1533 ( .A1(n428), .A2(n2540), .B1(n380), .B2(n2539), .ZN(n2017) );
  OAI22_X2 U1534 ( .A1(n2541), .A2(n428), .B1(n380), .B2(n2540), .ZN(n2018) );
  OAI22_X2 U1535 ( .A1(n2541), .A2(n380), .B1(n428), .B2(n2542), .ZN(n2019) );
  OAI22_X2 U1536 ( .A1(n428), .A2(n2543), .B1(n380), .B2(n2542), .ZN(n2020) );
  OAI22_X2 U1537 ( .A1(n2544), .A2(n428), .B1(n380), .B2(n2543), .ZN(n2021) );
  OAI22_X2 U1538 ( .A1(n2544), .A2(n380), .B1(n428), .B2(n2545), .ZN(n2022) );
  OAI22_X2 U1539 ( .A1(n428), .A2(n2546), .B1(n380), .B2(n2545), .ZN(n2023) );
  OAI22_X2 U1540 ( .A1(n2547), .A2(n428), .B1(n380), .B2(n2546), .ZN(n2024) );
  OAI22_X2 U1541 ( .A1(n2547), .A2(n380), .B1(n428), .B2(n2548), .ZN(n2025) );
  OAI22_X2 U1542 ( .A1(n428), .A2(n2549), .B1(n380), .B2(n2548), .ZN(n2026) );
  OAI22_X2 U1543 ( .A1(n2550), .A2(n428), .B1(n380), .B2(n2549), .ZN(n2027) );
  OAI22_X2 U1544 ( .A1(n2550), .A2(n380), .B1(n428), .B2(n2551), .ZN(n2028) );
  OAI22_X2 U1545 ( .A1(n428), .A2(n2552), .B1(n380), .B2(n2551), .ZN(n2029) );
  OAI22_X2 U1546 ( .A1(n2553), .A2(n428), .B1(n380), .B2(n2552), .ZN(n2030) );
  OAI22_X2 U1547 ( .A1(n2553), .A2(n380), .B1(n428), .B2(n2554), .ZN(n2031) );
  OAI22_X2 U1549 ( .A1(n2556), .A2(n428), .B1(n380), .B2(n2555), .ZN(n2033) );
  OAI22_X2 U1550 ( .A1(n2556), .A2(n380), .B1(n428), .B2(n2557), .ZN(n2034) );
  OAI22_X2 U1551 ( .A1(n428), .A2(n2558), .B1(n380), .B2(n2557), .ZN(n2035) );
  OAI22_X2 U1552 ( .A1(n2559), .A2(n428), .B1(n380), .B2(n2558), .ZN(n2036) );
  OAI22_X2 U1553 ( .A1(n2559), .A2(n380), .B1(n428), .B2(n2560), .ZN(n2037) );
  OAI22_X2 U1554 ( .A1(n428), .A2(n2561), .B1(n380), .B2(n2560), .ZN(n2038) );
  OAI22_X2 U1555 ( .A1(n2562), .A2(n428), .B1(n380), .B2(n2561), .ZN(n2039) );
  OAI22_X2 U1556 ( .A1(n2562), .A2(n380), .B1(n428), .B2(n2563), .ZN(n2040) );
  OAI22_X2 U1591 ( .A1(n2566), .A2(n3208), .B1(n425), .B2(n2567), .ZN(n2044)
         );
  OAI22_X2 U1592 ( .A1(n2568), .A2(n425), .B1(n3208), .B2(n2567), .ZN(n2045)
         );
  OAI22_X2 U1593 ( .A1(n2568), .A2(n3209), .B1(n425), .B2(n2569), .ZN(n2046)
         );
  OAI22_X2 U1594 ( .A1(n425), .A2(n2570), .B1(n3208), .B2(n2569), .ZN(n2047)
         );
  OAI22_X2 U1595 ( .A1(n2571), .A2(n425), .B1(n3208), .B2(n2570), .ZN(n2048)
         );
  OAI22_X2 U1596 ( .A1(n2571), .A2(n3209), .B1(n425), .B2(n2572), .ZN(n2049)
         );
  OAI22_X2 U1597 ( .A1(n425), .A2(n2573), .B1(n3209), .B2(n2572), .ZN(n1103)
         );
  OAI22_X2 U1598 ( .A1(n2574), .A2(n425), .B1(n3209), .B2(n2573), .ZN(n2050)
         );
  OAI22_X2 U1599 ( .A1(n2574), .A2(n3209), .B1(n425), .B2(n2575), .ZN(n2051)
         );
  OAI22_X2 U1600 ( .A1(n425), .A2(n2576), .B1(n3209), .B2(n2575), .ZN(n2052)
         );
  OAI22_X2 U1601 ( .A1(n2577), .A2(n425), .B1(n3209), .B2(n2576), .ZN(n2053)
         );
  OAI22_X2 U1602 ( .A1(n2577), .A2(n3208), .B1(n425), .B2(n2578), .ZN(n2054)
         );
  OAI22_X2 U1603 ( .A1(n425), .A2(n2579), .B1(n3208), .B2(n2578), .ZN(n1229)
         );
  OAI22_X2 U1604 ( .A1(n2580), .A2(n425), .B1(n3209), .B2(n2579), .ZN(n2055)
         );
  OAI22_X2 U1605 ( .A1(n2580), .A2(n3208), .B1(n425), .B2(n2581), .ZN(n2056)
         );
  OAI22_X2 U1606 ( .A1(n425), .A2(n2582), .B1(n3208), .B2(n2581), .ZN(n2057)
         );
  OAI22_X2 U1607 ( .A1(n2583), .A2(n425), .B1(n3209), .B2(n2582), .ZN(n2058)
         );
  OAI22_X2 U1608 ( .A1(n2583), .A2(n3208), .B1(n425), .B2(n2584), .ZN(n2059)
         );
  OAI22_X2 U1609 ( .A1(n425), .A2(n2585), .B1(n3208), .B2(n2584), .ZN(n1391)
         );
  OAI22_X2 U1610 ( .A1(n2586), .A2(n425), .B1(n3209), .B2(n2585), .ZN(n2060)
         );
  OAI22_X2 U1611 ( .A1(n2586), .A2(n3208), .B1(n425), .B2(n2587), .ZN(n2061)
         );
  OAI22_X2 U1612 ( .A1(n425), .A2(n2588), .B1(n3208), .B2(n2587), .ZN(n2062)
         );
  OAI22_X2 U1613 ( .A1(n2589), .A2(n425), .B1(n3208), .B2(n2588), .ZN(n2063)
         );
  OAI22_X2 U1614 ( .A1(n2589), .A2(n3209), .B1(n425), .B2(n2590), .ZN(n2064)
         );
  OAI22_X2 U1615 ( .A1(n425), .A2(n2591), .B1(n3209), .B2(n2590), .ZN(n2065)
         );
  OAI22_X2 U1616 ( .A1(n2592), .A2(n425), .B1(n3208), .B2(n2591), .ZN(n2066)
         );
  OAI22_X2 U1617 ( .A1(n2592), .A2(n3209), .B1(n425), .B2(n2593), .ZN(n2067)
         );
  OAI22_X2 U1618 ( .A1(n425), .A2(n2594), .B1(n3209), .B2(n2593), .ZN(n2068)
         );
  OAI22_X2 U1619 ( .A1(n2595), .A2(n425), .B1(n3209), .B2(n2594), .ZN(n2069)
         );
  OAI22_X2 U1620 ( .A1(n2595), .A2(n3208), .B1(n425), .B2(n2596), .ZN(n2070)
         );
  OAI22_X2 U1621 ( .A1(n425), .A2(n2597), .B1(n3209), .B2(n2596), .ZN(n2071)
         );
  OAI22_X2 U1655 ( .A1(n2599), .A2(n3193), .B1(n422), .B2(n2600), .ZN(n2074)
         );
  OAI22_X2 U1656 ( .A1(n2601), .A2(n422), .B1(n3193), .B2(n2600), .ZN(n2075)
         );
  OAI22_X2 U1657 ( .A1(n2601), .A2(n3193), .B1(n422), .B2(n2602), .ZN(n2076)
         );
  OAI22_X2 U1659 ( .A1(n2604), .A2(n422), .B1(n3193), .B2(n2603), .ZN(n2078)
         );
  OAI22_X2 U1660 ( .A1(n2604), .A2(n3193), .B1(n422), .B2(n2605), .ZN(n2079)
         );
  OAI22_X2 U1661 ( .A1(n422), .A2(n2606), .B1(n3193), .B2(n2605), .ZN(n2080)
         );
  OAI22_X2 U1662 ( .A1(n2607), .A2(n422), .B1(n3193), .B2(n2606), .ZN(n2081)
         );
  OAI22_X2 U1663 ( .A1(n2607), .A2(n3193), .B1(n422), .B2(n2608), .ZN(n2082)
         );
  OAI22_X2 U1665 ( .A1(n2610), .A2(n422), .B1(n3193), .B2(n2609), .ZN(n2084)
         );
  OAI22_X2 U1666 ( .A1(n2610), .A2(n3193), .B1(n422), .B2(n2611), .ZN(n2085)
         );
  OAI22_X2 U1668 ( .A1(n2613), .A2(n422), .B1(n3193), .B2(n2612), .ZN(n2087)
         );
  OAI22_X2 U1669 ( .A1(n2613), .A2(n3193), .B1(n422), .B2(n2614), .ZN(n2088)
         );
  OAI22_X2 U1671 ( .A1(n2616), .A2(n422), .B1(n3193), .B2(n2615), .ZN(n2090)
         );
  OAI22_X2 U1672 ( .A1(n2616), .A2(n3193), .B1(n422), .B2(n2617), .ZN(n2091)
         );
  OAI22_X2 U1674 ( .A1(n2619), .A2(n422), .B1(n3193), .B2(n2618), .ZN(n2093)
         );
  OAI22_X2 U1675 ( .A1(n2619), .A2(n3193), .B1(n422), .B2(n2620), .ZN(n2094)
         );
  OAI22_X2 U1678 ( .A1(n2622), .A2(n3193), .B1(n422), .B2(n2623), .ZN(n2097)
         );
  OAI22_X2 U1680 ( .A1(n2625), .A2(n422), .B1(n3193), .B2(n2624), .ZN(n2099)
         );
  OAI22_X2 U1683 ( .A1(n2628), .A2(n422), .B1(n3193), .B2(n2627), .ZN(n2102)
         );
  OAI22_X2 U1684 ( .A1(n2628), .A2(n3193), .B1(n422), .B2(n2629), .ZN(n2103)
         );
  OAI22_X2 U1718 ( .A1(n419), .A2(n3016), .B1(n3235), .B2(n2664), .ZN(n1880)
         );
  OAI22_X2 U1719 ( .A1(n2632), .A2(n3235), .B1(n419), .B2(n2633), .ZN(n2107)
         );
  OAI22_X2 U1720 ( .A1(n2634), .A2(n419), .B1(n3235), .B2(n2633), .ZN(n2108)
         );
  OAI22_X2 U1721 ( .A1(n2634), .A2(n3234), .B1(n419), .B2(n2635), .ZN(n2109)
         );
  OAI22_X2 U1722 ( .A1(n419), .A2(n2636), .B1(n3234), .B2(n2635), .ZN(n2110)
         );
  OAI22_X2 U1723 ( .A1(n2637), .A2(n419), .B1(n3234), .B2(n2636), .ZN(n2111)
         );
  OAI22_X2 U1724 ( .A1(n2637), .A2(n3234), .B1(n419), .B2(n2638), .ZN(n2112)
         );
  OAI22_X2 U1725 ( .A1(n419), .A2(n2639), .B1(n3234), .B2(n2638), .ZN(n2113)
         );
  OAI22_X2 U1726 ( .A1(n2640), .A2(n419), .B1(n3235), .B2(n2639), .ZN(n2114)
         );
  OAI22_X2 U1727 ( .A1(n2640), .A2(n3235), .B1(n419), .B2(n2641), .ZN(n2115)
         );
  OAI22_X2 U1728 ( .A1(n419), .A2(n2642), .B1(n3234), .B2(n2641), .ZN(n2116)
         );
  OAI22_X2 U1729 ( .A1(n2643), .A2(n419), .B1(n3235), .B2(n2642), .ZN(n2117)
         );
  OAI22_X2 U1730 ( .A1(n2643), .A2(n3234), .B1(n419), .B2(n2644), .ZN(n2118)
         );
  OAI22_X2 U1731 ( .A1(n419), .A2(n2645), .B1(n3235), .B2(n2644), .ZN(n2119)
         );
  OAI22_X2 U1732 ( .A1(n2646), .A2(n419), .B1(n3234), .B2(n2645), .ZN(n2120)
         );
  OAI22_X2 U1733 ( .A1(n2646), .A2(n3235), .B1(n419), .B2(n2647), .ZN(n2121)
         );
  OAI22_X2 U1734 ( .A1(n419), .A2(n2648), .B1(n3235), .B2(n2647), .ZN(n2122)
         );
  OAI22_X2 U1735 ( .A1(n2649), .A2(n419), .B1(n3234), .B2(n2648), .ZN(n2123)
         );
  OAI22_X2 U1736 ( .A1(n2649), .A2(n3235), .B1(n419), .B2(n2650), .ZN(n2124)
         );
  OAI22_X2 U1737 ( .A1(n419), .A2(n2651), .B1(n3234), .B2(n2650), .ZN(n2125)
         );
  OAI22_X2 U1738 ( .A1(n2652), .A2(n419), .B1(n3234), .B2(n2651), .ZN(n2126)
         );
  OAI22_X2 U1739 ( .A1(n2652), .A2(n3234), .B1(n419), .B2(n2653), .ZN(n2127)
         );
  OAI22_X2 U1740 ( .A1(n419), .A2(n2654), .B1(n3235), .B2(n2653), .ZN(n2128)
         );
  OAI22_X2 U1741 ( .A1(n2655), .A2(n419), .B1(n3235), .B2(n2654), .ZN(n2129)
         );
  OAI22_X2 U1742 ( .A1(n2655), .A2(n3235), .B1(n419), .B2(n2656), .ZN(n2130)
         );
  OAI22_X2 U1744 ( .A1(n2658), .A2(n419), .B1(n3234), .B2(n2657), .ZN(n2132)
         );
  OAI22_X2 U1745 ( .A1(n2658), .A2(n3235), .B1(n419), .B2(n2659), .ZN(n2133)
         );
  OAI22_X2 U1746 ( .A1(n419), .A2(n2660), .B1(n3235), .B2(n2659), .ZN(n2134)
         );
  OAI22_X2 U1747 ( .A1(n2661), .A2(n419), .B1(n3234), .B2(n2660), .ZN(n2135)
         );
  OAI22_X2 U1748 ( .A1(n2661), .A2(n3234), .B1(n419), .B2(n2662), .ZN(n2136)
         );
  OAI22_X2 U1749 ( .A1(n419), .A2(n2663), .B1(n3234), .B2(n2662), .ZN(n2137)
         );
  OAI22_X2 U1782 ( .A1(n416), .A2(n3017), .B1(n3198), .B2(n2697), .ZN(n1881)
         );
  OAI22_X2 U1783 ( .A1(n2665), .A2(n3197), .B1(n416), .B2(n2666), .ZN(n2140)
         );
  OAI22_X2 U1784 ( .A1(n2667), .A2(n416), .B1(n3198), .B2(n2666), .ZN(n2141)
         );
  OAI22_X2 U1785 ( .A1(n2667), .A2(n3198), .B1(n416), .B2(n2668), .ZN(n2142)
         );
  OAI22_X2 U1786 ( .A1(n416), .A2(n2669), .B1(n3198), .B2(n2668), .ZN(n2143)
         );
  OAI22_X2 U1787 ( .A1(n2670), .A2(n416), .B1(n3197), .B2(n2669), .ZN(n2144)
         );
  OAI22_X2 U1788 ( .A1(n2670), .A2(n3197), .B1(n416), .B2(n2671), .ZN(n2145)
         );
  OAI22_X2 U1789 ( .A1(n416), .A2(n2672), .B1(n3198), .B2(n2671), .ZN(n2146)
         );
  OAI22_X2 U1790 ( .A1(n2673), .A2(n416), .B1(n3198), .B2(n2672), .ZN(n2147)
         );
  OAI22_X2 U1791 ( .A1(n2673), .A2(n3197), .B1(n416), .B2(n2674), .ZN(n2148)
         );
  OAI22_X2 U1792 ( .A1(n416), .A2(n2675), .B1(n3197), .B2(n2674), .ZN(n2149)
         );
  OAI22_X2 U1793 ( .A1(n2676), .A2(n416), .B1(n3197), .B2(n2675), .ZN(n2150)
         );
  OAI22_X2 U1794 ( .A1(n2676), .A2(n3198), .B1(n416), .B2(n2677), .ZN(n2151)
         );
  OAI22_X2 U1795 ( .A1(n416), .A2(n2678), .B1(n3197), .B2(n2677), .ZN(n2152)
         );
  OAI22_X2 U1796 ( .A1(n2679), .A2(n416), .B1(n3197), .B2(n2678), .ZN(n2153)
         );
  OAI22_X2 U1797 ( .A1(n2679), .A2(n3197), .B1(n416), .B2(n2680), .ZN(n2154)
         );
  OAI22_X2 U1798 ( .A1(n416), .A2(n2681), .B1(n3197), .B2(n2680), .ZN(n2155)
         );
  OAI22_X2 U1799 ( .A1(n2682), .A2(n416), .B1(n3197), .B2(n2681), .ZN(n2156)
         );
  OAI22_X2 U1800 ( .A1(n2682), .A2(n3198), .B1(n416), .B2(n2683), .ZN(n2157)
         );
  OAI22_X2 U1801 ( .A1(n416), .A2(n2684), .B1(n3197), .B2(n2683), .ZN(n2158)
         );
  OAI22_X2 U1802 ( .A1(n2685), .A2(n416), .B1(n3198), .B2(n2684), .ZN(n2159)
         );
  OAI22_X2 U1803 ( .A1(n2685), .A2(n3197), .B1(n416), .B2(n2686), .ZN(n2160)
         );
  OAI22_X2 U1805 ( .A1(n2688), .A2(n416), .B1(n3198), .B2(n2687), .ZN(n2162)
         );
  OAI22_X2 U1806 ( .A1(n2688), .A2(n3197), .B1(n416), .B2(n2689), .ZN(n2163)
         );
  OAI22_X2 U1807 ( .A1(n416), .A2(n2690), .B1(n3197), .B2(n2689), .ZN(n2164)
         );
  OAI22_X2 U1808 ( .A1(n2691), .A2(n416), .B1(n3198), .B2(n2690), .ZN(n2165)
         );
  OAI22_X2 U1809 ( .A1(n2691), .A2(n3198), .B1(n416), .B2(n2692), .ZN(n2166)
         );
  OAI22_X2 U1810 ( .A1(n416), .A2(n2693), .B1(n3198), .B2(n2692), .ZN(n2167)
         );
  OAI22_X2 U1811 ( .A1(n2694), .A2(n416), .B1(n3198), .B2(n2693), .ZN(n2168)
         );
  OAI22_X2 U1812 ( .A1(n2694), .A2(n3198), .B1(n416), .B2(n2695), .ZN(n2169)
         );
  OAI22_X2 U1813 ( .A1(n416), .A2(n2696), .B1(n3198), .B2(n2695), .ZN(n2170)
         );
  OAI22_X2 U1846 ( .A1(n3223), .A2(n3018), .B1(n365), .B2(n2730), .ZN(n1882)
         );
  OAI22_X2 U1847 ( .A1(n2698), .A2(n365), .B1(n3223), .B2(n2699), .ZN(n2173)
         );
  OAI22_X2 U1848 ( .A1(n2700), .A2(n3223), .B1(n2699), .B2(n365), .ZN(n2174)
         );
  OAI22_X2 U1849 ( .A1(n2700), .A2(n365), .B1(n3223), .B2(n2701), .ZN(n2175)
         );
  OAI22_X2 U1850 ( .A1(n3223), .A2(n2702), .B1(n2701), .B2(n365), .ZN(n2176)
         );
  OAI22_X2 U1851 ( .A1(n2703), .A2(n3223), .B1(n2702), .B2(n365), .ZN(n2177)
         );
  OAI22_X2 U1852 ( .A1(n2703), .A2(n365), .B1(n3223), .B2(n2704), .ZN(n2178)
         );
  OAI22_X2 U1853 ( .A1(n3222), .A2(n2705), .B1(n2704), .B2(n365), .ZN(n1279)
         );
  OAI22_X2 U1854 ( .A1(n2706), .A2(n3223), .B1(n2705), .B2(n365), .ZN(n2179)
         );
  OAI22_X2 U1855 ( .A1(n2706), .A2(n365), .B1(n3223), .B2(n2707), .ZN(n2180)
         );
  OAI22_X2 U1856 ( .A1(n3223), .A2(n2708), .B1(n2707), .B2(n365), .ZN(n2181)
         );
  OAI22_X2 U1857 ( .A1(n2709), .A2(n3223), .B1(n2708), .B2(n365), .ZN(n2182)
         );
  OAI22_X2 U1858 ( .A1(n2709), .A2(n365), .B1(n3223), .B2(n2710), .ZN(n2183)
         );
  OAI22_X2 U1859 ( .A1(n3223), .A2(n2711), .B1(n2710), .B2(n365), .ZN(n2184)
         );
  OAI22_X2 U1860 ( .A1(n2712), .A2(n3223), .B1(n2711), .B2(n365), .ZN(n2185)
         );
  OAI22_X2 U1861 ( .A1(n2712), .A2(n365), .B1(n3223), .B2(n2713), .ZN(n2186)
         );
  OAI22_X2 U1862 ( .A1(n3223), .A2(n2714), .B1(n2713), .B2(n365), .ZN(n2187)
         );
  OAI22_X2 U1863 ( .A1(n2715), .A2(n3223), .B1(n2714), .B2(n365), .ZN(n2188)
         );
  OAI22_X2 U1864 ( .A1(n2715), .A2(n365), .B1(n3223), .B2(n2716), .ZN(n2189)
         );
  OAI22_X2 U1865 ( .A1(n3223), .A2(n2717), .B1(n2716), .B2(n365), .ZN(n2190)
         );
  OAI22_X2 U1866 ( .A1(n2718), .A2(n3223), .B1(n2717), .B2(n365), .ZN(n2191)
         );
  OAI22_X2 U1867 ( .A1(n2718), .A2(n365), .B1(n3223), .B2(n2719), .ZN(n2192)
         );
  OAI22_X2 U1868 ( .A1(n3222), .A2(n2720), .B1(n2719), .B2(n365), .ZN(n2193)
         );
  OAI22_X2 U1869 ( .A1(n2721), .A2(n3223), .B1(n2720), .B2(n365), .ZN(n2194)
         );
  OAI22_X2 U1870 ( .A1(n2721), .A2(n365), .B1(n3223), .B2(n2722), .ZN(n2195)
         );
  OAI22_X2 U1871 ( .A1(n3222), .A2(n2723), .B1(n2722), .B2(n365), .ZN(n2196)
         );
  OAI22_X2 U1872 ( .A1(n2724), .A2(n3223), .B1(n2723), .B2(n365), .ZN(n2197)
         );
  OAI22_X2 U1873 ( .A1(n2724), .A2(n365), .B1(n3223), .B2(n2725), .ZN(n2198)
         );
  OAI22_X2 U1874 ( .A1(n3223), .A2(n2726), .B1(n2725), .B2(n365), .ZN(n2199)
         );
  OAI22_X2 U1875 ( .A1(n2727), .A2(n3223), .B1(n2726), .B2(n365), .ZN(n2200)
         );
  OAI22_X2 U1876 ( .A1(n2727), .A2(n365), .B1(n3223), .B2(n2728), .ZN(n2201)
         );
  OAI22_X2 U1877 ( .A1(n3223), .A2(n2729), .B1(n2728), .B2(n365), .ZN(n2202)
         );
  OAI22_X2 U1910 ( .A1(n3183), .A2(n3019), .B1(n362), .B2(n2763), .ZN(n1883)
         );
  OAI22_X2 U1911 ( .A1(n2731), .A2(n362), .B1(n3183), .B2(n2732), .ZN(n2205)
         );
  OAI22_X2 U1912 ( .A1(n2733), .A2(n3183), .B1(n362), .B2(n2732), .ZN(n2206)
         );
  OAI22_X2 U1913 ( .A1(n2733), .A2(n362), .B1(n3182), .B2(n2734), .ZN(n2207)
         );
  OAI22_X2 U1914 ( .A1(n3183), .A2(n2735), .B1(n362), .B2(n2734), .ZN(n2208)
         );
  OAI22_X2 U1915 ( .A1(n2736), .A2(n3182), .B1(n362), .B2(n2735), .ZN(n2209)
         );
  OAI22_X2 U1916 ( .A1(n2736), .A2(n362), .B1(n3183), .B2(n2737), .ZN(n2210)
         );
  OAI22_X2 U1917 ( .A1(n3182), .A2(n2738), .B1(n362), .B2(n2737), .ZN(n2211)
         );
  OAI22_X2 U1918 ( .A1(n2739), .A2(n3183), .B1(n362), .B2(n2738), .ZN(n2212)
         );
  OAI22_X2 U1919 ( .A1(n2739), .A2(n362), .B1(n3182), .B2(n2740), .ZN(n2213)
         );
  OAI22_X2 U1920 ( .A1(n410), .A2(n2741), .B1(n362), .B2(n2740), .ZN(n2214) );
  OAI22_X2 U1921 ( .A1(n2742), .A2(n3183), .B1(n362), .B2(n2741), .ZN(n2215)
         );
  OAI22_X2 U1922 ( .A1(n2742), .A2(n362), .B1(n3182), .B2(n2743), .ZN(n2216)
         );
  OAI22_X2 U1923 ( .A1(n3183), .A2(n2744), .B1(n362), .B2(n2743), .ZN(n2217)
         );
  OAI22_X2 U1924 ( .A1(n2745), .A2(n3183), .B1(n362), .B2(n2744), .ZN(n2218)
         );
  OAI22_X2 U1925 ( .A1(n2745), .A2(n362), .B1(n3183), .B2(n2746), .ZN(n2219)
         );
  OAI22_X2 U1927 ( .A1(n2748), .A2(n3183), .B1(n362), .B2(n2747), .ZN(n2221)
         );
  OAI22_X2 U1928 ( .A1(n2748), .A2(n362), .B1(n3182), .B2(n2749), .ZN(n2222)
         );
  OAI22_X2 U1930 ( .A1(n2751), .A2(n3182), .B1(n362), .B2(n2750), .ZN(n2224)
         );
  OAI22_X2 U1931 ( .A1(n2751), .A2(n362), .B1(n3183), .B2(n2752), .ZN(n2225)
         );
  OAI22_X2 U1932 ( .A1(n3182), .A2(n2753), .B1(n362), .B2(n2752), .ZN(n2226)
         );
  OAI22_X2 U1933 ( .A1(n2754), .A2(n3182), .B1(n362), .B2(n2753), .ZN(n2227)
         );
  OAI22_X2 U1934 ( .A1(n2754), .A2(n362), .B1(n3183), .B2(n2755), .ZN(n2228)
         );
  OAI22_X2 U1935 ( .A1(n3183), .A2(n2756), .B1(n362), .B2(n2755), .ZN(n2229)
         );
  OAI22_X2 U1936 ( .A1(n2757), .A2(n3183), .B1(n362), .B2(n2756), .ZN(n2230)
         );
  OAI22_X2 U1937 ( .A1(n2757), .A2(n362), .B1(n3182), .B2(n2758), .ZN(n2231)
         );
  OAI22_X2 U1938 ( .A1(n3183), .A2(n2759), .B1(n362), .B2(n2758), .ZN(n2232)
         );
  OAI22_X2 U1939 ( .A1(n2760), .A2(n3182), .B1(n362), .B2(n2759), .ZN(n2233)
         );
  OAI22_X2 U1940 ( .A1(n2760), .A2(n362), .B1(n3183), .B2(n2761), .ZN(n2234)
         );
  OAI22_X2 U1941 ( .A1(n3182), .A2(n2762), .B1(n362), .B2(n2761), .ZN(n2235)
         );
  OAI22_X2 U1974 ( .A1(n407), .A2(n3020), .B1(n359), .B2(n2796), .ZN(n1884) );
  OAI22_X2 U1975 ( .A1(n2764), .A2(n359), .B1(n407), .B2(n2765), .ZN(n2238) );
  OAI22_X2 U1976 ( .A1(n2766), .A2(n407), .B1(n359), .B2(n2765), .ZN(n2239) );
  OAI22_X2 U1977 ( .A1(n2766), .A2(n359), .B1(n407), .B2(n2767), .ZN(n2240) );
  OAI22_X2 U1978 ( .A1(n407), .A2(n2768), .B1(n359), .B2(n2767), .ZN(n2241) );
  OAI22_X2 U1979 ( .A1(n2769), .A2(n407), .B1(n359), .B2(n2768), .ZN(n2242) );
  OAI22_X2 U1980 ( .A1(n2769), .A2(n359), .B1(n407), .B2(n2770), .ZN(n2243) );
  OAI22_X2 U1981 ( .A1(n407), .A2(n2771), .B1(n359), .B2(n2770), .ZN(n2244) );
  OAI22_X2 U1982 ( .A1(n2772), .A2(n407), .B1(n359), .B2(n2771), .ZN(n2245) );
  OAI22_X2 U1983 ( .A1(n2772), .A2(n359), .B1(n407), .B2(n2773), .ZN(n2246) );
  OAI22_X2 U1984 ( .A1(n407), .A2(n2774), .B1(n359), .B2(n2773), .ZN(n2247) );
  OAI22_X2 U1985 ( .A1(n2775), .A2(n407), .B1(n359), .B2(n2774), .ZN(n2248) );
  OAI22_X2 U1986 ( .A1(n2775), .A2(n359), .B1(n407), .B2(n2776), .ZN(n2249) );
  OAI22_X2 U1987 ( .A1(n407), .A2(n2777), .B1(n359), .B2(n2776), .ZN(n2250) );
  OAI22_X2 U1988 ( .A1(n2778), .A2(n407), .B1(n359), .B2(n2777), .ZN(n2251) );
  OAI22_X2 U1989 ( .A1(n2778), .A2(n359), .B1(n407), .B2(n2779), .ZN(n2252) );
  OAI22_X2 U1990 ( .A1(n407), .A2(n2780), .B1(n359), .B2(n2779), .ZN(n2253) );
  OAI22_X2 U1991 ( .A1(n2781), .A2(n407), .B1(n359), .B2(n2780), .ZN(n2254) );
  OAI22_X2 U1992 ( .A1(n2781), .A2(n359), .B1(n407), .B2(n2782), .ZN(n2255) );
  OAI22_X2 U1994 ( .A1(n2784), .A2(n407), .B1(n359), .B2(n2783), .ZN(n2257) );
  OAI22_X2 U1995 ( .A1(n2784), .A2(n359), .B1(n407), .B2(n2785), .ZN(n2258) );
  OAI22_X2 U1996 ( .A1(n407), .A2(n2786), .B1(n359), .B2(n2785), .ZN(n2259) );
  OAI22_X2 U1997 ( .A1(n2787), .A2(n407), .B1(n359), .B2(n2786), .ZN(n2260) );
  OAI22_X2 U1998 ( .A1(n2787), .A2(n359), .B1(n407), .B2(n2788), .ZN(n2261) );
  OAI22_X2 U1999 ( .A1(n407), .A2(n2789), .B1(n359), .B2(n2788), .ZN(n2262) );
  OAI22_X2 U2000 ( .A1(n2790), .A2(n407), .B1(n359), .B2(n2789), .ZN(n2263) );
  OAI22_X2 U2001 ( .A1(n2790), .A2(n359), .B1(n407), .B2(n2791), .ZN(n2264) );
  OAI22_X2 U2002 ( .A1(n407), .A2(n2792), .B1(n359), .B2(n2791), .ZN(n2265) );
  OAI22_X2 U2003 ( .A1(n2793), .A2(n407), .B1(n359), .B2(n2792), .ZN(n2266) );
  OAI22_X2 U2004 ( .A1(n2793), .A2(n359), .B1(n407), .B2(n2794), .ZN(n2267) );
  OAI22_X2 U2005 ( .A1(n407), .A2(n2795), .B1(n359), .B2(n2794), .ZN(n2268) );
  OAI22_X2 U2038 ( .A1(n404), .A2(n3021), .B1(n3231), .B2(n2829), .ZN(n1885)
         );
  OAI22_X2 U2039 ( .A1(n2797), .A2(n3231), .B1(n404), .B2(n2798), .ZN(n2271)
         );
  OAI22_X2 U2040 ( .A1(n2799), .A2(n404), .B1(n3231), .B2(n2798), .ZN(n2272)
         );
  OAI22_X2 U2041 ( .A1(n2799), .A2(n3231), .B1(n404), .B2(n2800), .ZN(n2273)
         );
  OAI22_X2 U2042 ( .A1(n404), .A2(n2801), .B1(n3231), .B2(n2800), .ZN(n2274)
         );
  OAI22_X2 U2043 ( .A1(n2802), .A2(n404), .B1(n3231), .B2(n2801), .ZN(n2275)
         );
  OAI22_X2 U2044 ( .A1(n2802), .A2(n3231), .B1(n404), .B2(n2803), .ZN(n2276)
         );
  OAI22_X2 U2045 ( .A1(n404), .A2(n2804), .B1(n3231), .B2(n2803), .ZN(n2277)
         );
  OAI22_X2 U2046 ( .A1(n2805), .A2(n404), .B1(n3231), .B2(n2804), .ZN(n2278)
         );
  OAI22_X2 U2047 ( .A1(n2805), .A2(n3231), .B1(n404), .B2(n2806), .ZN(n2279)
         );
  OAI22_X2 U2048 ( .A1(n404), .A2(n2807), .B1(n3231), .B2(n2806), .ZN(n2280)
         );
  OAI22_X2 U2049 ( .A1(n2808), .A2(n404), .B1(n3231), .B2(n2807), .ZN(n2281)
         );
  OAI22_X2 U2050 ( .A1(n2808), .A2(n3231), .B1(n404), .B2(n2809), .ZN(n2282)
         );
  OAI22_X2 U2051 ( .A1(n404), .A2(n2810), .B1(n3231), .B2(n2809), .ZN(n2283)
         );
  OAI22_X2 U2052 ( .A1(n2811), .A2(n404), .B1(n3231), .B2(n2810), .ZN(n2284)
         );
  OAI22_X2 U2053 ( .A1(n2811), .A2(n3231), .B1(n404), .B2(n2812), .ZN(n2285)
         );
  OAI22_X2 U2054 ( .A1(n404), .A2(n2813), .B1(n3231), .B2(n2812), .ZN(n2286)
         );
  OAI22_X2 U2055 ( .A1(n2814), .A2(n404), .B1(n3231), .B2(n2813), .ZN(n2287)
         );
  OAI22_X2 U2056 ( .A1(n2814), .A2(n3231), .B1(n404), .B2(n2815), .ZN(n2288)
         );
  OAI22_X2 U2057 ( .A1(n404), .A2(n2816), .B1(n3231), .B2(n2815), .ZN(n2289)
         );
  OAI22_X2 U2058 ( .A1(n2817), .A2(n404), .B1(n3231), .B2(n2816), .ZN(n2290)
         );
  OAI22_X2 U2059 ( .A1(n2817), .A2(n3231), .B1(n404), .B2(n2818), .ZN(n2291)
         );
  OAI22_X2 U2060 ( .A1(n404), .A2(n2819), .B1(n3231), .B2(n2818), .ZN(n2292)
         );
  OAI22_X2 U2061 ( .A1(n2820), .A2(n404), .B1(n3231), .B2(n2819), .ZN(n2293)
         );
  OAI22_X2 U2062 ( .A1(n2820), .A2(n3231), .B1(n404), .B2(n2821), .ZN(n2294)
         );
  OAI22_X2 U2063 ( .A1(n404), .A2(n2822), .B1(n3231), .B2(n2821), .ZN(n2295)
         );
  OAI22_X2 U2064 ( .A1(n2823), .A2(n404), .B1(n3231), .B2(n2822), .ZN(n2296)
         );
  OAI22_X2 U2065 ( .A1(n2823), .A2(n3231), .B1(n404), .B2(n2824), .ZN(n2297)
         );
  OAI22_X2 U2066 ( .A1(n404), .A2(n2825), .B1(n3231), .B2(n2824), .ZN(n2298)
         );
  OAI22_X2 U2067 ( .A1(n2826), .A2(n404), .B1(n3231), .B2(n2825), .ZN(n2299)
         );
  OAI22_X2 U2068 ( .A1(n2826), .A2(n3231), .B1(n404), .B2(n2827), .ZN(n2300)
         );
  OAI22_X2 U2069 ( .A1(n404), .A2(n2828), .B1(n3231), .B2(n2827), .ZN(n2301)
         );
  OAI22_X2 U2102 ( .A1(n401), .A2(n3022), .B1(n3227), .B2(n2862), .ZN(n1886)
         );
  OAI22_X2 U2103 ( .A1(n2830), .A2(n3226), .B1(n401), .B2(n2831), .ZN(n2304)
         );
  OAI22_X2 U2104 ( .A1(n2832), .A2(n401), .B1(n2831), .B2(n3227), .ZN(n2305)
         );
  OAI22_X2 U2105 ( .A1(n2832), .A2(n3227), .B1(n401), .B2(n2833), .ZN(n2306)
         );
  OAI22_X2 U2106 ( .A1(n401), .A2(n2834), .B1(n2833), .B2(n3226), .ZN(n2307)
         );
  OAI22_X2 U2107 ( .A1(n2835), .A2(n401), .B1(n2834), .B2(n3226), .ZN(n2308)
         );
  OAI22_X2 U2108 ( .A1(n2835), .A2(n3226), .B1(n401), .B2(n2836), .ZN(n2309)
         );
  OAI22_X2 U2109 ( .A1(n401), .A2(n2837), .B1(n2836), .B2(n3226), .ZN(n2310)
         );
  OAI22_X2 U2110 ( .A1(n2838), .A2(n401), .B1(n2837), .B2(n3226), .ZN(n2311)
         );
  OAI22_X2 U2111 ( .A1(n2838), .A2(n3226), .B1(n401), .B2(n2839), .ZN(n2312)
         );
  OAI22_X2 U2112 ( .A1(n401), .A2(n2840), .B1(n2839), .B2(n3226), .ZN(n2313)
         );
  OAI22_X2 U2113 ( .A1(n2841), .A2(n401), .B1(n2840), .B2(n3226), .ZN(n2314)
         );
  OAI22_X2 U2114 ( .A1(n2841), .A2(n3227), .B1(n401), .B2(n2842), .ZN(n2315)
         );
  OAI22_X2 U2116 ( .A1(n2844), .A2(n401), .B1(n2843), .B2(n3227), .ZN(n2317)
         );
  OAI22_X2 U2117 ( .A1(n2844), .A2(n3226), .B1(n401), .B2(n2845), .ZN(n2318)
         );
  OAI22_X2 U2118 ( .A1(n401), .A2(n2846), .B1(n2845), .B2(n3227), .ZN(n2319)
         );
  OAI22_X2 U2119 ( .A1(n2847), .A2(n401), .B1(n2846), .B2(n3227), .ZN(n2320)
         );
  OAI22_X2 U2120 ( .A1(n2847), .A2(n3226), .B1(n401), .B2(n2848), .ZN(n2321)
         );
  OAI22_X2 U2121 ( .A1(n401), .A2(n2849), .B1(n2848), .B2(n3226), .ZN(n2322)
         );
  OAI22_X2 U2122 ( .A1(n2850), .A2(n401), .B1(n2849), .B2(n3226), .ZN(n2323)
         );
  OAI22_X2 U2123 ( .A1(n2850), .A2(n3227), .B1(n401), .B2(n2851), .ZN(n2324)
         );
  OAI22_X2 U2124 ( .A1(n401), .A2(n2852), .B1(n2851), .B2(n3227), .ZN(n2325)
         );
  OAI22_X2 U2125 ( .A1(n2853), .A2(n401), .B1(n2852), .B2(n3227), .ZN(n2326)
         );
  OAI22_X2 U2126 ( .A1(n2853), .A2(n3227), .B1(n401), .B2(n2854), .ZN(n2327)
         );
  OAI22_X2 U2127 ( .A1(n401), .A2(n2855), .B1(n2854), .B2(n3227), .ZN(n2328)
         );
  OAI22_X2 U2128 ( .A1(n2856), .A2(n401), .B1(n2855), .B2(n3227), .ZN(n2329)
         );
  OAI22_X2 U2129 ( .A1(n2856), .A2(n3227), .B1(n401), .B2(n2857), .ZN(n2330)
         );
  OAI22_X2 U2130 ( .A1(n401), .A2(n2858), .B1(n2857), .B2(n3226), .ZN(n2331)
         );
  OAI22_X2 U2131 ( .A1(n2859), .A2(n401), .B1(n2858), .B2(n3226), .ZN(n2332)
         );
  OAI22_X2 U2132 ( .A1(n2859), .A2(n3227), .B1(n401), .B2(n2860), .ZN(n2333)
         );
  OAI22_X2 U2133 ( .A1(n401), .A2(n2861), .B1(n2860), .B2(n3227), .ZN(n2334)
         );
  OAI22_X2 U2166 ( .A1(n398), .A2(n3023), .B1(n350), .B2(n2895), .ZN(n1887) );
  OAI22_X2 U2167 ( .A1(n2863), .A2(n350), .B1(n398), .B2(n2864), .ZN(n2337) );
  OAI22_X2 U2168 ( .A1(n2865), .A2(n398), .B1(n350), .B2(n2864), .ZN(n2338) );
  OAI22_X2 U2169 ( .A1(n2865), .A2(n350), .B1(n398), .B2(n2866), .ZN(n2339) );
  OAI22_X2 U2170 ( .A1(n398), .A2(n2867), .B1(n350), .B2(n2866), .ZN(n2340) );
  OAI22_X2 U2171 ( .A1(n2868), .A2(n398), .B1(n350), .B2(n2867), .ZN(n2341) );
  OAI22_X2 U2172 ( .A1(n2868), .A2(n350), .B1(n398), .B2(n2869), .ZN(n2342) );
  OAI22_X2 U2173 ( .A1(n398), .A2(n2870), .B1(n350), .B2(n2869), .ZN(n2343) );
  OAI22_X2 U2174 ( .A1(n2871), .A2(n398), .B1(n350), .B2(n2870), .ZN(n2344) );
  OAI22_X2 U2175 ( .A1(n2871), .A2(n350), .B1(n398), .B2(n2872), .ZN(n2345) );
  OAI22_X2 U2176 ( .A1(n398), .A2(n2873), .B1(n350), .B2(n2872), .ZN(n2346) );
  OAI22_X2 U2177 ( .A1(n2874), .A2(n398), .B1(n350), .B2(n2873), .ZN(n2347) );
  OAI22_X2 U2178 ( .A1(n2874), .A2(n350), .B1(n398), .B2(n2875), .ZN(n2348) );
  OAI22_X2 U2180 ( .A1(n2877), .A2(n398), .B1(n350), .B2(n2876), .ZN(n2350) );
  OAI22_X2 U2181 ( .A1(n2877), .A2(n350), .B1(n398), .B2(n2878), .ZN(n2351) );
  OAI22_X2 U2182 ( .A1(n398), .A2(n2879), .B1(n350), .B2(n2878), .ZN(n2352) );
  OAI22_X2 U2183 ( .A1(n2880), .A2(n398), .B1(n350), .B2(n2879), .ZN(n2353) );
  OAI22_X2 U2184 ( .A1(n2880), .A2(n350), .B1(n398), .B2(n2881), .ZN(n2354) );
  OAI22_X2 U2185 ( .A1(n398), .A2(n2882), .B1(n350), .B2(n2881), .ZN(n2355) );
  OAI22_X2 U2186 ( .A1(n2883), .A2(n398), .B1(n350), .B2(n2882), .ZN(n2356) );
  OAI22_X2 U2187 ( .A1(n2883), .A2(n350), .B1(n398), .B2(n2884), .ZN(n2357) );
  OAI22_X2 U2188 ( .A1(n398), .A2(n2885), .B1(n350), .B2(n2884), .ZN(n2358) );
  OAI22_X2 U2189 ( .A1(n2886), .A2(n398), .B1(n350), .B2(n2885), .ZN(n2359) );
  OAI22_X2 U2190 ( .A1(n2886), .A2(n350), .B1(n398), .B2(n2887), .ZN(n2360) );
  OAI22_X2 U2191 ( .A1(n398), .A2(n2888), .B1(n350), .B2(n2887), .ZN(n2361) );
  OAI22_X2 U2192 ( .A1(n2889), .A2(n398), .B1(n350), .B2(n2888), .ZN(n2362) );
  OAI22_X2 U2193 ( .A1(n2889), .A2(n350), .B1(n398), .B2(n2890), .ZN(n2363) );
  OAI22_X2 U2194 ( .A1(n398), .A2(n2891), .B1(n350), .B2(n2890), .ZN(n2364) );
  OAI22_X2 U2195 ( .A1(n2892), .A2(n398), .B1(n350), .B2(n2891), .ZN(n2365) );
  OAI22_X2 U2196 ( .A1(n2892), .A2(n350), .B1(n398), .B2(n2893), .ZN(n2366) );
  OAI22_X2 U2197 ( .A1(n398), .A2(n2894), .B1(n350), .B2(n2893), .ZN(n2367) );
  OAI22_X2 U2230 ( .A1(n395), .A2(n3024), .B1(n2928), .B2(n347), .ZN(n1888) );
  OAI22_X2 U2231 ( .A1(n2896), .A2(n347), .B1(n395), .B2(n2897), .ZN(n2370) );
  OAI22_X2 U2232 ( .A1(n2898), .A2(n395), .B1(n2897), .B2(n347), .ZN(n2371) );
  OAI22_X2 U2233 ( .A1(n2898), .A2(n347), .B1(n395), .B2(n2899), .ZN(n2372) );
  OAI22_X2 U2234 ( .A1(n395), .A2(n2900), .B1(n2899), .B2(n347), .ZN(n2373) );
  OAI22_X2 U2235 ( .A1(n2901), .A2(n395), .B1(n2900), .B2(n347), .ZN(n2374) );
  OAI22_X2 U2236 ( .A1(n2901), .A2(n347), .B1(n395), .B2(n2902), .ZN(n2375) );
  OAI22_X2 U2237 ( .A1(n395), .A2(n2903), .B1(n2902), .B2(n347), .ZN(n2376) );
  OAI22_X2 U2238 ( .A1(n2904), .A2(n395), .B1(n2903), .B2(n347), .ZN(n2377) );
  OAI22_X2 U2239 ( .A1(n2904), .A2(n347), .B1(n395), .B2(n2905), .ZN(n2378) );
  OAI22_X2 U2240 ( .A1(n395), .A2(n2906), .B1(n2905), .B2(n347), .ZN(n2379) );
  OAI22_X2 U2241 ( .A1(n2907), .A2(n395), .B1(n2906), .B2(n347), .ZN(n2380) );
  OAI22_X2 U2242 ( .A1(n2907), .A2(n347), .B1(n395), .B2(n2908), .ZN(n2381) );
  OAI22_X2 U2243 ( .A1(n395), .A2(n2909), .B1(n2908), .B2(n347), .ZN(n2382) );
  OAI22_X2 U2244 ( .A1(n2910), .A2(n395), .B1(n2909), .B2(n347), .ZN(n2383) );
  OAI22_X2 U2245 ( .A1(n2910), .A2(n347), .B1(n395), .B2(n2911), .ZN(n2384) );
  OAI22_X2 U2246 ( .A1(n395), .A2(n2912), .B1(n2911), .B2(n347), .ZN(n2385) );
  OAI22_X2 U2247 ( .A1(n2913), .A2(n395), .B1(n2912), .B2(n347), .ZN(n2386) );
  OAI22_X2 U2248 ( .A1(n2913), .A2(n347), .B1(n395), .B2(n2914), .ZN(n2387) );
  OAI22_X2 U2249 ( .A1(n395), .A2(n2915), .B1(n2914), .B2(n347), .ZN(n2388) );
  OAI22_X2 U2250 ( .A1(n2916), .A2(n395), .B1(n2915), .B2(n347), .ZN(n2389) );
  OAI22_X2 U2251 ( .A1(n2916), .A2(n347), .B1(n395), .B2(n2917), .ZN(n2390) );
  OAI22_X2 U2252 ( .A1(n395), .A2(n2918), .B1(n2917), .B2(n347), .ZN(n2391) );
  OAI22_X2 U2253 ( .A1(n2919), .A2(n395), .B1(n2918), .B2(n347), .ZN(n2392) );
  OAI22_X2 U2254 ( .A1(n2919), .A2(n347), .B1(n395), .B2(n2920), .ZN(n2393) );
  OAI22_X2 U2255 ( .A1(n395), .A2(n2921), .B1(n2920), .B2(n347), .ZN(n2394) );
  OAI22_X2 U2256 ( .A1(n2922), .A2(n395), .B1(n2921), .B2(n347), .ZN(n2395) );
  OAI22_X2 U2257 ( .A1(n2922), .A2(n347), .B1(n395), .B2(n2923), .ZN(n2396) );
  OAI22_X2 U2258 ( .A1(n395), .A2(n2924), .B1(n2923), .B2(n347), .ZN(n2397) );
  OAI22_X2 U2259 ( .A1(n2925), .A2(n395), .B1(n2924), .B2(n347), .ZN(n2398) );
  OAI22_X2 U2260 ( .A1(n2925), .A2(n347), .B1(n395), .B2(n2926), .ZN(n2399) );
  OAI22_X2 U2261 ( .A1(n395), .A2(n2927), .B1(n2926), .B2(n347), .ZN(n2400) );
  NAND2_X4 U2356 ( .A1(n2961), .A2(n3185), .ZN(n440) );
  XOR2_X2 U2357 ( .A(n342), .B(b[30]), .Z(n2961) );
  NAND2_X4 U2365 ( .A1(n2964), .A2(n3211), .ZN(n431) );
  XOR2_X2 U2366 ( .A(b[24]), .B(n335), .Z(n2964) );
  XOR2_X2 U2378 ( .A(b[16]), .B(n323), .Z(n2968) );
  NAND2_X4 U2383 ( .A1(n2970), .A2(n365), .ZN(n413) );
  XOR2_X2 U2384 ( .A(n317), .B(b[12]), .Z(n2970) );
  XOR2_X2 U2387 ( .A(b[10]), .B(n314), .Z(n2971) );
  NAND2_X4 U2392 ( .A1(n2973), .A2(n3230), .ZN(n404) );
  XOR2_X2 U2393 ( .A(b[6]), .B(n308), .Z(n2973) );
  XOR2_X2 U2396 ( .A(b[4]), .B(n305), .Z(n2974) );
  XOR2_X2 U2399 ( .A(b[2]), .B(n302), .Z(n2975) );
  NAND2_X4 U2401 ( .A1(n2976), .A2(n347), .ZN(n395) );
  XOR2_X2 U2402 ( .A(n299), .B(b[0]), .Z(n2976) );
  XNOR2_X1 U2406 ( .A(n342), .B(n2940), .ZN(n2412) );
  XNOR2_X1 U2407 ( .A(n2940), .B(n338), .ZN(n2478) );
  XNOR2_X1 U2408 ( .A(n2940), .B(n3173), .ZN(n2445) );
  XNOR2_X1 U2409 ( .A(n2940), .B(n323), .ZN(n2643) );
  XNOR2_X1 U2410 ( .A(n2940), .B(n320), .ZN(n2676) );
  XNOR2_X1 U2411 ( .A(n2940), .B(n326), .ZN(n2610) );
  XNOR2_X1 U2412 ( .A(n2940), .B(n305), .ZN(n2841) );
  XNOR2_X1 U2413 ( .A(n2940), .B(n329), .ZN(n2577) );
  XNOR2_X1 U2414 ( .A(n2940), .B(n335), .ZN(n2511) );
  XNOR2_X1 U2415 ( .A(n2940), .B(n332), .ZN(n2544) );
  XNOR2_X1 U2416 ( .A(n2940), .B(n314), .ZN(n2742) );
  XNOR2_X1 U2417 ( .A(n2940), .B(n317), .ZN(n2709) );
  XNOR2_X1 U2418 ( .A(n2940), .B(n302), .ZN(n2874) );
  XNOR2_X1 U2419 ( .A(n2940), .B(n308), .ZN(n2808) );
  XNOR2_X1 U2420 ( .A(n2940), .B(n311), .ZN(n2775) );
  XNOR2_X1 U2421 ( .A(n2940), .B(n3218), .ZN(n2907) );
  XNOR2_X1 U2422 ( .A(n2929), .B(n342), .ZN(n2401) );
  XNOR2_X1 U2423 ( .A(n2929), .B(n3173), .ZN(n2434) );
  XNOR2_X1 U2424 ( .A(n2929), .B(n338), .ZN(n2467) );
  XNOR2_X1 U2425 ( .A(n2929), .B(n335), .ZN(n2500) );
  XNOR2_X1 U2426 ( .A(n2929), .B(n332), .ZN(n2533) );
  XNOR2_X1 U2427 ( .A(n2929), .B(n329), .ZN(n2566) );
  XNOR2_X1 U2428 ( .A(n2929), .B(n326), .ZN(n2599) );
  XNOR2_X1 U2429 ( .A(n2929), .B(n317), .ZN(n2698) );
  XNOR2_X1 U2430 ( .A(n2929), .B(n320), .ZN(n2665) );
  XNOR2_X1 U2431 ( .A(n2929), .B(n305), .ZN(n2830) );
  XNOR2_X1 U2432 ( .A(n2929), .B(n323), .ZN(n2632) );
  XNOR2_X1 U2433 ( .A(n2929), .B(n302), .ZN(n2863) );
  XNOR2_X1 U2434 ( .A(n2929), .B(n314), .ZN(n2731) );
  XNOR2_X1 U2435 ( .A(n2929), .B(n311), .ZN(n2764) );
  XNOR2_X1 U2436 ( .A(n2929), .B(n308), .ZN(n2797) );
  XNOR2_X1 U2437 ( .A(n2929), .B(n3218), .ZN(n2896) );
  XNOR2_X1 U2438 ( .A(n342), .B(n2955), .ZN(n2427) );
  XNOR2_X1 U2439 ( .A(n2955), .B(n3218), .ZN(n2922) );
  XNOR2_X1 U2440 ( .A(n2955), .B(n302), .ZN(n2889) );
  XNOR2_X1 U2441 ( .A(n2955), .B(n305), .ZN(n2856) );
  XNOR2_X1 U2442 ( .A(n2955), .B(n338), .ZN(n2493) );
  XNOR2_X1 U2443 ( .A(n2955), .B(n311), .ZN(n2790) );
  XNOR2_X1 U2444 ( .A(n2955), .B(n329), .ZN(n2592) );
  XNOR2_X1 U2445 ( .A(n2955), .B(n341), .ZN(n2460) );
  XNOR2_X1 U2446 ( .A(n2955), .B(n308), .ZN(n2823) );
  XNOR2_X1 U2447 ( .A(n2955), .B(n332), .ZN(n2559) );
  XNOR2_X1 U2448 ( .A(n2955), .B(n323), .ZN(n2658) );
  XNOR2_X1 U2449 ( .A(n2955), .B(n317), .ZN(n2724) );
  XNOR2_X1 U2450 ( .A(n2955), .B(n326), .ZN(n2625) );
  XNOR2_X1 U2451 ( .A(n2955), .B(n335), .ZN(n2526) );
  XNOR2_X1 U2452 ( .A(n2955), .B(n314), .ZN(n2757) );
  XNOR2_X1 U2453 ( .A(n2955), .B(n320), .ZN(n2691) );
  XNOR2_X1 U2454 ( .A(n342), .B(n2934), .ZN(n2406) );
  XNOR2_X1 U2455 ( .A(n2934), .B(n3173), .ZN(n2439) );
  XNOR2_X1 U2456 ( .A(n2934), .B(n329), .ZN(n2571) );
  XNOR2_X1 U2457 ( .A(n2934), .B(n314), .ZN(n2736) );
  XNOR2_X1 U2458 ( .A(n2934), .B(n332), .ZN(n2538) );
  XNOR2_X1 U2459 ( .A(n2934), .B(n323), .ZN(n2637) );
  XNOR2_X1 U2460 ( .A(n2934), .B(n338), .ZN(n2472) );
  XNOR2_X1 U2461 ( .A(n2934), .B(n326), .ZN(n2604) );
  XNOR2_X1 U2462 ( .A(n2934), .B(n335), .ZN(n2505) );
  XNOR2_X1 U2463 ( .A(n2934), .B(n311), .ZN(n2769) );
  XNOR2_X1 U2464 ( .A(n2934), .B(n317), .ZN(n2703) );
  XNOR2_X1 U2465 ( .A(n2934), .B(n320), .ZN(n2670) );
  XNOR2_X1 U2466 ( .A(n2934), .B(n305), .ZN(n2835) );
  XNOR2_X1 U2467 ( .A(n2934), .B(n308), .ZN(n2802) );
  XNOR2_X1 U2468 ( .A(n2934), .B(n3218), .ZN(n2901) );
  XNOR2_X1 U2469 ( .A(n2934), .B(n302), .ZN(n2868) );
  XNOR2_X1 U2470 ( .A(n342), .B(n2937), .ZN(n2409) );
  XNOR2_X1 U2471 ( .A(n2937), .B(n320), .ZN(n2673) );
  XNOR2_X1 U2472 ( .A(n2937), .B(n338), .ZN(n2475) );
  XNOR2_X1 U2473 ( .A(n2937), .B(n317), .ZN(n2706) );
  XNOR2_X1 U2474 ( .A(n2937), .B(n335), .ZN(n2508) );
  XNOR2_X1 U2475 ( .A(n2937), .B(n3173), .ZN(n2442) );
  XNOR2_X1 U2476 ( .A(n2937), .B(n326), .ZN(n2607) );
  XNOR2_X1 U2477 ( .A(n2937), .B(n329), .ZN(n2574) );
  XNOR2_X1 U2478 ( .A(n2937), .B(n332), .ZN(n2541) );
  XNOR2_X1 U2479 ( .A(n2937), .B(n323), .ZN(n2640) );
  XNOR2_X1 U2480 ( .A(n2937), .B(n311), .ZN(n2772) );
  XNOR2_X1 U2481 ( .A(n2937), .B(n305), .ZN(n2838) );
  XNOR2_X1 U2482 ( .A(n2937), .B(n314), .ZN(n2739) );
  XNOR2_X1 U2483 ( .A(n2937), .B(n308), .ZN(n2805) );
  XNOR2_X1 U2484 ( .A(n2937), .B(n302), .ZN(n2871) );
  XNOR2_X1 U2485 ( .A(n2937), .B(n3218), .ZN(n2904) );
  XNOR2_X1 U2486 ( .A(n342), .B(n2946), .ZN(n2418) );
  XNOR2_X1 U2487 ( .A(n2946), .B(n335), .ZN(n2517) );
  XNOR2_X1 U2488 ( .A(n2946), .B(n332), .ZN(n2550) );
  XNOR2_X1 U2489 ( .A(n2946), .B(n3173), .ZN(n2451) );
  XNOR2_X1 U2490 ( .A(n2946), .B(n338), .ZN(n2484) );
  XNOR2_X1 U2491 ( .A(n2946), .B(n314), .ZN(n2748) );
  XNOR2_X1 U2492 ( .A(n2946), .B(n311), .ZN(n2781) );
  XNOR2_X1 U2493 ( .A(n2946), .B(n3218), .ZN(n2913) );
  XNOR2_X1 U2494 ( .A(n2946), .B(n317), .ZN(n2715) );
  XNOR2_X1 U2495 ( .A(n2946), .B(n320), .ZN(n2682) );
  XNOR2_X1 U2496 ( .A(n2946), .B(n329), .ZN(n2583) );
  XNOR2_X1 U2497 ( .A(n2946), .B(n326), .ZN(n2616) );
  XNOR2_X1 U2498 ( .A(n2946), .B(n302), .ZN(n2880) );
  XNOR2_X1 U2499 ( .A(n2946), .B(n305), .ZN(n2847) );
  XNOR2_X1 U2500 ( .A(n2946), .B(n308), .ZN(n2814) );
  XNOR2_X1 U2501 ( .A(n2946), .B(n323), .ZN(n2649) );
  XNOR2_X1 U2502 ( .A(n342), .B(n2949), .ZN(n2421) );
  XNOR2_X1 U2503 ( .A(n2949), .B(n335), .ZN(n2520) );
  XNOR2_X1 U2504 ( .A(n2949), .B(n338), .ZN(n2487) );
  XNOR2_X1 U2505 ( .A(n2949), .B(n3218), .ZN(n2916) );
  XNOR2_X1 U2506 ( .A(n2949), .B(n329), .ZN(n2586) );
  XNOR2_X1 U2507 ( .A(n2949), .B(n302), .ZN(n2883) );
  XNOR2_X1 U2508 ( .A(n2949), .B(n341), .ZN(n2454) );
  XNOR2_X1 U2509 ( .A(n2949), .B(n317), .ZN(n2718) );
  XNOR2_X1 U2510 ( .A(n2949), .B(n320), .ZN(n2685) );
  XNOR2_X1 U2511 ( .A(n2949), .B(n332), .ZN(n2553) );
  XNOR2_X1 U2512 ( .A(n2949), .B(n308), .ZN(n2817) );
  XNOR2_X1 U2513 ( .A(n2949), .B(n314), .ZN(n2751) );
  XNOR2_X1 U2514 ( .A(n2949), .B(n305), .ZN(n2850) );
  XNOR2_X1 U2515 ( .A(n2949), .B(n326), .ZN(n2619) );
  XNOR2_X1 U2516 ( .A(n2949), .B(n311), .ZN(n2784) );
  XNOR2_X1 U2517 ( .A(n2949), .B(n323), .ZN(n2652) );
  XNOR2_X1 U2518 ( .A(n342), .B(n2931), .ZN(n2403) );
  XNOR2_X1 U2519 ( .A(n2931), .B(n3173), .ZN(n2436) );
  XNOR2_X1 U2520 ( .A(n2931), .B(n338), .ZN(n2469) );
  XNOR2_X1 U2521 ( .A(n2931), .B(n332), .ZN(n2535) );
  XNOR2_X1 U2522 ( .A(n2931), .B(n335), .ZN(n2502) );
  XNOR2_X1 U2523 ( .A(n2931), .B(n323), .ZN(n2634) );
  XNOR2_X1 U2524 ( .A(n2931), .B(n326), .ZN(n2601) );
  XNOR2_X1 U2525 ( .A(n2931), .B(n329), .ZN(n2568) );
  XNOR2_X1 U2526 ( .A(n2931), .B(n311), .ZN(n2766) );
  XNOR2_X1 U2527 ( .A(n2931), .B(n314), .ZN(n2733) );
  XNOR2_X1 U2528 ( .A(n2931), .B(n308), .ZN(n2799) );
  XNOR2_X1 U2529 ( .A(n2931), .B(n320), .ZN(n2667) );
  XNOR2_X1 U2530 ( .A(n2931), .B(n317), .ZN(n2700) );
  XNOR2_X1 U2531 ( .A(n2931), .B(n302), .ZN(n2865) );
  XNOR2_X1 U2532 ( .A(n2931), .B(n305), .ZN(n2832) );
  XNOR2_X1 U2533 ( .A(n2931), .B(n3218), .ZN(n2898) );
  XNOR2_X1 U2534 ( .A(n2958), .B(n305), .ZN(n2859) );
  XNOR2_X1 U2535 ( .A(n2958), .B(n308), .ZN(n2826) );
  XNOR2_X1 U2536 ( .A(n2958), .B(n314), .ZN(n2760) );
  XNOR2_X1 U2537 ( .A(n2958), .B(n302), .ZN(n2892) );
  XNOR2_X1 U2538 ( .A(n2958), .B(n323), .ZN(n2661) );
  XNOR2_X1 U2539 ( .A(n2958), .B(n3218), .ZN(n2925) );
  XNOR2_X1 U2540 ( .A(n2958), .B(n311), .ZN(n2793) );
  XNOR2_X1 U2541 ( .A(n2958), .B(n332), .ZN(n2562) );
  XNOR2_X1 U2542 ( .A(n342), .B(n2958), .ZN(n2430) );
  XNOR2_X1 U2543 ( .A(n2958), .B(n320), .ZN(n2694) );
  XNOR2_X1 U2544 ( .A(n2958), .B(n329), .ZN(n2595) );
  XNOR2_X1 U2545 ( .A(n2958), .B(n341), .ZN(n2463) );
  XNOR2_X1 U2546 ( .A(n2958), .B(n326), .ZN(n2628) );
  XNOR2_X1 U2547 ( .A(n2958), .B(n317), .ZN(n2727) );
  XNOR2_X1 U2548 ( .A(n2958), .B(n338), .ZN(n2496) );
  XNOR2_X1 U2549 ( .A(n2958), .B(n335), .ZN(n2529) );
  XNOR2_X1 U2550 ( .A(n342), .B(n2952), .ZN(n2424) );
  XNOR2_X1 U2551 ( .A(n2952), .B(n3173), .ZN(n2457) );
  XNOR2_X1 U2552 ( .A(n2952), .B(n305), .ZN(n2853) );
  XNOR2_X1 U2553 ( .A(n2952), .B(n302), .ZN(n2886) );
  XNOR2_X1 U2554 ( .A(n2952), .B(n3218), .ZN(n2919) );
  XNOR2_X1 U2555 ( .A(n2952), .B(n332), .ZN(n2556) );
  XNOR2_X1 U2556 ( .A(n2952), .B(n323), .ZN(n2655) );
  XNOR2_X1 U2557 ( .A(n2952), .B(n308), .ZN(n2820) );
  XNOR2_X1 U2558 ( .A(n2952), .B(n329), .ZN(n2589) );
  XNOR2_X1 U2559 ( .A(n2952), .B(n338), .ZN(n2490) );
  XNOR2_X1 U2560 ( .A(n2952), .B(n311), .ZN(n2787) );
  XNOR2_X1 U2561 ( .A(n2952), .B(n335), .ZN(n2523) );
  XNOR2_X1 U2562 ( .A(n2952), .B(n320), .ZN(n2688) );
  XNOR2_X1 U2563 ( .A(n2952), .B(n314), .ZN(n2754) );
  XNOR2_X1 U2564 ( .A(n2952), .B(n326), .ZN(n2622) );
  XNOR2_X1 U2565 ( .A(n2952), .B(n317), .ZN(n2721) );
  XNOR2_X1 U2566 ( .A(n2943), .B(n3173), .ZN(n2448) );
  XNOR2_X1 U2567 ( .A(n342), .B(n2943), .ZN(n2415) );
  XNOR2_X1 U2568 ( .A(n2943), .B(n329), .ZN(n2580) );
  XNOR2_X1 U2569 ( .A(n2943), .B(n308), .ZN(n2811) );
  XNOR2_X1 U2570 ( .A(n2943), .B(n338), .ZN(n2481) );
  XNOR2_X1 U2571 ( .A(n2943), .B(n332), .ZN(n2547) );
  XNOR2_X1 U2572 ( .A(n2943), .B(n335), .ZN(n2514) );
  XNOR2_X1 U2573 ( .A(n2943), .B(n3218), .ZN(n2910) );
  XNOR2_X1 U2574 ( .A(n2943), .B(n320), .ZN(n2679) );
  XNOR2_X1 U2575 ( .A(n2943), .B(n317), .ZN(n2712) );
  XNOR2_X1 U2576 ( .A(n2943), .B(n326), .ZN(n2613) );
  XNOR2_X1 U2577 ( .A(n2943), .B(n302), .ZN(n2877) );
  XNOR2_X1 U2578 ( .A(n2943), .B(n311), .ZN(n2778) );
  XNOR2_X1 U2579 ( .A(n2943), .B(n314), .ZN(n2745) );
  XNOR2_X1 U2580 ( .A(n2943), .B(n323), .ZN(n2646) );
  XNOR2_X1 U2581 ( .A(n2943), .B(n305), .ZN(n2844) );
  XNOR2_X1 U2582 ( .A(n342), .B(n2954), .ZN(n2426) );
  XNOR2_X1 U2583 ( .A(n308), .B(n2954), .ZN(n2822) );
  XNOR2_X1 U2584 ( .A(n326), .B(n2954), .ZN(n2624) );
  XNOR2_X1 U2585 ( .A(n311), .B(n2954), .ZN(n2789) );
  XNOR2_X1 U2586 ( .A(n314), .B(n2954), .ZN(n2756) );
  XNOR2_X1 U2587 ( .A(n302), .B(n2954), .ZN(n2888) );
  XNOR2_X1 U2588 ( .A(n3218), .B(n2954), .ZN(n2921) );
  XNOR2_X1 U2589 ( .A(n305), .B(n2954), .ZN(n2855) );
  XNOR2_X1 U2590 ( .A(n320), .B(n2954), .ZN(n2690) );
  XNOR2_X1 U2591 ( .A(n335), .B(n2954), .ZN(n2525) );
  XNOR2_X1 U2592 ( .A(n338), .B(n2954), .ZN(n2492) );
  XNOR2_X1 U2593 ( .A(n332), .B(n2954), .ZN(n2558) );
  XNOR2_X1 U2594 ( .A(n329), .B(n2954), .ZN(n2591) );
  XNOR2_X1 U2595 ( .A(n323), .B(n2954), .ZN(n2657) );
  XNOR2_X1 U2596 ( .A(n317), .B(n2954), .ZN(n2723) );
  XNOR2_X1 U2597 ( .A(n342), .B(n2948), .ZN(n2420) );
  XNOR2_X1 U2598 ( .A(n332), .B(n2948), .ZN(n2552) );
  XNOR2_X1 U2599 ( .A(n326), .B(n2948), .ZN(n2618) );
  XNOR2_X1 U2600 ( .A(n308), .B(n2948), .ZN(n2816) );
  XNOR2_X1 U2601 ( .A(n320), .B(n2948), .ZN(n2684) );
  XNOR2_X1 U2602 ( .A(n3218), .B(n2948), .ZN(n2915) );
  XNOR2_X1 U2603 ( .A(n311), .B(n2948), .ZN(n2783) );
  XNOR2_X1 U2604 ( .A(n317), .B(n2948), .ZN(n2717) );
  XNOR2_X1 U2605 ( .A(n338), .B(n2948), .ZN(n2486) );
  XNOR2_X1 U2606 ( .A(n335), .B(n2948), .ZN(n2519) );
  XNOR2_X1 U2607 ( .A(n302), .B(n2948), .ZN(n2882) );
  XNOR2_X1 U2608 ( .A(n323), .B(n2948), .ZN(n2651) );
  XNOR2_X1 U2609 ( .A(n305), .B(n2948), .ZN(n2849) );
  XNOR2_X1 U2610 ( .A(n314), .B(n2948), .ZN(n2750) );
  XNOR2_X1 U2611 ( .A(n341), .B(n2948), .ZN(n2453) );
  XNOR2_X1 U2612 ( .A(n329), .B(n2948), .ZN(n2585) );
  XNOR2_X1 U2613 ( .A(n342), .B(n2947), .ZN(n2419) );
  XNOR2_X1 U2614 ( .A(n332), .B(n2947), .ZN(n2551) );
  XNOR2_X1 U2615 ( .A(n326), .B(n2947), .ZN(n2617) );
  XNOR2_X1 U2616 ( .A(n3218), .B(n2947), .ZN(n2914) );
  XNOR2_X1 U2617 ( .A(n308), .B(n2947), .ZN(n2815) );
  XNOR2_X1 U2618 ( .A(n338), .B(n2947), .ZN(n2485) );
  XNOR2_X1 U2619 ( .A(n320), .B(n2947), .ZN(n2683) );
  XNOR2_X1 U2620 ( .A(n311), .B(n2947), .ZN(n2782) );
  XNOR2_X1 U2621 ( .A(n317), .B(n2947), .ZN(n2716) );
  XNOR2_X1 U2622 ( .A(n335), .B(n2947), .ZN(n2518) );
  XNOR2_X1 U2623 ( .A(n302), .B(n2947), .ZN(n2881) );
  XNOR2_X1 U2624 ( .A(n305), .B(n2947), .ZN(n2848) );
  XNOR2_X1 U2625 ( .A(n323), .B(n2947), .ZN(n2650) );
  XNOR2_X1 U2626 ( .A(n314), .B(n2947), .ZN(n2749) );
  XNOR2_X1 U2627 ( .A(n341), .B(n2947), .ZN(n2452) );
  XNOR2_X1 U2628 ( .A(n329), .B(n2947), .ZN(n2584) );
  XNOR2_X1 U2629 ( .A(n342), .B(n2950), .ZN(n2422) );
  XNOR2_X1 U2630 ( .A(n338), .B(n2950), .ZN(n2488) );
  XNOR2_X1 U2631 ( .A(n341), .B(n2950), .ZN(n2455) );
  XNOR2_X1 U2632 ( .A(n323), .B(n2950), .ZN(n2653) );
  XNOR2_X1 U2633 ( .A(n311), .B(n2950), .ZN(n2785) );
  XNOR2_X1 U2634 ( .A(n3218), .B(n2950), .ZN(n2917) );
  XNOR2_X1 U2635 ( .A(n320), .B(n2950), .ZN(n2686) );
  XNOR2_X1 U2636 ( .A(n302), .B(n2950), .ZN(n2884) );
  XNOR2_X1 U2637 ( .A(n335), .B(n2950), .ZN(n2521) );
  XNOR2_X1 U2638 ( .A(n305), .B(n2950), .ZN(n2851) );
  XNOR2_X1 U2639 ( .A(n308), .B(n2950), .ZN(n2818) );
  XNOR2_X1 U2640 ( .A(n326), .B(n2950), .ZN(n2620) );
  XNOR2_X1 U2641 ( .A(n314), .B(n2950), .ZN(n2752) );
  XNOR2_X1 U2642 ( .A(n317), .B(n2950), .ZN(n2719) );
  XNOR2_X1 U2643 ( .A(n329), .B(n2950), .ZN(n2587) );
  XNOR2_X1 U2644 ( .A(n332), .B(n2950), .ZN(n2554) );
  XNOR2_X1 U2645 ( .A(n342), .B(n2951), .ZN(n2423) );
  XNOR2_X1 U2646 ( .A(n338), .B(n2951), .ZN(n2489) );
  XNOR2_X1 U2647 ( .A(n3173), .B(n2951), .ZN(n2456) );
  XNOR2_X1 U2648 ( .A(n311), .B(n2951), .ZN(n2786) );
  XNOR2_X1 U2649 ( .A(n323), .B(n2951), .ZN(n2654) );
  XNOR2_X1 U2650 ( .A(n3218), .B(n2951), .ZN(n2918) );
  XNOR2_X1 U2651 ( .A(n302), .B(n2951), .ZN(n2885) );
  XNOR2_X1 U2652 ( .A(n320), .B(n2951), .ZN(n2687) );
  XNOR2_X1 U2653 ( .A(n308), .B(n2951), .ZN(n2819) );
  XNOR2_X1 U2654 ( .A(n326), .B(n2951), .ZN(n2621) );
  XNOR2_X1 U2655 ( .A(n335), .B(n2951), .ZN(n2522) );
  XNOR2_X1 U2656 ( .A(n305), .B(n2951), .ZN(n2852) );
  XNOR2_X1 U2657 ( .A(n317), .B(n2951), .ZN(n2720) );
  XNOR2_X1 U2658 ( .A(n314), .B(n2951), .ZN(n2753) );
  XNOR2_X1 U2659 ( .A(n329), .B(n2951), .ZN(n2588) );
  XNOR2_X1 U2660 ( .A(n332), .B(n2951), .ZN(n2555) );
  XNOR2_X1 U2661 ( .A(n342), .B(n2945), .ZN(n2417) );
  XNOR2_X1 U2662 ( .A(n341), .B(n2945), .ZN(n2450) );
  XNOR2_X1 U2663 ( .A(n302), .B(n2945), .ZN(n2879) );
  XNOR2_X1 U2664 ( .A(n329), .B(n2945), .ZN(n2582) );
  XNOR2_X1 U2665 ( .A(n335), .B(n2945), .ZN(n2516) );
  XNOR2_X1 U2666 ( .A(n317), .B(n2945), .ZN(n2714) );
  XNOR2_X1 U2667 ( .A(n311), .B(n2945), .ZN(n2780) );
  XNOR2_X1 U2668 ( .A(n326), .B(n2945), .ZN(n2615) );
  XNOR2_X1 U2669 ( .A(n338), .B(n2945), .ZN(n2483) );
  XNOR2_X1 U2670 ( .A(n3218), .B(n2945), .ZN(n2912) );
  XNOR2_X1 U2671 ( .A(n332), .B(n2945), .ZN(n2549) );
  XNOR2_X1 U2672 ( .A(n308), .B(n2945), .ZN(n2813) );
  XNOR2_X1 U2673 ( .A(n323), .B(n2945), .ZN(n2648) );
  XNOR2_X1 U2674 ( .A(n320), .B(n2945), .ZN(n2681) );
  XNOR2_X1 U2675 ( .A(n314), .B(n2945), .ZN(n2747) );
  XNOR2_X1 U2676 ( .A(n305), .B(n2945), .ZN(n2846) );
  XNOR2_X1 U2677 ( .A(n342), .B(n2944), .ZN(n2416) );
  XNOR2_X1 U2678 ( .A(n341), .B(n2944), .ZN(n2449) );
  XNOR2_X1 U2679 ( .A(n335), .B(n2944), .ZN(n2515) );
  XNOR2_X1 U2680 ( .A(n311), .B(n2944), .ZN(n2779) );
  XNOR2_X1 U2681 ( .A(n338), .B(n2944), .ZN(n2482) );
  XNOR2_X1 U2682 ( .A(n302), .B(n2944), .ZN(n2878) );
  XNOR2_X1 U2683 ( .A(n317), .B(n2944), .ZN(n2713) );
  XNOR2_X1 U2684 ( .A(n329), .B(n2944), .ZN(n2581) );
  XNOR2_X1 U2685 ( .A(n332), .B(n2944), .ZN(n2548) );
  XNOR2_X1 U2686 ( .A(n3218), .B(n2944), .ZN(n2911) );
  XNOR2_X1 U2687 ( .A(n326), .B(n2944), .ZN(n2614) );
  XNOR2_X1 U2688 ( .A(n308), .B(n2944), .ZN(n2812) );
  XNOR2_X1 U2689 ( .A(n320), .B(n2944), .ZN(n2680) );
  XNOR2_X1 U2690 ( .A(n305), .B(n2944), .ZN(n2845) );
  XNOR2_X1 U2691 ( .A(n314), .B(n2944), .ZN(n2746) );
  XNOR2_X1 U2692 ( .A(n323), .B(n2944), .ZN(n2647) );
  XNOR2_X1 U2693 ( .A(n342), .B(n2953), .ZN(n2425) );
  XNOR2_X1 U2694 ( .A(n314), .B(n2953), .ZN(n2755) );
  XNOR2_X1 U2695 ( .A(n308), .B(n2953), .ZN(n2821) );
  XNOR2_X1 U2696 ( .A(n326), .B(n2953), .ZN(n2623) );
  XNOR2_X1 U2697 ( .A(n305), .B(n2953), .ZN(n2854) );
  XNOR2_X1 U2698 ( .A(n302), .B(n2953), .ZN(n2887) );
  XNOR2_X1 U2699 ( .A(n311), .B(n2953), .ZN(n2788) );
  XNOR2_X1 U2700 ( .A(n3218), .B(n2953), .ZN(n2920) );
  XNOR2_X1 U2701 ( .A(n335), .B(n2953), .ZN(n2524) );
  XNOR2_X1 U2702 ( .A(n320), .B(n2953), .ZN(n2689) );
  XNOR2_X1 U2703 ( .A(n332), .B(n2953), .ZN(n2557) );
  XNOR2_X1 U2704 ( .A(n341), .B(n2953), .ZN(n2458) );
  XNOR2_X1 U2705 ( .A(n338), .B(n2953), .ZN(n2491) );
  XNOR2_X1 U2706 ( .A(n323), .B(n2953), .ZN(n2656) );
  XNOR2_X1 U2707 ( .A(n329), .B(n2953), .ZN(n2590) );
  XNOR2_X1 U2708 ( .A(n317), .B(n2953), .ZN(n2722) );
  XNOR2_X1 U2709 ( .A(n342), .B(n2957), .ZN(n2429) );
  XNOR2_X1 U2710 ( .A(n3218), .B(n2957), .ZN(n2924) );
  XNOR2_X1 U2711 ( .A(n302), .B(n2957), .ZN(n2891) );
  XNOR2_X1 U2712 ( .A(n305), .B(n2957), .ZN(n2858) );
  XNOR2_X1 U2713 ( .A(n311), .B(n2957), .ZN(n2792) );
  XNOR2_X1 U2714 ( .A(n320), .B(n2957), .ZN(n2693) );
  XNOR2_X1 U2715 ( .A(n308), .B(n2957), .ZN(n2825) );
  XNOR2_X1 U2716 ( .A(n326), .B(n2957), .ZN(n2627) );
  XNOR2_X1 U2717 ( .A(n323), .B(n2957), .ZN(n2660) );
  XNOR2_X1 U2718 ( .A(n314), .B(n2957), .ZN(n2759) );
  XNOR2_X1 U2719 ( .A(n335), .B(n2957), .ZN(n2528) );
  XNOR2_X1 U2720 ( .A(n317), .B(n2957), .ZN(n2726) );
  XNOR2_X1 U2721 ( .A(n338), .B(n2957), .ZN(n2495) );
  XNOR2_X1 U2722 ( .A(n332), .B(n2957), .ZN(n2561) );
  XNOR2_X1 U2723 ( .A(n329), .B(n2957), .ZN(n2594) );
  XNOR2_X1 U2724 ( .A(n341), .B(n2957), .ZN(n2462) );
  XNOR2_X1 U2725 ( .A(n342), .B(n2942), .ZN(n2414) );
  XNOR2_X1 U2726 ( .A(n338), .B(n2942), .ZN(n2480) );
  XNOR2_X1 U2727 ( .A(n320), .B(n2942), .ZN(n2678) );
  XNOR2_X1 U2728 ( .A(n308), .B(n2942), .ZN(n2810) );
  XNOR2_X1 U2729 ( .A(n323), .B(n2942), .ZN(n2645) );
  XNOR2_X1 U2730 ( .A(n341), .B(n2942), .ZN(n2447) );
  XNOR2_X1 U2731 ( .A(n332), .B(n2942), .ZN(n2546) );
  XNOR2_X1 U2732 ( .A(n335), .B(n2942), .ZN(n2513) );
  XNOR2_X1 U2733 ( .A(n311), .B(n2942), .ZN(n2777) );
  XNOR2_X1 U2734 ( .A(n326), .B(n2942), .ZN(n2612) );
  XNOR2_X1 U2735 ( .A(n317), .B(n2942), .ZN(n2711) );
  XNOR2_X1 U2736 ( .A(n314), .B(n2942), .ZN(n2744) );
  XNOR2_X1 U2737 ( .A(n305), .B(n2942), .ZN(n2843) );
  XNOR2_X1 U2738 ( .A(n299), .B(n2942), .ZN(n2909) );
  XNOR2_X1 U2739 ( .A(n302), .B(n2942), .ZN(n2876) );
  XNOR2_X1 U2740 ( .A(n329), .B(n2942), .ZN(n2579) );
  XNOR2_X1 U2741 ( .A(n342), .B(n2941), .ZN(n2413) );
  XNOR2_X1 U2742 ( .A(n338), .B(n2941), .ZN(n2479) );
  XNOR2_X1 U2743 ( .A(n320), .B(n2941), .ZN(n2677) );
  XNOR2_X1 U2744 ( .A(n308), .B(n2941), .ZN(n2809) );
  XNOR2_X1 U2745 ( .A(n323), .B(n2941), .ZN(n2644) );
  XNOR2_X1 U2746 ( .A(n341), .B(n2941), .ZN(n2446) );
  XNOR2_X1 U2747 ( .A(n332), .B(n2941), .ZN(n2545) );
  XNOR2_X1 U2748 ( .A(n311), .B(n2941), .ZN(n2776) );
  XNOR2_X1 U2749 ( .A(n335), .B(n2941), .ZN(n2512) );
  XNOR2_X1 U2750 ( .A(n317), .B(n2941), .ZN(n2710) );
  XNOR2_X1 U2751 ( .A(n326), .B(n2941), .ZN(n2611) );
  XNOR2_X1 U2752 ( .A(n314), .B(n2941), .ZN(n2743) );
  XNOR2_X1 U2753 ( .A(n305), .B(n2941), .ZN(n2842) );
  XNOR2_X1 U2754 ( .A(n299), .B(n2941), .ZN(n2908) );
  XNOR2_X1 U2755 ( .A(n302), .B(n2941), .ZN(n2875) );
  XNOR2_X1 U2756 ( .A(n329), .B(n2941), .ZN(n2578) );
  XNOR2_X1 U2757 ( .A(n342), .B(n2933), .ZN(n2405) );
  XNOR2_X1 U2758 ( .A(n3173), .B(n2933), .ZN(n2438) );
  XNOR2_X1 U2759 ( .A(n338), .B(n2933), .ZN(n2471) );
  XNOR2_X1 U2760 ( .A(n335), .B(n2933), .ZN(n2504) );
  XNOR2_X1 U2761 ( .A(n323), .B(n2933), .ZN(n2636) );
  XNOR2_X1 U2762 ( .A(n332), .B(n2933), .ZN(n2537) );
  XNOR2_X1 U2763 ( .A(n308), .B(n2933), .ZN(n2801) );
  XNOR2_X1 U2764 ( .A(n329), .B(n2933), .ZN(n2570) );
  XNOR2_X1 U2765 ( .A(n311), .B(n2933), .ZN(n2768) );
  XNOR2_X1 U2766 ( .A(n320), .B(n2933), .ZN(n2669) );
  XNOR2_X1 U2767 ( .A(n326), .B(n2933), .ZN(n2603) );
  XNOR2_X1 U2768 ( .A(n317), .B(n2933), .ZN(n2702) );
  XNOR2_X1 U2769 ( .A(n3218), .B(n2933), .ZN(n2900) );
  XNOR2_X1 U2770 ( .A(n314), .B(n2933), .ZN(n2735) );
  XNOR2_X1 U2771 ( .A(n302), .B(n2933), .ZN(n2867) );
  XNOR2_X1 U2772 ( .A(n305), .B(n2933), .ZN(n2834) );
  XNOR2_X1 U2773 ( .A(n342), .B(n2956), .ZN(n2428) );
  XNOR2_X1 U2774 ( .A(n3218), .B(n2956), .ZN(n2923) );
  XNOR2_X1 U2775 ( .A(n305), .B(n2956), .ZN(n2857) );
  XNOR2_X1 U2776 ( .A(n302), .B(n2956), .ZN(n2890) );
  XNOR2_X1 U2777 ( .A(n326), .B(n2956), .ZN(n2626) );
  XNOR2_X1 U2778 ( .A(n308), .B(n2956), .ZN(n2824) );
  XNOR2_X1 U2779 ( .A(n311), .B(n2956), .ZN(n2791) );
  XNOR2_X1 U2780 ( .A(n320), .B(n2956), .ZN(n2692) );
  XNOR2_X1 U2781 ( .A(n314), .B(n2956), .ZN(n2758) );
  XNOR2_X1 U2782 ( .A(n317), .B(n2956), .ZN(n2725) );
  XNOR2_X1 U2783 ( .A(n323), .B(n2956), .ZN(n2659) );
  XNOR2_X1 U2784 ( .A(n335), .B(n2956), .ZN(n2527) );
  XNOR2_X1 U2785 ( .A(n332), .B(n2956), .ZN(n2560) );
  XNOR2_X1 U2786 ( .A(n329), .B(n2956), .ZN(n2593) );
  XNOR2_X1 U2787 ( .A(n338), .B(n2956), .ZN(n2494) );
  XNOR2_X1 U2788 ( .A(n341), .B(n2956), .ZN(n2461) );
  XNOR2_X1 U2789 ( .A(n342), .B(n2939), .ZN(n2411) );
  XNOR2_X1 U2790 ( .A(n323), .B(n2939), .ZN(n2642) );
  XNOR2_X1 U2791 ( .A(n341), .B(n2939), .ZN(n2444) );
  XNOR2_X1 U2792 ( .A(n332), .B(n2939), .ZN(n2543) );
  XNOR2_X1 U2793 ( .A(n326), .B(n2939), .ZN(n2609) );
  XNOR2_X1 U2794 ( .A(n338), .B(n2939), .ZN(n2477) );
  XNOR2_X1 U2795 ( .A(n320), .B(n2939), .ZN(n2675) );
  XNOR2_X1 U2796 ( .A(n308), .B(n2939), .ZN(n2807) );
  XNOR2_X1 U2797 ( .A(n317), .B(n2939), .ZN(n2708) );
  XNOR2_X1 U2798 ( .A(n335), .B(n2939), .ZN(n2510) );
  XNOR2_X1 U2799 ( .A(n329), .B(n2939), .ZN(n2576) );
  XNOR2_X1 U2800 ( .A(n299), .B(n2939), .ZN(n2906) );
  XNOR2_X1 U2801 ( .A(n311), .B(n2939), .ZN(n2774) );
  XNOR2_X1 U2802 ( .A(n302), .B(n2939), .ZN(n2873) );
  XNOR2_X1 U2803 ( .A(n305), .B(n2939), .ZN(n2840) );
  XNOR2_X1 U2804 ( .A(n314), .B(n2939), .ZN(n2741) );
  XNOR2_X1 U2805 ( .A(n342), .B(n2938), .ZN(n2410) );
  XNOR2_X1 U2806 ( .A(n323), .B(n2938), .ZN(n2641) );
  XNOR2_X1 U2807 ( .A(n332), .B(n2938), .ZN(n2542) );
  XNOR2_X1 U2808 ( .A(n341), .B(n2938), .ZN(n2443) );
  XNOR2_X1 U2809 ( .A(n338), .B(n2938), .ZN(n2476) );
  XNOR2_X1 U2810 ( .A(n326), .B(n2938), .ZN(n2608) );
  XNOR2_X1 U2811 ( .A(n320), .B(n2938), .ZN(n2674) );
  XNOR2_X1 U2812 ( .A(n329), .B(n2938), .ZN(n2575) );
  XNOR2_X1 U2813 ( .A(n335), .B(n2938), .ZN(n2509) );
  XNOR2_X1 U2814 ( .A(n317), .B(n2938), .ZN(n2707) );
  XNOR2_X1 U2815 ( .A(n308), .B(n2938), .ZN(n2806) );
  XNOR2_X1 U2816 ( .A(n311), .B(n2938), .ZN(n2773) );
  XNOR2_X1 U2817 ( .A(n302), .B(n2938), .ZN(n2872) );
  XNOR2_X1 U2818 ( .A(n299), .B(n2938), .ZN(n2905) );
  XNOR2_X1 U2819 ( .A(n305), .B(n2938), .ZN(n2839) );
  XNOR2_X1 U2820 ( .A(n314), .B(n2938), .ZN(n2740) );
  XNOR2_X1 U2821 ( .A(n342), .B(n2959), .ZN(n2431) );
  XNOR2_X1 U2822 ( .A(n3218), .B(n2959), .ZN(n2926) );
  XNOR2_X1 U2823 ( .A(n308), .B(n2959), .ZN(n2827) );
  XNOR2_X1 U2824 ( .A(n311), .B(n2959), .ZN(n2794) );
  XNOR2_X1 U2825 ( .A(n317), .B(n2959), .ZN(n2728) );
  XNOR2_X1 U2826 ( .A(n323), .B(n2959), .ZN(n2662) );
  XNOR2_X1 U2827 ( .A(n314), .B(n2959), .ZN(n2761) );
  XNOR2_X1 U2828 ( .A(n335), .B(n2959), .ZN(n2530) );
  XNOR2_X1 U2829 ( .A(n302), .B(n2959), .ZN(n2893) );
  XNOR2_X1 U2830 ( .A(n320), .B(n2959), .ZN(n2695) );
  XNOR2_X1 U2831 ( .A(n305), .B(n2959), .ZN(n2860) );
  XNOR2_X1 U2832 ( .A(n338), .B(n2959), .ZN(n2497) );
  XNOR2_X1 U2833 ( .A(n329), .B(n2959), .ZN(n2596) );
  XNOR2_X1 U2834 ( .A(n326), .B(n2959), .ZN(n2629) );
  XNOR2_X1 U2835 ( .A(n341), .B(n2959), .ZN(n2464) );
  XNOR2_X1 U2836 ( .A(n332), .B(n2959), .ZN(n2563) );
  XNOR2_X1 U2837 ( .A(n342), .B(n2932), .ZN(n2404) );
  XNOR2_X1 U2838 ( .A(n3173), .B(n2932), .ZN(n2437) );
  XNOR2_X1 U2839 ( .A(n338), .B(n2932), .ZN(n2470) );
  XNOR2_X1 U2840 ( .A(n335), .B(n2932), .ZN(n2503) );
  XNOR2_X1 U2841 ( .A(n323), .B(n2932), .ZN(n2635) );
  XNOR2_X1 U2842 ( .A(n332), .B(n2932), .ZN(n2536) );
  XNOR2_X1 U2843 ( .A(n308), .B(n2932), .ZN(n2800) );
  XNOR2_X1 U2844 ( .A(n329), .B(n2932), .ZN(n2569) );
  XNOR2_X1 U2845 ( .A(n320), .B(n2932), .ZN(n2668) );
  XNOR2_X1 U2846 ( .A(n317), .B(n2932), .ZN(n2701) );
  XNOR2_X1 U2847 ( .A(n311), .B(n2932), .ZN(n2767) );
  XNOR2_X1 U2848 ( .A(n3218), .B(n2932), .ZN(n2899) );
  XNOR2_X1 U2849 ( .A(n326), .B(n2932), .ZN(n2602) );
  XNOR2_X1 U2850 ( .A(n314), .B(n2932), .ZN(n2734) );
  XNOR2_X1 U2851 ( .A(n302), .B(n2932), .ZN(n2866) );
  XNOR2_X1 U2852 ( .A(n305), .B(n2932), .ZN(n2833) );
  XNOR2_X1 U2853 ( .A(n342), .B(n2936), .ZN(n2408) );
  XNOR2_X1 U2854 ( .A(n3173), .B(n2936), .ZN(n2441) );
  XNOR2_X1 U2855 ( .A(n332), .B(n2936), .ZN(n2540) );
  XNOR2_X1 U2856 ( .A(n314), .B(n2936), .ZN(n2738) );
  XNOR2_X1 U2857 ( .A(n326), .B(n2936), .ZN(n2606) );
  XNOR2_X1 U2858 ( .A(n335), .B(n2936), .ZN(n2507) );
  XNOR2_X1 U2859 ( .A(n305), .B(n2936), .ZN(n2837) );
  XNOR2_X1 U2860 ( .A(n338), .B(n2936), .ZN(n2474) );
  XNOR2_X1 U2861 ( .A(n323), .B(n2936), .ZN(n2639) );
  XNOR2_X1 U2862 ( .A(n320), .B(n2936), .ZN(n2672) );
  XNOR2_X1 U2863 ( .A(n311), .B(n2936), .ZN(n2771) );
  XNOR2_X1 U2864 ( .A(n3218), .B(n2936), .ZN(n2903) );
  XNOR2_X1 U2865 ( .A(n308), .B(n2936), .ZN(n2804) );
  XNOR2_X1 U2866 ( .A(n329), .B(n2936), .ZN(n2573) );
  XNOR2_X1 U2867 ( .A(n302), .B(n2936), .ZN(n2870) );
  XNOR2_X1 U2868 ( .A(n317), .B(n2936), .ZN(n2705) );
  XNOR2_X1 U2869 ( .A(n342), .B(n2935), .ZN(n2407) );
  XNOR2_X1 U2870 ( .A(n341), .B(n2935), .ZN(n2440) );
  XNOR2_X1 U2871 ( .A(n332), .B(n2935), .ZN(n2539) );
  XNOR2_X1 U2872 ( .A(n314), .B(n2935), .ZN(n2737) );
  XNOR2_X1 U2873 ( .A(n305), .B(n2935), .ZN(n2836) );
  XNOR2_X1 U2874 ( .A(n326), .B(n2935), .ZN(n2605) );
  XNOR2_X1 U2875 ( .A(n335), .B(n2935), .ZN(n2506) );
  XNOR2_X1 U2876 ( .A(n338), .B(n2935), .ZN(n2473) );
  XNOR2_X1 U2877 ( .A(n323), .B(n2935), .ZN(n2638) );
  XNOR2_X1 U2878 ( .A(n320), .B(n2935), .ZN(n2671) );
  XNOR2_X1 U2879 ( .A(n311), .B(n2935), .ZN(n2770) );
  XNOR2_X1 U2880 ( .A(n3218), .B(n2935), .ZN(n2902) );
  XNOR2_X1 U2881 ( .A(n329), .B(n2935), .ZN(n2572) );
  XNOR2_X1 U2882 ( .A(n308), .B(n2935), .ZN(n2803) );
  XNOR2_X1 U2883 ( .A(n302), .B(n2935), .ZN(n2869) );
  XNOR2_X1 U2884 ( .A(n317), .B(n2935), .ZN(n2704) );
  XNOR2_X1 U2885 ( .A(n342), .B(n2930), .ZN(n2402) );
  XNOR2_X1 U2886 ( .A(n3173), .B(n2930), .ZN(n2435) );
  XNOR2_X1 U2887 ( .A(n338), .B(n2930), .ZN(n2468) );
  XNOR2_X1 U2888 ( .A(n332), .B(n2930), .ZN(n2534) );
  XNOR2_X1 U2889 ( .A(n335), .B(n2930), .ZN(n2501) );
  XNOR2_X1 U2890 ( .A(n323), .B(n2930), .ZN(n2633) );
  XNOR2_X1 U2891 ( .A(n317), .B(n2930), .ZN(n2699) );
  XNOR2_X1 U2892 ( .A(n326), .B(n2930), .ZN(n2600) );
  XNOR2_X1 U2893 ( .A(n329), .B(n2930), .ZN(n2567) );
  XNOR2_X1 U2894 ( .A(n308), .B(n2930), .ZN(n2798) );
  XNOR2_X1 U2895 ( .A(n305), .B(n2930), .ZN(n2831) );
  XNOR2_X1 U2896 ( .A(n302), .B(n2930), .ZN(n2864) );
  XNOR2_X1 U2897 ( .A(n311), .B(n2930), .ZN(n2765) );
  XNOR2_X1 U2898 ( .A(n320), .B(n2930), .ZN(n2666) );
  XNOR2_X1 U2899 ( .A(n314), .B(n2930), .ZN(n2732) );
  XNOR2_X1 U2900 ( .A(n3218), .B(n2930), .ZN(n2897) );
  INV_X4 U2901 ( .A(b[0]), .ZN(n347) );
  NOR2_X1 U2902 ( .A1(n1482), .A2(n1509), .ZN(n724) );
  INV_X8 U2903 ( .A(n3263), .ZN(n365) );
  OAI21_X2 U2904 ( .B1(n699), .B2(n678), .A(n3172), .ZN(n677) );
  NAND2_X1 U2905 ( .A1(n1762), .A2(n1775), .ZN(n816) );
  OAI21_X1 U2906 ( .B1(n3284), .B2(n3263), .A(n3285), .ZN(n2172) );
  INV_X2 U2907 ( .A(n3265), .ZN(n353) );
  AND2_X2 U2908 ( .A1(n2965), .A2(n380), .ZN(n3171) );
  INV_X8 U2909 ( .A(n3171), .ZN(n428) );
  CLKBUF_X1 U2910 ( .A(n679), .Z(n3172) );
  INV_X4 U2911 ( .A(n3010), .ZN(n3173) );
  INV_X1 U2912 ( .A(n341), .ZN(n3010) );
  XOR2_X1 U2913 ( .A(n1262), .B(n1287), .Z(n3174) );
  XOR2_X1 U2914 ( .A(n1285), .B(n3174), .Z(n1258) );
  NAND2_X1 U2915 ( .A1(n1285), .A2(n1262), .ZN(n3175) );
  NAND2_X1 U2916 ( .A1(n1285), .A2(n1287), .ZN(n3176) );
  NAND2_X1 U2917 ( .A1(n1262), .A2(n1287), .ZN(n3177) );
  NAND3_X1 U2918 ( .A1(n3175), .A2(n3177), .A3(n3176), .ZN(n1257) );
  XOR2_X1 U2919 ( .A(n1563), .B(n1540), .Z(n3178) );
  XOR2_X1 U2920 ( .A(n1538), .B(n3178), .Z(n1536) );
  NAND2_X1 U2921 ( .A1(n1538), .A2(n1563), .ZN(n3179) );
  NAND2_X1 U2922 ( .A1(n1538), .A2(n1540), .ZN(n3180) );
  NAND2_X1 U2923 ( .A1(n1563), .A2(n1540), .ZN(n3181) );
  NAND3_X1 U2924 ( .A1(n3179), .A2(n3181), .A3(n3180), .ZN(n1535) );
  XOR2_X1 U2925 ( .A(n474), .B(n721), .Z(product[30]) );
  INV_X1 U2926 ( .A(n1183), .ZN(n1184) );
  NAND2_X1 U2927 ( .A1(n1072), .A2(n1087), .ZN(n619) );
  NAND2_X1 U2928 ( .A1(n1536), .A2(n1561), .ZN(n744) );
  BUF_X2 U2929 ( .A(n727), .Z(n3274) );
  NAND2_X1 U2930 ( .A1(n680), .A2(n692), .ZN(n678) );
  AOI21_X2 U2931 ( .B1(n670), .B2(n652), .A(n653), .ZN(n651) );
  INV_X1 U2932 ( .A(n700), .ZN(n699) );
  NOR2_X1 U2933 ( .A1(n687), .A2(n682), .ZN(n680) );
  NOR2_X2 U2934 ( .A1(n1282), .A2(n1307), .ZN(n682) );
  OAI22_X1 U2935 ( .A1(n428), .A2(n2555), .B1(n380), .B2(n2554), .ZN(n2032) );
  OAI21_X1 U2936 ( .B1(n671), .B2(n675), .A(n672), .ZN(n670) );
  INV_X4 U2937 ( .A(n437), .ZN(n3202) );
  XNOR2_X1 U2938 ( .A(n341), .B(n2954), .ZN(n2459) );
  NAND2_X2 U2939 ( .A1(n1256), .A2(n1281), .ZN(n675) );
  INV_X4 U2940 ( .A(n3228), .ZN(n3183) );
  INV_X2 U2941 ( .A(n3228), .ZN(n3182) );
  INV_X1 U2942 ( .A(n3228), .ZN(n410) );
  AND2_X1 U2943 ( .A1(n2971), .A2(n362), .ZN(n3228) );
  NOR2_X1 U2944 ( .A1(n1746), .A2(n1761), .ZN(n810) );
  NAND2_X1 U2945 ( .A1(n1746), .A2(n1761), .ZN(n811) );
  OAI21_X2 U2946 ( .B1(n785), .B2(n765), .A(n766), .ZN(n764) );
  XNOR2_X1 U2947 ( .A(n341), .B(n3247), .ZN(n3246) );
  INV_X1 U2948 ( .A(n3246), .ZN(n392) );
  OAI21_X1 U2949 ( .B1(n730), .B2(n747), .A(n731), .ZN(n729) );
  INV_X2 U2950 ( .A(n743), .ZN(n916) );
  INV_X2 U2951 ( .A(n392), .ZN(n3184) );
  INV_X1 U2952 ( .A(n3184), .ZN(n3185) );
  INV_X8 U2953 ( .A(n3184), .ZN(n3186) );
  NOR2_X1 U2954 ( .A1(n3185), .A2(n3275), .ZN(n1920) );
  INV_X1 U2955 ( .A(b[18]), .ZN(n3261) );
  XOR2_X1 U2956 ( .A(b[18]), .B(n326), .Z(n2967) );
  NOR2_X2 U2957 ( .A1(n654), .A2(n666), .ZN(n652) );
  NAND2_X1 U2958 ( .A1(n1164), .A2(n1185), .ZN(n659) );
  NOR2_X2 U2959 ( .A1(n1164), .A2(n1185), .ZN(n658) );
  NAND2_X1 U2960 ( .A1(n2962), .A2(n389), .ZN(n437) );
  INV_X1 U2961 ( .A(n1333), .ZN(n1334) );
  INV_X2 U2962 ( .A(n440), .ZN(n3187) );
  INV_X1 U2963 ( .A(n3187), .ZN(n3188) );
  INV_X4 U2964 ( .A(n3187), .ZN(n3190) );
  INV_X4 U2965 ( .A(n3187), .ZN(n3189) );
  OAI22_X1 U2966 ( .A1(n3205), .A2(n2462), .B1(n389), .B2(n2461), .ZN(n3191)
         );
  OR2_X1 U2967 ( .A1(n2122), .A2(n1943), .ZN(n1421) );
  OAI21_X1 U2968 ( .B1(n679), .B2(n650), .A(n651), .ZN(n649) );
  AOI21_X2 U2969 ( .B1(n680), .B2(n693), .A(n681), .ZN(n679) );
  AND2_X1 U2970 ( .A1(n441), .A2(b[0]), .ZN(product[0]) );
  XNOR2_X1 U2971 ( .A(n342), .B(n441), .ZN(n2432) );
  XNOR2_X1 U2972 ( .A(n3218), .B(n441), .ZN(n2927) );
  XNOR2_X1 U2973 ( .A(n308), .B(n441), .ZN(n2828) );
  XNOR2_X1 U2974 ( .A(n311), .B(n441), .ZN(n2795) );
  XNOR2_X1 U2975 ( .A(n317), .B(n441), .ZN(n2729) );
  XNOR2_X1 U2976 ( .A(n323), .B(n441), .ZN(n2663) );
  XNOR2_X1 U2977 ( .A(n314), .B(n441), .ZN(n2762) );
  XNOR2_X1 U2978 ( .A(n335), .B(n441), .ZN(n2531) );
  XNOR2_X1 U2979 ( .A(n302), .B(n441), .ZN(n2894) );
  XNOR2_X1 U2980 ( .A(n305), .B(n441), .ZN(n2861) );
  XNOR2_X1 U2981 ( .A(n338), .B(n441), .ZN(n2498) );
  XNOR2_X1 U2982 ( .A(n320), .B(n441), .ZN(n2696) );
  XNOR2_X1 U2983 ( .A(n326), .B(n441), .ZN(n2630) );
  XNOR2_X1 U2984 ( .A(n329), .B(n441), .ZN(n2597) );
  XNOR2_X1 U2985 ( .A(n341), .B(n441), .ZN(n2465) );
  XNOR2_X1 U2986 ( .A(n332), .B(n441), .ZN(n2564) );
  INV_X4 U2987 ( .A(n441), .ZN(n3275) );
  NAND2_X1 U2988 ( .A1(n1814), .A2(n1823), .ZN(n838) );
  NOR2_X1 U2989 ( .A1(n1814), .A2(n1823), .ZN(n837) );
  INV_X1 U2990 ( .A(b[20]), .ZN(n3271) );
  XOR2_X1 U2991 ( .A(b[20]), .B(n329), .Z(n2966) );
  OAI21_X1 U2992 ( .B1(n604), .B2(n598), .A(n599), .ZN(n597) );
  AOI21_X1 U2993 ( .B1(n515), .B2(n883), .A(n510), .ZN(n508) );
  INV_X1 U2994 ( .A(n598), .ZN(n895) );
  XOR2_X1 U2995 ( .A(n660), .B(n463), .Z(product[41]) );
  XOR2_X1 U2996 ( .A(n668), .B(n465), .Z(product[39]) );
  INV_X1 U2997 ( .A(n719), .ZN(n913) );
  OAI21_X2 U2998 ( .B1(n719), .B2(n725), .A(n720), .ZN(n718) );
  NAND2_X1 U2999 ( .A1(n1454), .A2(n1481), .ZN(n720) );
  NOR2_X2 U3000 ( .A1(n1454), .A2(n1481), .ZN(n719) );
  AOI21_X2 U3001 ( .B1(n902), .B2(n662), .A(n657), .ZN(n655) );
  INV_X1 U3002 ( .A(n659), .ZN(n657) );
  NAND2_X1 U3003 ( .A1(n903), .A2(n902), .ZN(n654) );
  XOR2_X1 U3004 ( .A(b[28]), .B(n341), .Z(n2962) );
  INV_X4 U3005 ( .A(b[28]), .ZN(n3252) );
  INV_X1 U3006 ( .A(b[22]), .ZN(n3267) );
  XOR2_X1 U3007 ( .A(b[22]), .B(n332), .Z(n2965) );
  XNOR2_X1 U3008 ( .A(n531), .B(n446), .ZN(product[58]) );
  OAI21_X1 U3009 ( .B1(n699), .B2(n697), .A(n698), .ZN(n696) );
  NAND2_X1 U3010 ( .A1(n910), .A2(n698), .ZN(n471) );
  AOI21_X1 U3011 ( .B1(n609), .B2(n542), .A(n543), .ZN(n541) );
  AOI21_X1 U3012 ( .B1(n609), .B2(n896), .A(n606), .ZN(n604) );
  INV_X1 U3013 ( .A(b[14]), .ZN(n3255) );
  XOR2_X1 U3014 ( .A(b[14]), .B(n320), .Z(n2969) );
  OAI22_X1 U3015 ( .A1(n422), .A2(n2624), .B1(n374), .B2(n2623), .ZN(n2098) );
  OAI22_X1 U3016 ( .A1(n2625), .A2(n374), .B1(n422), .B2(n2626), .ZN(n2100) );
  OAI22_X1 U3017 ( .A1(n2622), .A2(n422), .B1(n374), .B2(n2621), .ZN(n2096) );
  OAI22_X1 U3018 ( .A1(n422), .A2(n2609), .B1(n374), .B2(n2608), .ZN(n2083) );
  OAI22_X1 U3019 ( .A1(n422), .A2(n2630), .B1(n374), .B2(n2629), .ZN(n2104) );
  OAI22_X1 U3020 ( .A1(n422), .A2(n3015), .B1(n374), .B2(n2631), .ZN(n1879) );
  OAI22_X1 U3021 ( .A1(n422), .A2(n2615), .B1(n374), .B2(n2614), .ZN(n2089) );
  OAI22_X1 U3022 ( .A1(n422), .A2(n2603), .B1(n374), .B2(n2602), .ZN(n2077) );
  OAI22_X1 U3023 ( .A1(n422), .A2(n2612), .B1(n374), .B2(n2611), .ZN(n2086) );
  NOR2_X2 U3024 ( .A1(n1308), .A2(n1335), .ZN(n687) );
  INV_X4 U3025 ( .A(n3256), .ZN(n359) );
  XOR2_X1 U3026 ( .A(b[8]), .B(n311), .Z(n2972) );
  INV_X4 U3027 ( .A(b[8]), .ZN(n3257) );
  INV_X2 U3028 ( .A(n3260), .ZN(n3193) );
  INV_X2 U3029 ( .A(n3260), .ZN(n374) );
  AOI21_X1 U3030 ( .B1(n677), .B2(n669), .A(n670), .ZN(n668) );
  INV_X4 U3031 ( .A(n3249), .ZN(n386) );
  XOR2_X1 U3032 ( .A(b[26]), .B(n338), .Z(n2963) );
  INV_X4 U3033 ( .A(b[26]), .ZN(n3250) );
  INV_X1 U3034 ( .A(n666), .ZN(n904) );
  OAI21_X2 U3035 ( .B1(n668), .B2(n666), .A(n667), .ZN(n665) );
  NAND2_X2 U3036 ( .A1(n1208), .A2(n1231), .ZN(n667) );
  NOR2_X2 U3037 ( .A1(n1208), .A2(n1231), .ZN(n666) );
  XNOR2_X2 U3038 ( .A(n326), .B(n3271), .ZN(n3270) );
  NOR2_X1 U3039 ( .A1(n1336), .A2(n1363), .ZN(n3192) );
  NOR2_X1 U3040 ( .A1(n1336), .A2(n1363), .ZN(n694) );
  OAI21_X1 U3041 ( .B1(n694), .B2(n698), .A(n695), .ZN(n693) );
  OAI22_X1 U3042 ( .A1(n434), .A2(n2495), .B1(n386), .B2(n2494), .ZN(n1974) );
  OAI21_X2 U3043 ( .B1(n3274), .B2(n701), .A(n702), .ZN(n700) );
  AOI21_X2 U3044 ( .B1(n726), .B2(n914), .A(n723), .ZN(n721) );
  OAI22_X1 U3045 ( .A1(n3188), .A2(n2431), .B1(n2430), .B2(n3186), .ZN(n1918)
         );
  INV_X2 U3046 ( .A(n3206), .ZN(n3209) );
  INV_X1 U3047 ( .A(n682), .ZN(n907) );
  OAI21_X1 U3048 ( .B1(n682), .B2(n688), .A(n683), .ZN(n681) );
  OAI22_X1 U3049 ( .A1(n422), .A2(n2618), .B1(n374), .B2(n2617), .ZN(n2092) );
  OAI22_X1 U3050 ( .A1(n422), .A2(n2621), .B1(n374), .B2(n2620), .ZN(n2095) );
  OAI21_X1 U3051 ( .B1(n785), .B2(n765), .A(n766), .ZN(n3194) );
  NAND2_X2 U3052 ( .A1(n1042), .A2(n1055), .ZN(n599) );
  NOR2_X2 U3053 ( .A1(n1042), .A2(n1055), .ZN(n598) );
  OAI21_X1 U3054 ( .B1(n545), .B2(n525), .A(n526), .ZN(n524) );
  AOI21_X2 U3055 ( .B1(n613), .B2(n523), .A(n524), .ZN(n522) );
  OAI21_X1 U3056 ( .B1(n522), .B2(n516), .A(n517), .ZN(n515) );
  INV_X4 U3057 ( .A(n3268), .ZN(n362) );
  INV_X1 U3058 ( .A(b[10]), .ZN(n3269) );
  INV_X1 U3059 ( .A(b[12]), .ZN(n3264) );
  XOR2_X1 U3060 ( .A(n763), .B(n479), .Z(product[25]) );
  NAND2_X1 U3061 ( .A1(n903), .A2(n664), .ZN(n464) );
  AOI21_X1 U3062 ( .B1(n665), .B2(n903), .A(n662), .ZN(n660) );
  INV_X1 U3063 ( .A(n663), .ZN(n903) );
  OAI21_X1 U3064 ( .B1(n3273), .B2(n3249), .A(n3293), .ZN(n1948) );
  OAI21_X1 U3065 ( .B1(n3199), .B2(n3260), .A(n3288), .ZN(n2073) );
  XNOR2_X1 U3066 ( .A(n756), .B(n478), .ZN(product[26]) );
  OAI21_X1 U3067 ( .B1(n3201), .B2(n3256), .A(n3282), .ZN(n2237) );
  OAI21_X1 U3068 ( .B1(n654), .B2(n667), .A(n655), .ZN(n653) );
  AOI21_X2 U3069 ( .B1(n703), .B2(n718), .A(n704), .ZN(n702) );
  AOI21_X2 U3070 ( .B1(n915), .B2(n742), .A(n733), .ZN(n731) );
  INV_X1 U3071 ( .A(n744), .ZN(n742) );
  OAI22_X1 U3072 ( .A1(n407), .A2(n2783), .B1(n359), .B2(n2782), .ZN(n2256) );
  NAND2_X1 U3073 ( .A1(n1586), .A2(n1609), .ZN(n758) );
  INV_X1 U3074 ( .A(n758), .ZN(n760) );
  NAND2_X1 U3075 ( .A1(n918), .A2(n758), .ZN(n479) );
  OAI21_X1 U3076 ( .B1(n763), .B2(n757), .A(n758), .ZN(n756) );
  INV_X2 U3077 ( .A(n368), .ZN(n3195) );
  INV_X1 U3078 ( .A(n3195), .ZN(n3196) );
  INV_X8 U3079 ( .A(n3195), .ZN(n3198) );
  INV_X4 U3080 ( .A(n3195), .ZN(n3197) );
  OAI21_X1 U3081 ( .B1(n541), .B2(n539), .A(n540), .ZN(n538) );
  OAI21_X1 U3082 ( .B1(n541), .B2(n532), .A(n533), .ZN(n531) );
  XOR2_X1 U3083 ( .A(n541), .B(n448), .Z(product[56]) );
  NOR2_X2 U3084 ( .A1(n1364), .A2(n1393), .ZN(n697) );
  NAND2_X2 U3085 ( .A1(n1364), .A2(n1393), .ZN(n698) );
  OAI22_X1 U3086 ( .A1(n2434), .A2(n389), .B1(n3205), .B2(n2435), .ZN(n949) );
  OAI22_X1 U3087 ( .A1(n3205), .A2(n2438), .B1(n389), .B2(n2437), .ZN(n1923)
         );
  OAI22_X1 U3088 ( .A1(n2439), .A2(n3205), .B1(n389), .B2(n2438), .ZN(n1924)
         );
  OAI22_X1 U3089 ( .A1(n2442), .A2(n3205), .B1(n389), .B2(n2441), .ZN(n1926)
         );
  OAI22_X1 U3090 ( .A1(n3205), .A2(n2441), .B1(n389), .B2(n2440), .ZN(n991) );
  OAI22_X1 U3091 ( .A1(n2445), .A2(n389), .B1(n3205), .B2(n2446), .ZN(n1930)
         );
  OAI22_X1 U3092 ( .A1(n2445), .A2(n3205), .B1(n389), .B2(n2444), .ZN(n1929)
         );
  OAI22_X1 U3093 ( .A1(n2451), .A2(n3205), .B1(n389), .B2(n2450), .ZN(n1934)
         );
  OAI22_X1 U3094 ( .A1(n2454), .A2(n389), .B1(n3205), .B2(n2455), .ZN(n1937)
         );
  OAI22_X1 U3095 ( .A1(n3205), .A2(n2444), .B1(n389), .B2(n2443), .ZN(n1928)
         );
  OAI22_X1 U3096 ( .A1(n2454), .A2(n3205), .B1(n389), .B2(n2453), .ZN(n1936)
         );
  OAI22_X1 U3097 ( .A1(n2460), .A2(n3205), .B1(n389), .B2(n2459), .ZN(n1941)
         );
  OAI22_X1 U3098 ( .A1(n2460), .A2(n389), .B1(n3205), .B2(n2461), .ZN(n1942)
         );
  OAI22_X1 U3099 ( .A1(n3205), .A2(n2447), .B1(n389), .B2(n2446), .ZN(n1069)
         );
  OAI22_X1 U3100 ( .A1(n3205), .A2(n2465), .B1(n389), .B2(n2464), .ZN(n1946)
         );
  AND2_X2 U3101 ( .A1(n2967), .A2(n374), .ZN(n3199) );
  INV_X8 U3102 ( .A(n3199), .ZN(n422) );
  INV_X4 U3103 ( .A(n3254), .ZN(n368) );
  OAI21_X2 U3104 ( .B1(n806), .B2(n823), .A(n807), .ZN(n805) );
  INV_X1 U3105 ( .A(n3274), .ZN(n3200) );
  NAND2_X2 U3106 ( .A1(n915), .A2(n916), .ZN(n730) );
  INV_X1 U3107 ( .A(n3270), .ZN(n377) );
  OAI21_X1 U3108 ( .B1(n3236), .B2(n3270), .A(n3289), .ZN(n2043) );
  NAND2_X2 U3109 ( .A1(n1632), .A2(n1653), .ZN(n773) );
  AND2_X2 U3110 ( .A1(n2972), .A2(n359), .ZN(n3201) );
  INV_X8 U3111 ( .A(n3201), .ZN(n407) );
  NAND2_X1 U3112 ( .A1(n909), .A2(n695), .ZN(n470) );
  OAI21_X1 U3113 ( .B1(n3294), .B2(n3251), .A(n3295), .ZN(n1921) );
  INV_X1 U3114 ( .A(n671), .ZN(n905) );
  NOR2_X2 U3115 ( .A1(n674), .A2(n671), .ZN(n669) );
  NAND2_X2 U3116 ( .A1(n1232), .A2(n1255), .ZN(n672) );
  NOR2_X2 U3117 ( .A1(n1232), .A2(n1255), .ZN(n671) );
  INV_X1 U3118 ( .A(n693), .ZN(n691) );
  INV_X1 U3119 ( .A(n796), .ZN(n794) );
  NAND2_X1 U3120 ( .A1(n924), .A2(n796), .ZN(n485) );
  INV_X1 U3121 ( .A(n769), .ZN(n919) );
  INV_X1 U3122 ( .A(n3202), .ZN(n3203) );
  INV_X4 U3123 ( .A(n3202), .ZN(n3205) );
  INV_X4 U3124 ( .A(n3202), .ZN(n3204) );
  NAND2_X2 U3125 ( .A1(n1308), .A2(n1335), .ZN(n688) );
  XOR2_X1 U3126 ( .A(n3239), .B(n1564), .Z(n1562) );
  NAND2_X1 U3127 ( .A1(n1562), .A2(n1585), .ZN(n755) );
  NOR2_X1 U3128 ( .A1(n1562), .A2(n1585), .ZN(n754) );
  NAND2_X1 U3129 ( .A1(n915), .A2(n735), .ZN(n476) );
  OAI22_X1 U3130 ( .A1(n3182), .A2(n2747), .B1(n362), .B2(n2746), .ZN(n2220)
         );
  INV_X2 U3131 ( .A(n377), .ZN(n3206) );
  INV_X1 U3132 ( .A(n3206), .ZN(n3207) );
  INV_X2 U3133 ( .A(n3206), .ZN(n3208) );
  OAI21_X1 U3134 ( .B1(n3219), .B2(n3254), .A(n3286), .ZN(n2139) );
  INV_X1 U3135 ( .A(n727), .ZN(n726) );
  XNOR2_X1 U3136 ( .A(n625), .B(n459), .ZN(product[45]) );
  AOI21_X1 U3137 ( .B1(n625), .B2(n898), .A(n622), .ZN(n620) );
  INV_X1 U3138 ( .A(n3192), .ZN(n909) );
  NOR2_X1 U3139 ( .A1(n697), .A2(n3192), .ZN(n692) );
  NOR2_X1 U3140 ( .A1(n1186), .A2(n1207), .ZN(n663) );
  NAND2_X2 U3141 ( .A1(n1186), .A2(n1207), .ZN(n664) );
  INV_X1 U3142 ( .A(n1391), .ZN(n1392) );
  INV_X4 U3143 ( .A(n383), .ZN(n3210) );
  INV_X1 U3144 ( .A(n3210), .ZN(n3211) );
  INV_X2 U3145 ( .A(n3210), .ZN(n3213) );
  INV_X4 U3146 ( .A(n3210), .ZN(n3212) );
  NAND2_X1 U3147 ( .A1(b[2]), .A2(n3215), .ZN(n3216) );
  NAND2_X1 U3148 ( .A1(n3214), .A2(n299), .ZN(n3217) );
  NAND2_X2 U3149 ( .A1(n3216), .A2(n3217), .ZN(n3272) );
  INV_X1 U3150 ( .A(b[2]), .ZN(n3214) );
  INV_X1 U3151 ( .A(n299), .ZN(n3215) );
  INV_X8 U3152 ( .A(n3024), .ZN(n3218) );
  INV_X8 U3153 ( .A(n3272), .ZN(n350) );
  AND2_X2 U3154 ( .A1(n2969), .A2(n3196), .ZN(n3219) );
  INV_X8 U3155 ( .A(n3219), .ZN(n416) );
  NAND2_X1 U3156 ( .A1(n1282), .A2(n1307), .ZN(n683) );
  CLKBUF_X1 U3157 ( .A(n784), .Z(n3220) );
  AOI21_X1 U3158 ( .B1(n3200), .B2(n708), .A(n709), .ZN(n707) );
  XNOR2_X1 U3159 ( .A(n745), .B(n477), .ZN(product[27]) );
  INV_X2 U3160 ( .A(n413), .ZN(n3221) );
  INV_X1 U3161 ( .A(n3221), .ZN(n3222) );
  INV_X8 U3162 ( .A(n3221), .ZN(n3223) );
  INV_X1 U3163 ( .A(n3223), .ZN(n3284) );
  OAI21_X1 U3164 ( .B1(n3228), .B2(n3268), .A(n3283), .ZN(n2204) );
  NAND2_X1 U3165 ( .A1(n1336), .A2(n1363), .ZN(n695) );
  INV_X2 U3166 ( .A(n353), .ZN(n3224) );
  INV_X1 U3167 ( .A(n3224), .ZN(n3225) );
  INV_X4 U3168 ( .A(n3224), .ZN(n3227) );
  INV_X2 U3169 ( .A(n3224), .ZN(n3226) );
  AOI21_X1 U3170 ( .B1(n784), .B2(n922), .A(n781), .ZN(n779) );
  XNOR2_X1 U3171 ( .A(n3220), .B(n483), .ZN(product[21]) );
  INV_X2 U3172 ( .A(n356), .ZN(n3229) );
  INV_X1 U3173 ( .A(n3229), .ZN(n3230) );
  INV_X4 U3174 ( .A(n3229), .ZN(n3231) );
  XNOR2_X1 U3175 ( .A(n726), .B(n475), .ZN(product[29]) );
  INV_X4 U3176 ( .A(n371), .ZN(n3232) );
  INV_X1 U3177 ( .A(n3232), .ZN(n3233) );
  INV_X4 U3178 ( .A(n3232), .ZN(n3235) );
  INV_X2 U3179 ( .A(n3232), .ZN(n3234) );
  NOR2_X2 U3180 ( .A1(n1510), .A2(n1535), .ZN(n734) );
  OAI21_X1 U3181 ( .B1(n769), .B2(n773), .A(n770), .ZN(n768) );
  NOR2_X2 U3182 ( .A1(n772), .A2(n769), .ZN(n767) );
  AND2_X2 U3183 ( .A1(n2966), .A2(n3207), .ZN(n3236) );
  INV_X8 U3184 ( .A(n3236), .ZN(n425) );
  NOR2_X2 U3185 ( .A1(n1610), .A2(n1631), .ZN(n769) );
  NAND2_X2 U3186 ( .A1(n1610), .A2(n1631), .ZN(n770) );
  INV_X1 U3187 ( .A(n404), .ZN(n3280) );
  NOR2_X2 U3188 ( .A1(n1586), .A2(n1609), .ZN(n757) );
  OAI21_X1 U3189 ( .B1(n3248), .B2(n3272), .A(n3278), .ZN(n2336) );
  OAI21_X1 U3190 ( .B1(n3237), .B2(n3265), .A(n3279), .ZN(n2303) );
  AND2_X2 U3191 ( .A1(n2974), .A2(n3225), .ZN(n3237) );
  INV_X8 U3192 ( .A(n3237), .ZN(n401) );
  XOR2_X1 U3193 ( .A(n1589), .B(n1570), .Z(n3238) );
  XOR2_X1 U3194 ( .A(n3238), .B(n1568), .Z(n1564) );
  XOR2_X1 U3195 ( .A(n1587), .B(n1566), .Z(n3239) );
  NAND2_X1 U3196 ( .A1(n1589), .A2(n1570), .ZN(n3240) );
  NAND2_X1 U3197 ( .A1(n1589), .A2(n1568), .ZN(n3241) );
  NAND2_X1 U3198 ( .A1(n1570), .A2(n1568), .ZN(n3242) );
  NAND3_X1 U3199 ( .A1(n3240), .A2(n3241), .A3(n3242), .ZN(n1563) );
  NAND2_X1 U3200 ( .A1(n1587), .A2(n1566), .ZN(n3243) );
  NAND2_X1 U3201 ( .A1(n1587), .A2(n1564), .ZN(n3244) );
  NAND2_X1 U3202 ( .A1(n1566), .A2(n1564), .ZN(n3245) );
  NAND3_X1 U3203 ( .A1(n3243), .A2(n3244), .A3(n3245), .ZN(n1561) );
  NAND2_X1 U3204 ( .A1(n767), .A2(n775), .ZN(n765) );
  AOI21_X2 U3205 ( .B1(n767), .B2(n776), .A(n768), .ZN(n766) );
  INV_X32 U3206 ( .A(b[30]), .ZN(n3247) );
  INV_X1 U3207 ( .A(n3189), .ZN(n3296) );
  AND2_X2 U3208 ( .A1(n2975), .A2(n350), .ZN(n3248) );
  INV_X8 U3209 ( .A(n3248), .ZN(n398) );
  XNOR2_X2 U3210 ( .A(n335), .B(n3250), .ZN(n3249) );
  XNOR2_X2 U3211 ( .A(n3252), .B(n338), .ZN(n3251) );
  INV_X8 U3212 ( .A(n3251), .ZN(n389) );
  XOR2_X2 U3213 ( .A(b[16]), .B(n320), .Z(n3253) );
  INV_X4 U3214 ( .A(n3253), .ZN(n371) );
  XNOR2_X2 U3215 ( .A(n317), .B(n3255), .ZN(n3254) );
  XNOR2_X2 U3216 ( .A(n3257), .B(n308), .ZN(n3256) );
  XOR2_X2 U3217 ( .A(b[24]), .B(n332), .Z(n3258) );
  INV_X4 U3218 ( .A(n3258), .ZN(n383) );
  XOR2_X2 U3219 ( .A(b[6]), .B(n305), .Z(n3259) );
  INV_X4 U3220 ( .A(n3259), .ZN(n356) );
  XNOR2_X2 U3221 ( .A(n3261), .B(n323), .ZN(n3260) );
  AND2_X2 U3222 ( .A1(n2968), .A2(n3233), .ZN(n3262) );
  INV_X8 U3223 ( .A(n3262), .ZN(n419) );
  XNOR2_X2 U3224 ( .A(n314), .B(n3264), .ZN(n3263) );
  OAI22_X1 U3225 ( .A1(n419), .A2(n2657), .B1(n3235), .B2(n2656), .ZN(n2131)
         );
  XOR2_X2 U3226 ( .A(b[4]), .B(n302), .Z(n3265) );
  OAI22_X1 U3227 ( .A1(n401), .A2(n2843), .B1(n2842), .B2(n3227), .ZN(n2316)
         );
  AOI21_X2 U3228 ( .B1(n749), .B2(n916), .A(n742), .ZN(n738) );
  NAND2_X1 U3229 ( .A1(n748), .A2(n916), .ZN(n737) );
  NAND2_X1 U3230 ( .A1(n916), .A2(n744), .ZN(n477) );
  XNOR2_X2 U3231 ( .A(n3267), .B(n329), .ZN(n3266) );
  INV_X8 U3232 ( .A(n3266), .ZN(n380) );
  XNOR2_X2 U3233 ( .A(n3269), .B(n311), .ZN(n3268) );
  OAI22_X1 U3234 ( .A1(n398), .A2(n2876), .B1(n350), .B2(n2875), .ZN(n2349) );
  AOI21_X2 U3235 ( .B1(n917), .B2(n760), .A(n753), .ZN(n747) );
  NAND2_X1 U3236 ( .A1(n917), .A2(n918), .ZN(n746) );
  NAND2_X1 U3237 ( .A1(n917), .A2(n755), .ZN(n478) );
  NAND2_X2 U3238 ( .A1(n669), .A2(n652), .ZN(n650) );
  XNOR2_X1 U3239 ( .A(n646), .B(n462), .ZN(product[42]) );
  XOR2_X1 U3240 ( .A(n632), .B(n460), .Z(product[44]) );
  AOI21_X1 U3241 ( .B1(n646), .B2(n514), .A(n515), .ZN(n513) );
  AOI21_X1 U3242 ( .B1(n646), .B2(n519), .A(n520), .ZN(n518) );
  AOI21_X1 U3243 ( .B1(n646), .B2(n901), .A(n643), .ZN(n641) );
  AOI21_X1 U3244 ( .B1(n646), .B2(n585), .A(n586), .ZN(n584) );
  OAI21_X2 U3245 ( .B1(n632), .B2(n626), .A(n627), .ZN(n625) );
  NAND2_X2 U3246 ( .A1(n1510), .A2(n1535), .ZN(n735) );
  AOI21_X2 U3247 ( .B1(n646), .B2(n633), .A(n634), .ZN(n632) );
  NOR2_X2 U3248 ( .A1(n1394), .A2(n1423), .ZN(n705) );
  NAND2_X2 U3249 ( .A1(n1394), .A2(n1423), .ZN(n706) );
  OAI21_X2 U3250 ( .B1(n705), .B2(n715), .A(n706), .ZN(n704) );
  XNOR2_X1 U3251 ( .A(n609), .B(n457), .ZN(product[47]) );
  AND2_X2 U3252 ( .A1(n2963), .A2(n386), .ZN(n3273) );
  INV_X8 U3253 ( .A(n3273), .ZN(n434) );
  OAI22_X1 U3254 ( .A1(n434), .A2(n3011), .B1(n386), .B2(n2499), .ZN(n1875) );
  INV_X1 U3255 ( .A(n785), .ZN(n784) );
  AOI21_X2 U3256 ( .B1(n786), .B2(n805), .A(n787), .ZN(n785) );
  OAI21_X1 U3257 ( .B1(n647), .B2(n567), .A(n568), .ZN(n566) );
  OAI21_X1 U3258 ( .B1(n647), .B2(n610), .A(n611), .ZN(n609) );
  OAI21_X1 U3259 ( .B1(n647), .B2(n507), .A(n508), .ZN(n506) );
  INV_X1 U3260 ( .A(n3204), .ZN(n3294) );
  XNOR2_X1 U3261 ( .A(n3191), .B(n2122), .ZN(n1422) );
  OAI22_X1 U3262 ( .A1(n3205), .A2(n2462), .B1(n389), .B2(n2461), .ZN(n1943)
         );
  NOR2_X1 U3263 ( .A1(n1536), .A2(n1561), .ZN(n743) );
  OAI22_X1 U3264 ( .A1(n416), .A2(n2687), .B1(n3198), .B2(n2686), .ZN(n2161)
         );
  OAI22_X1 U3265 ( .A1(n422), .A2(n2627), .B1(n374), .B2(n2626), .ZN(n2101) );
  NOR2_X1 U3266 ( .A1(n1712), .A2(n1729), .ZN(n795) );
  NAND2_X1 U3267 ( .A1(n1712), .A2(n1729), .ZN(n796) );
  AOI21_X2 U3268 ( .B1(n924), .B2(n801), .A(n794), .ZN(n792) );
  OAI21_X1 U3269 ( .B1(n792), .B2(n788), .A(n789), .ZN(n787) );
  OAI21_X1 U3270 ( .B1(n804), .B2(n791), .A(n792), .ZN(n790) );
  OAI22_X1 U3271 ( .A1(n410), .A2(n2750), .B1(n362), .B2(n2749), .ZN(n2223) );
  AOI21_X2 U3272 ( .B1(n3194), .B2(n728), .A(n729), .ZN(n727) );
  NOR2_X2 U3273 ( .A1(n730), .A2(n746), .ZN(n728) );
  OAI22_X1 U3274 ( .A1(n428), .A2(n2564), .B1(n380), .B2(n2563), .ZN(n2041) );
  OAI22_X1 U3275 ( .A1(n425), .A2(n3014), .B1(n3209), .B2(n2598), .ZN(n1878)
         );
  XOR2_X1 U3276 ( .A(n716), .B(n473), .Z(product[31]) );
  AOI21_X1 U3277 ( .B1(n726), .B2(n717), .A(n718), .ZN(n716) );
  OAI21_X1 U3278 ( .B1(n763), .B2(n746), .A(n747), .ZN(n745) );
  INV_X1 U3279 ( .A(n747), .ZN(n749) );
  INV_X2 U3280 ( .A(n504), .ZN(product[63]) );
  INV_X2 U3281 ( .A(n503), .ZN(product[1]) );
  INV_X2 U3282 ( .A(n991), .ZN(n992) );
  INV_X2 U3283 ( .A(n973), .ZN(n974) );
  INV_X2 U3284 ( .A(n959), .ZN(n960) );
  INV_X2 U3285 ( .A(n949), .ZN(n950) );
  INV_X2 U3286 ( .A(n943), .ZN(n944) );
  INV_X2 U3287 ( .A(n881), .ZN(n942) );
  INV_X2 U3288 ( .A(n879), .ZN(n941) );
  INV_X2 U3289 ( .A(n871), .ZN(n939) );
  INV_X2 U3290 ( .A(n863), .ZN(n937) );
  INV_X2 U3291 ( .A(n855), .ZN(n935) );
  INV_X2 U3292 ( .A(n851), .ZN(n934) );
  INV_X2 U3293 ( .A(n848), .ZN(n933) );
  INV_X2 U3294 ( .A(n829), .ZN(n930) );
  INV_X2 U3295 ( .A(n826), .ZN(n929) );
  INV_X2 U3296 ( .A(n815), .ZN(n927) );
  INV_X2 U3297 ( .A(n788), .ZN(n923) );
  INV_X2 U3298 ( .A(n777), .ZN(n921) );
  INV_X2 U3299 ( .A(n772), .ZN(n920) );
  INV_X2 U3300 ( .A(n705), .ZN(n911) );
  INV_X2 U3301 ( .A(n697), .ZN(n910) );
  INV_X2 U3302 ( .A(n674), .ZN(n906) );
  INV_X2 U3303 ( .A(n618), .ZN(n897) );
  INV_X2 U3304 ( .A(n563), .ZN(n891) );
  INV_X2 U3305 ( .A(n560), .ZN(n890) );
  INV_X2 U3306 ( .A(n555), .ZN(n889) );
  INV_X2 U3307 ( .A(n552), .ZN(n888) );
  INV_X2 U3308 ( .A(n539), .ZN(n887) );
  INV_X2 U3309 ( .A(n536), .ZN(n886) );
  INV_X2 U3310 ( .A(n516), .ZN(n884) );
  INV_X2 U3311 ( .A(n877), .ZN(n875) );
  INV_X2 U3312 ( .A(n876), .ZN(n940) );
  INV_X2 U3313 ( .A(n869), .ZN(n867) );
  INV_X2 U3314 ( .A(n868), .ZN(n938) );
  INV_X2 U3315 ( .A(n861), .ZN(n859) );
  INV_X2 U3316 ( .A(n860), .ZN(n936) );
  INV_X2 U3317 ( .A(n854), .ZN(n853) );
  INV_X2 U3318 ( .A(n845), .ZN(n844) );
  INV_X2 U3319 ( .A(n843), .ZN(n841) );
  INV_X2 U3320 ( .A(n842), .ZN(n932) );
  INV_X2 U3321 ( .A(n838), .ZN(n836) );
  INV_X2 U3322 ( .A(n837), .ZN(n931) );
  INV_X2 U3323 ( .A(n832), .ZN(n831) );
  INV_X2 U3324 ( .A(n823), .ZN(n822) );
  INV_X2 U3325 ( .A(n821), .ZN(n819) );
  INV_X2 U3326 ( .A(n820), .ZN(n928) );
  INV_X2 U3327 ( .A(n811), .ZN(n809) );
  INV_X2 U3328 ( .A(n810), .ZN(n926) );
  INV_X2 U3329 ( .A(n805), .ZN(n804) );
  INV_X2 U3330 ( .A(n799), .ZN(n801) );
  INV_X2 U3331 ( .A(n798), .ZN(n925) );
  INV_X2 U3332 ( .A(n795), .ZN(n924) );
  INV_X2 U3333 ( .A(n783), .ZN(n781) );
  INV_X2 U3334 ( .A(n782), .ZN(n922) );
  INV_X2 U3335 ( .A(n764), .ZN(n763) );
  INV_X2 U3336 ( .A(n757), .ZN(n918) );
  INV_X2 U3337 ( .A(n755), .ZN(n753) );
  INV_X2 U3338 ( .A(n754), .ZN(n917) );
  INV_X2 U3339 ( .A(n746), .ZN(n748) );
  INV_X2 U3340 ( .A(n735), .ZN(n733) );
  INV_X2 U3341 ( .A(n734), .ZN(n915) );
  INV_X2 U3342 ( .A(n725), .ZN(n723) );
  INV_X2 U3343 ( .A(n724), .ZN(n914) );
  INV_X2 U3344 ( .A(n715), .ZN(n713) );
  INV_X2 U3345 ( .A(n714), .ZN(n912) );
  INV_X2 U3346 ( .A(n711), .ZN(n709) );
  INV_X2 U3347 ( .A(n710), .ZN(n708) );
  INV_X2 U3348 ( .A(n692), .ZN(n690) );
  INV_X2 U3349 ( .A(n688), .ZN(n686) );
  INV_X2 U3350 ( .A(n687), .ZN(n908) );
  INV_X2 U3351 ( .A(n677), .ZN(n676) );
  INV_X2 U3352 ( .A(n664), .ZN(n662) );
  INV_X2 U3353 ( .A(n658), .ZN(n902) );
  INV_X2 U3354 ( .A(n647), .ZN(n646) );
  INV_X2 U3355 ( .A(n645), .ZN(n643) );
  INV_X2 U3356 ( .A(n644), .ZN(n901) );
  INV_X2 U3357 ( .A(n640), .ZN(n638) );
  INV_X2 U3358 ( .A(n639), .ZN(n900) );
  INV_X2 U3359 ( .A(n636), .ZN(n634) );
  INV_X2 U3360 ( .A(n635), .ZN(n633) );
  INV_X2 U3361 ( .A(n627), .ZN(n629) );
  INV_X2 U3362 ( .A(n626), .ZN(n899) );
  INV_X2 U3363 ( .A(n624), .ZN(n622) );
  INV_X2 U3364 ( .A(n623), .ZN(n898) );
  INV_X2 U3365 ( .A(n613), .ZN(n611) );
  INV_X2 U3366 ( .A(n612), .ZN(n610) );
  INV_X2 U3367 ( .A(n608), .ZN(n606) );
  INV_X2 U3368 ( .A(n607), .ZN(n896) );
  INV_X2 U3369 ( .A(n599), .ZN(n601) );
  INV_X2 U3370 ( .A(n596), .ZN(n594) );
  INV_X2 U3371 ( .A(n595), .ZN(n894) );
  INV_X2 U3372 ( .A(n590), .ZN(n588) );
  INV_X2 U3373 ( .A(n589), .ZN(n587) );
  INV_X2 U3374 ( .A(n579), .ZN(n581) );
  INV_X2 U3375 ( .A(n578), .ZN(n893) );
  INV_X2 U3376 ( .A(n576), .ZN(n574) );
  INV_X2 U3377 ( .A(n575), .ZN(n892) );
  INV_X2 U3378 ( .A(n572), .ZN(n570) );
  INV_X2 U3379 ( .A(n571), .ZN(n569) );
  INV_X2 U3380 ( .A(n566), .ZN(n565) );
  INV_X2 U3381 ( .A(n545), .ZN(n543) );
  INV_X2 U3382 ( .A(n544), .ZN(n542) );
  INV_X2 U3383 ( .A(n535), .ZN(n533) );
  INV_X2 U3384 ( .A(n534), .ZN(n532) );
  INV_X2 U3385 ( .A(n530), .ZN(n528) );
  INV_X2 U3386 ( .A(n529), .ZN(n885) );
  INV_X2 U3387 ( .A(n522), .ZN(n520) );
  INV_X2 U3388 ( .A(n521), .ZN(n519) );
  INV_X2 U3389 ( .A(n512), .ZN(n510) );
  INV_X2 U3390 ( .A(n511), .ZN(n883) );
  INV_X2 U3391 ( .A(n299), .ZN(n3024) );
  INV_X2 U3392 ( .A(n302), .ZN(n3023) );
  INV_X2 U3393 ( .A(n305), .ZN(n3022) );
  INV_X2 U3394 ( .A(n308), .ZN(n3021) );
  INV_X2 U3395 ( .A(n311), .ZN(n3020) );
  INV_X2 U3396 ( .A(n314), .ZN(n3019) );
  INV_X2 U3397 ( .A(n317), .ZN(n3018) );
  INV_X2 U3398 ( .A(n320), .ZN(n3017) );
  INV_X2 U3399 ( .A(n323), .ZN(n3016) );
  INV_X2 U3400 ( .A(n326), .ZN(n3015) );
  INV_X2 U3401 ( .A(n329), .ZN(n3014) );
  INV_X2 U3402 ( .A(n332), .ZN(n3013) );
  INV_X2 U3403 ( .A(n335), .ZN(n3012) );
  INV_X2 U3404 ( .A(n338), .ZN(n3011) );
  INV_X2 U3405 ( .A(n342), .ZN(n3009) );
  NAND2_X2 U3406 ( .A1(n3218), .A2(n3275), .ZN(n2928) );
  NAND2_X2 U3407 ( .A1(n302), .A2(n3275), .ZN(n2895) );
  NAND2_X2 U3408 ( .A1(n305), .A2(n3275), .ZN(n2862) );
  NAND2_X2 U3409 ( .A1(n308), .A2(n3275), .ZN(n2829) );
  NAND2_X2 U3410 ( .A1(n311), .A2(n3275), .ZN(n2796) );
  NAND2_X2 U3411 ( .A1(n314), .A2(n3275), .ZN(n2763) );
  NAND2_X2 U3412 ( .A1(n317), .A2(n3275), .ZN(n2730) );
  NAND2_X2 U3413 ( .A1(n320), .A2(n3275), .ZN(n2697) );
  NAND2_X2 U3414 ( .A1(n323), .A2(n3275), .ZN(n2664) );
  NAND2_X2 U3415 ( .A1(n326), .A2(n3275), .ZN(n2631) );
  NAND2_X2 U3416 ( .A1(n329), .A2(n3275), .ZN(n2598) );
  NAND2_X2 U3417 ( .A1(n332), .A2(n3275), .ZN(n2565) );
  NAND2_X2 U3418 ( .A1(n335), .A2(n3275), .ZN(n2532) );
  NAND2_X2 U3419 ( .A1(n338), .A2(n3275), .ZN(n2499) );
  NAND2_X2 U3420 ( .A1(n341), .A2(n3275), .ZN(n2466) );
  NAND2_X2 U3421 ( .A1(n342), .A2(n3275), .ZN(n2433) );
  OAI21_X2 U3422 ( .B1(b[0]), .B2(n3276), .A(n3277), .ZN(n2369) );
  INV_X2 U3423 ( .A(n2896), .ZN(n3277) );
  INV_X2 U3424 ( .A(n395), .ZN(n3276) );
  NOR2_X2 U3425 ( .A1(n350), .A2(n3275), .ZN(n2368) );
  INV_X2 U3426 ( .A(n2863), .ZN(n3278) );
  NOR2_X2 U3427 ( .A1(n3226), .A2(n3275), .ZN(n2335) );
  INV_X2 U3428 ( .A(n2830), .ZN(n3279) );
  NOR2_X2 U3429 ( .A1(n3231), .A2(n3275), .ZN(n2302) );
  OAI21_X2 U3430 ( .B1(n3280), .B2(n3259), .A(n3281), .ZN(n2270) );
  INV_X2 U3431 ( .A(n2797), .ZN(n3281) );
  NOR2_X2 U3432 ( .A1(n359), .A2(n3275), .ZN(n2269) );
  INV_X2 U3433 ( .A(n2764), .ZN(n3282) );
  NOR2_X2 U3434 ( .A1(n362), .A2(n3275), .ZN(n2236) );
  INV_X2 U3435 ( .A(n2731), .ZN(n3283) );
  NOR2_X2 U3436 ( .A1(n365), .A2(n3275), .ZN(n2203) );
  INV_X2 U3437 ( .A(n2698), .ZN(n3285) );
  NOR2_X2 U3438 ( .A1(n3197), .A2(n3275), .ZN(n2171) );
  INV_X2 U3439 ( .A(n2665), .ZN(n3286) );
  NOR2_X2 U3440 ( .A1(n3234), .A2(n3275), .ZN(n2138) );
  OAI21_X2 U3441 ( .B1(n3262), .B2(n3253), .A(n3287), .ZN(n2106) );
  INV_X2 U3442 ( .A(n2632), .ZN(n3287) );
  NOR2_X2 U3443 ( .A1(n3193), .A2(n3275), .ZN(n2105) );
  INV_X2 U3444 ( .A(n2599), .ZN(n3288) );
  NOR2_X2 U3445 ( .A1(n3208), .A2(n3275), .ZN(n2072) );
  INV_X2 U3446 ( .A(n2566), .ZN(n3289) );
  NOR2_X2 U3447 ( .A1(n380), .A2(n3275), .ZN(n2042) );
  OAI21_X2 U3448 ( .B1(n3171), .B2(n3266), .A(n3290), .ZN(n2010) );
  INV_X2 U3449 ( .A(n2533), .ZN(n3290) );
  NOR2_X2 U3450 ( .A1(n3212), .A2(n3275), .ZN(n2009) );
  OAI21_X2 U3451 ( .B1(n3291), .B2(n3258), .A(n3292), .ZN(n1979) );
  INV_X2 U3452 ( .A(n2500), .ZN(n3292) );
  INV_X2 U3453 ( .A(n431), .ZN(n3291) );
  NOR2_X2 U3454 ( .A1(n386), .A2(n3275), .ZN(n1978) );
  INV_X2 U3455 ( .A(n2467), .ZN(n3293) );
  NOR2_X2 U3456 ( .A1(n389), .A2(n3275), .ZN(n1947) );
  INV_X2 U3457 ( .A(n2434), .ZN(n3295) );
  OAI21_X2 U3458 ( .B1(n3296), .B2(n3246), .A(n3297), .ZN(n1889) );
  INV_X2 U3459 ( .A(n2401), .ZN(n3297) );
  INV_X2 U3460 ( .A(n1279), .ZN(n1280) );
  INV_X2 U3461 ( .A(n1229), .ZN(n1230) );
  INV_X2 U3462 ( .A(n1141), .ZN(n1142) );
  INV_X2 U3463 ( .A(n1103), .ZN(n1104) );
  INV_X2 U3464 ( .A(n1069), .ZN(n1070) );
  INV_X2 U3465 ( .A(n1039), .ZN(n1040) );
  INV_X2 U3466 ( .A(n1013), .ZN(n1014) );
endmodule


module up_island_DW01_sub_1 ( A, B, DIFF, CI, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n123, n124, n126,
         n127, n128, n129, n130, n131, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n148, n149, n150, n151, n152, n153, n154, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n176, n177, n178, n179, n180,
         n181, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n200, n201, n202, n203, n204, n205, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n228, n229, n230, n231, n232,
         n233, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n252, n253, n254, n255, n256, n257, n261,
         n262, n263, n264, n265, n266, n267, n268, n271, n272, n273, n274,
         n277, n278, n279, n280, n281, n282, n284, n285, n286, n287, n288,
         n289, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n308, n309, n310, n311, n312, n313, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n331, n333, n337, n338, n339, n340, n341, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n363, n364, n365, n366, n368, n370, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n388,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  NAND2_X4 U6 ( .A1(n386), .A2(n37), .ZN(n5) );
  NAND2_X4 U20 ( .A1(n45), .A2(n48), .ZN(n6) );
  NAND2_X4 U32 ( .A1(n388), .A2(n57), .ZN(n7) );
  NAND2_X4 U38 ( .A1(n413), .A2(n61), .ZN(n59) );
  AOI21_X4 U39 ( .B1(n370), .B2(n61), .A(n62), .ZN(n60) );
  NOR2_X4 U46 ( .A1(n69), .A2(n93), .ZN(n67) );
  OAI21_X4 U47 ( .B1(n94), .B2(n69), .A(n70), .ZN(n68) );
  NAND2_X4 U48 ( .A1(n80), .A2(n71), .ZN(n69) );
  AOI21_X4 U49 ( .B1(n71), .B2(n81), .A(n72), .ZN(n70) );
  NAND2_X4 U52 ( .A1(n71), .A2(n74), .ZN(n8) );
  XNOR2_X2 U56 ( .A(n84), .B(n9), .ZN(DIFF[27]) );
  NAND2_X4 U58 ( .A1(n87), .A2(n80), .ZN(n76) );
  NAND2_X4 U64 ( .A1(n80), .A2(n83), .ZN(n9) );
  XNOR2_X2 U68 ( .A(n99), .B(n10), .ZN(DIFF[26]) );
  NOR2_X4 U72 ( .A1(n4), .A2(n89), .ZN(n87) );
  NAND2_X4 U78 ( .A1(n392), .A2(n95), .ZN(n93) );
  AOI21_X4 U79 ( .B1(n95), .B2(n105), .A(n96), .ZN(n94) );
  NAND2_X4 U82 ( .A1(n95), .A2(n98), .ZN(n10) );
  NAND2_X4 U88 ( .A1(n111), .A2(n392), .ZN(n100) );
  AOI21_X4 U89 ( .B1(n112), .B2(n392), .A(n105), .ZN(n101) );
  NAND2_X4 U94 ( .A1(n392), .A2(n107), .ZN(n11) );
  XNOR2_X2 U98 ( .A(n129), .B(n12), .ZN(DIFF[24]) );
  NAND2_X4 U114 ( .A1(n394), .A2(n393), .ZN(n123) );
  AOI21_X4 U115 ( .B1(n135), .B2(n393), .A(n126), .ZN(n124) );
  NAND2_X4 U118 ( .A1(n393), .A2(n128), .ZN(n12) );
  XNOR2_X2 U122 ( .A(n138), .B(n13), .ZN(DIFF[23]) );
  NAND2_X4 U124 ( .A1(n141), .A2(n394), .ZN(n130) );
  AOI21_X4 U125 ( .B1(n142), .B2(n394), .A(n135), .ZN(n131) );
  NAND2_X4 U130 ( .A1(n394), .A2(n137), .ZN(n13) );
  XNOR2_X2 U134 ( .A(n151), .B(n14), .ZN(DIFF[22]) );
  NAND2_X4 U146 ( .A1(n395), .A2(n150), .ZN(n14) );
  XNOR2_X2 U150 ( .A(n160), .B(n15), .ZN(DIFF[21]) );
  NOR2_X4 U156 ( .A1(n165), .A2(n158), .ZN(n154) );
  NAND2_X4 U158 ( .A1(n396), .A2(n159), .ZN(n15) );
  XNOR2_X2 U162 ( .A(n179), .B(n16), .ZN(DIFF[20]) );
  NAND2_X4 U164 ( .A1(n413), .A2(n163), .ZN(n161) );
  AOI21_X4 U165 ( .B1(n370), .B2(n163), .A(n164), .ZN(n162) );
  AOI21_X4 U177 ( .B1(n397), .B2(n185), .A(n176), .ZN(n174) );
  XNOR2_X2 U184 ( .A(n188), .B(n17), .ZN(DIFF[19]) );
  NAND2_X4 U186 ( .A1(n191), .A2(n398), .ZN(n180) );
  AOI21_X4 U187 ( .B1(n192), .B2(n398), .A(n185), .ZN(n181) );
  NAND2_X4 U192 ( .A1(n398), .A2(n187), .ZN(n17) );
  XNOR2_X2 U196 ( .A(n203), .B(n18), .ZN(DIFF[18]) );
  NOR2_X4 U200 ( .A1(n4), .A2(n193), .ZN(n191) );
  OAI21_X4 U201 ( .B1(n368), .B2(n193), .A(n194), .ZN(n192) );
  NAND2_X4 U202 ( .A1(n219), .A2(n195), .ZN(n193) );
  AOI21_X4 U203 ( .B1(n220), .B2(n195), .A(n196), .ZN(n194) );
  AOI21_X4 U207 ( .B1(n399), .B2(n209), .A(n200), .ZN(n198) );
  XNOR2_X2 U214 ( .A(n212), .B(n19), .ZN(DIFF[17]) );
  NAND2_X4 U216 ( .A1(n215), .A2(n400), .ZN(n204) );
  AOI21_X4 U217 ( .B1(n216), .B2(n400), .A(n209), .ZN(n205) );
  XNOR2_X2 U226 ( .A(n231), .B(n20), .ZN(DIFF[16]) );
  NOR2_X4 U230 ( .A1(n4), .A2(n217), .ZN(n215) );
  OAI21_X4 U231 ( .B1(n368), .B2(n217), .A(n218), .ZN(n216) );
  NOR2_X4 U234 ( .A1(n273), .A2(n221), .ZN(n219) );
  NOR2_X4 U238 ( .A1(n249), .A2(n225), .ZN(n223) );
  AOI21_X4 U241 ( .B1(n401), .B2(n237), .A(n228), .ZN(n226) );
  XNOR2_X2 U248 ( .A(n240), .B(n21), .ZN(DIFF[15]) );
  XNOR2_X2 U260 ( .A(n255), .B(n22), .ZN(DIFF[14]) );
  NOR2_X4 U264 ( .A1(n4), .A2(n245), .ZN(n243) );
  AOI21_X4 U271 ( .B1(n403), .B2(n261), .A(n252), .ZN(n250) );
  XNOR2_X2 U278 ( .A(n264), .B(n23), .ZN(DIFF[13]) );
  XNOR2_X2 U290 ( .A(n287), .B(n24), .ZN(DIFF[12]) );
  NOR2_X4 U294 ( .A1(n4), .A2(n273), .ZN(n267) );
  AOI21_X4 U309 ( .B1(n405), .B2(n293), .A(n284), .ZN(n282) );
  XNOR2_X2 U316 ( .A(n296), .B(n25), .ZN(DIFF[11]) );
  XNOR2_X2 U328 ( .A(n311), .B(n26), .ZN(DIFF[10]) );
  NOR2_X4 U332 ( .A1(n4), .A2(n301), .ZN(n299) );
  OAI21_X4 U333 ( .B1(n368), .B2(n301), .A(n302), .ZN(n300) );
  NAND2_X4 U334 ( .A1(n327), .A2(n303), .ZN(n301) );
  AOI21_X4 U339 ( .B1(n407), .B2(n317), .A(n308), .ZN(n306) );
  XNOR2_X2 U346 ( .A(n320), .B(n27), .ZN(DIFF[9]) );
  XNOR2_X2 U358 ( .A(n339), .B(n28), .ZN(DIFF[8]) );
  XNOR2_X2 U380 ( .A(n348), .B(n29), .ZN(DIFF[7]) );
  XNOR2_X2 U392 ( .A(n359), .B(n30), .ZN(DIFF[6]) );
  NOR2_X4 U396 ( .A1(n4), .A2(n353), .ZN(n351) );
  OAI21_X4 U397 ( .B1(n368), .B2(n353), .A(n354), .ZN(n352) );
  NAND2_X4 U402 ( .A1(n411), .A2(n358), .ZN(n30) );
  XNOR2_X2 U406 ( .A(n366), .B(n31), .ZN(DIFF[5]) );
  NAND2_X4 U408 ( .A1(n413), .A2(n412), .ZN(n360) );
  AOI21_X4 U409 ( .B1(n370), .B2(n412), .A(n363), .ZN(n361) );
  NAND2_X4 U412 ( .A1(n412), .A2(n567), .ZN(n31) );
  NAND2_X4 U422 ( .A1(n413), .A2(n368), .ZN(n32) );
  NOR2_X4 U424 ( .A1(n584), .A2(A[4]), .ZN(n4) );
  NAND2_X4 U425 ( .A1(n584), .A2(A[4]), .ZN(n368) );
  XNOR2_X2 U426 ( .A(n378), .B(n33), .ZN(DIFF[3]) );
  AOI21_X4 U427 ( .B1(n374), .B2(n382), .A(n375), .ZN(n2) );
  OAI21_X4 U429 ( .B1(n380), .B2(n376), .A(n377), .ZN(n375) );
  NAND2_X4 U430 ( .A1(n414), .A2(n377), .ZN(n33) );
  NOR2_X4 U432 ( .A1(n585), .A2(A[3]), .ZN(n376) );
  XOR2_X2 U434 ( .A(n34), .B(n381), .Z(DIFF[2]) );
  OAI21_X4 U435 ( .B1(n381), .B2(n379), .A(n380), .ZN(n378) );
  NAND2_X4 U436 ( .A1(n415), .A2(n380), .ZN(n34) );
  XOR2_X2 U440 ( .A(n35), .B(n385), .Z(DIFF[1]) );
  NAND2_X4 U443 ( .A1(n416), .A2(n384), .ZN(n35) );
  NOR2_X4 U445 ( .A1(n587), .A2(A[1]), .ZN(n383) );
  INV_X1 U484 ( .A(B[31]), .ZN(n417) );
  NAND2_X1 U485 ( .A1(A[29]), .A2(n419), .ZN(n57) );
  NOR2_X1 U486 ( .A1(A[29]), .A2(n419), .ZN(n56) );
  AOI21_X2 U487 ( .B1(n554), .B2(n395), .A(n148), .ZN(n577) );
  NAND2_X2 U488 ( .A1(n551), .A2(n552), .ZN(n553) );
  NAND2_X1 U489 ( .A1(n553), .A2(n40), .ZN(n38) );
  INV_X4 U490 ( .A(n2), .ZN(n551) );
  INV_X1 U491 ( .A(n39), .ZN(n552) );
  OAI21_X1 U492 ( .B1(n166), .B2(n158), .A(n159), .ZN(n554) );
  AOI21_X1 U493 ( .B1(n116), .B2(n67), .A(n68), .ZN(n64) );
  INV_X2 U494 ( .A(n186), .ZN(n398) );
  CLKBUF_X1 U495 ( .A(n399), .Z(n555) );
  OAI21_X2 U496 ( .B1(n559), .B2(n347), .A(n338), .ZN(n569) );
  AOI21_X2 U497 ( .B1(n272), .B2(n167), .A(n168), .ZN(n166) );
  AOI21_X1 U498 ( .B1(n157), .B2(n395), .A(n148), .ZN(n578) );
  XNOR2_X1 U499 ( .A(n588), .B(A[0]), .ZN(DIFF[0]) );
  NOR2_X1 U500 ( .A1(n588), .A2(A[0]), .ZN(n385) );
  NAND2_X1 U501 ( .A1(n556), .A2(n557), .ZN(n558) );
  NAND2_X1 U502 ( .A1(n558), .A2(n90), .ZN(n88) );
  INV_X1 U503 ( .A(n368), .ZN(n556) );
  INV_X1 U504 ( .A(n89), .ZN(n557) );
  AOI21_X1 U505 ( .B1(n579), .B2(n91), .A(n92), .ZN(n90) );
  NOR2_X1 U506 ( .A1(n586), .A2(A[2]), .ZN(n379) );
  NAND2_X1 U507 ( .A1(n586), .A2(A[2]), .ZN(n380) );
  NOR2_X1 U508 ( .A1(A[8]), .A2(n440), .ZN(n559) );
  NOR2_X1 U509 ( .A1(n440), .A2(A[8]), .ZN(n337) );
  NAND2_X1 U510 ( .A1(n397), .A2(n178), .ZN(n16) );
  INV_X1 U511 ( .A(n178), .ZN(n176) );
  INV_X1 U512 ( .A(n355), .ZN(n353) );
  AOI21_X1 U513 ( .B1(n356), .B2(n331), .A(n569), .ZN(n560) );
  AOI21_X1 U514 ( .B1(n356), .B2(n331), .A(n569), .ZN(n326) );
  NAND2_X1 U515 ( .A1(n400), .A2(n211), .ZN(n19) );
  OAI21_X1 U516 ( .B1(n560), .B2(n277), .A(n278), .ZN(n561) );
  OAI21_X1 U517 ( .B1(n326), .B2(n277), .A(n278), .ZN(n272) );
  NOR2_X2 U518 ( .A1(n4), .A2(n113), .ZN(n111) );
  OAI21_X2 U519 ( .B1(n368), .B2(n113), .A(n114), .ZN(n112) );
  XNOR2_X1 U520 ( .A(n108), .B(n11), .ZN(DIFF[25]) );
  AOI21_X1 U521 ( .B1(n561), .B2(n247), .A(n248), .ZN(n246) );
  OAI21_X1 U522 ( .B1(n368), .B2(n245), .A(n246), .ZN(n244) );
  OAI21_X1 U523 ( .B1(n274), .B2(n221), .A(n222), .ZN(n220) );
  OAI21_X1 U524 ( .B1(n368), .B2(n273), .A(n274), .ZN(n268) );
  AOI21_X2 U525 ( .B1(n328), .B2(n303), .A(n304), .ZN(n302) );
  NAND2_X1 U526 ( .A1(n408), .A2(n407), .ZN(n305) );
  CLKBUF_X1 U527 ( .A(n560), .Z(n562) );
  INV_X1 U528 ( .A(n357), .ZN(n563) );
  INV_X1 U529 ( .A(n563), .ZN(n564) );
  NAND2_X1 U530 ( .A1(n405), .A2(n286), .ZN(n24) );
  INV_X1 U531 ( .A(n286), .ZN(n284) );
  INV_X1 U532 ( .A(B[18]), .ZN(n565) );
  INV_X1 U533 ( .A(n200), .ZN(n566) );
  NAND2_X1 U534 ( .A1(n407), .A2(n310), .ZN(n26) );
  INV_X1 U535 ( .A(n310), .ZN(n308) );
  AOI21_X1 U536 ( .B1(n244), .B2(n402), .A(n237), .ZN(n233) );
  NAND2_X1 U537 ( .A1(n243), .A2(n402), .ZN(n232) );
  NAND2_X2 U538 ( .A1(n402), .A2(n401), .ZN(n225) );
  INV_X1 U539 ( .A(n363), .ZN(n567) );
  INV_X1 U540 ( .A(n365), .ZN(n363) );
  AOI21_X1 U541 ( .B1(n324), .B2(n408), .A(n317), .ZN(n313) );
  NAND2_X1 U542 ( .A1(n323), .A2(n408), .ZN(n312) );
  XNOR2_X1 U543 ( .A(n58), .B(n7), .ZN(DIFF[29]) );
  XNOR2_X1 U544 ( .A(n75), .B(n8), .ZN(DIFF[28]) );
  INV_X1 U545 ( .A(n88), .ZN(n86) );
  AOI21_X1 U546 ( .B1(n88), .B2(n80), .A(n81), .ZN(n77) );
  INV_X1 U547 ( .A(n346), .ZN(n568) );
  NOR2_X1 U548 ( .A1(n305), .A2(n281), .ZN(n279) );
  INV_X1 U549 ( .A(n202), .ZN(n200) );
  INV_X1 U550 ( .A(n356), .ZN(n354) );
  NAND2_X1 U551 ( .A1(n398), .A2(n397), .ZN(n173) );
  NAND2_X1 U552 ( .A1(n400), .A2(n399), .ZN(n197) );
  NAND2_X1 U553 ( .A1(n403), .A2(n254), .ZN(n22) );
  INV_X1 U554 ( .A(n254), .ZN(n252) );
  AOI21_X2 U555 ( .B1(n224), .B2(n171), .A(n172), .ZN(n170) );
  NAND2_X1 U556 ( .A1(n171), .A2(n223), .ZN(n169) );
  INV_X1 U557 ( .A(n337), .ZN(n409) );
  INV_X1 U558 ( .A(n347), .ZN(n345) );
  NAND2_X1 U559 ( .A1(n351), .A2(n568), .ZN(n340) );
  AOI21_X1 U560 ( .B1(n352), .B2(n568), .A(n345), .ZN(n341) );
  INV_X1 U561 ( .A(n346), .ZN(n410) );
  NAND2_X1 U562 ( .A1(n408), .A2(n319), .ZN(n27) );
  INV_X1 U563 ( .A(n280), .ZN(n278) );
  NAND2_X1 U564 ( .A1(n355), .A2(n331), .ZN(n325) );
  NOR2_X1 U565 ( .A1(n143), .A2(n123), .ZN(n570) );
  AND2_X2 U566 ( .A1(n570), .A2(n571), .ZN(n52) );
  AND2_X1 U567 ( .A1(n572), .A2(n67), .ZN(n571) );
  INV_X1 U568 ( .A(n56), .ZN(n572) );
  OR2_X2 U569 ( .A1(n143), .A2(n573), .ZN(n89) );
  OR2_X1 U570 ( .A1(n123), .A2(n574), .ZN(n573) );
  INV_X1 U571 ( .A(n91), .ZN(n574) );
  NOR2_X1 U572 ( .A1(n277), .A2(n325), .ZN(n575) );
  INV_X1 U573 ( .A(n279), .ZN(n277) );
  NOR2_X1 U574 ( .A1(n325), .A2(n277), .ZN(n271) );
  INV_X1 U575 ( .A(n328), .ZN(n576) );
  NAND2_X1 U576 ( .A1(n568), .A2(n347), .ZN(n29) );
  NAND2_X1 U577 ( .A1(n409), .A2(n338), .ZN(n28) );
  OAI21_X1 U578 ( .B1(n198), .B2(n173), .A(n174), .ZN(n172) );
  NOR2_X2 U579 ( .A1(n197), .A2(n173), .ZN(n171) );
  NOR2_X1 U580 ( .A1(n4), .A2(n325), .ZN(n323) );
  INV_X1 U581 ( .A(n325), .ZN(n327) );
  NOR2_X1 U582 ( .A1(n4), .A2(n143), .ZN(n141) );
  NOR2_X2 U583 ( .A1(n143), .A2(n123), .ZN(n115) );
  INV_X1 U584 ( .A(n333), .ZN(n331) );
  INV_X1 U585 ( .A(n63), .ZN(n61) );
  NAND2_X2 U586 ( .A1(n154), .A2(n395), .ZN(n143) );
  NAND2_X1 U587 ( .A1(n413), .A2(n154), .ZN(n152) );
  NAND2_X1 U588 ( .A1(n555), .A2(n566), .ZN(n18) );
  INV_X1 U589 ( .A(n201), .ZN(n399) );
  NAND2_X1 U590 ( .A1(n267), .A2(n404), .ZN(n256) );
  AOI21_X1 U591 ( .B1(n268), .B2(n404), .A(n261), .ZN(n257) );
  NAND2_X1 U592 ( .A1(n404), .A2(n263), .ZN(n23) );
  NAND2_X2 U593 ( .A1(n404), .A2(n403), .ZN(n249) );
  OAI21_X1 U594 ( .B1(n368), .B2(n325), .A(n576), .ZN(n324) );
  INV_X1 U595 ( .A(n562), .ZN(n328) );
  INV_X1 U596 ( .A(B[6]), .ZN(n442) );
  OAI21_X1 U597 ( .B1(n2), .B2(n312), .A(n313), .ZN(n311) );
  XOR2_X1 U598 ( .A(n2), .B(n32), .Z(DIFF[4]) );
  OAI21_X1 U599 ( .B1(n2), .B2(n321), .A(n322), .ZN(n320) );
  OAI21_X1 U600 ( .B1(n2), .B2(n232), .A(n233), .ZN(n231) );
  OAI21_X1 U601 ( .B1(n2), .B2(n256), .A(n257), .ZN(n255) );
  OAI21_X1 U602 ( .B1(n2), .B2(n241), .A(n242), .ZN(n240) );
  OAI21_X1 U603 ( .B1(n2), .B2(n189), .A(n190), .ZN(n188) );
  OAI21_X1 U604 ( .B1(n2), .B2(n297), .A(n298), .ZN(n296) );
  OAI21_X1 U605 ( .B1(n2), .B2(n4), .A(n368), .ZN(n366) );
  OAI21_X1 U606 ( .B1(n2), .B2(n360), .A(n361), .ZN(n359) );
  OAI21_X1 U607 ( .B1(n2), .B2(n288), .A(n289), .ZN(n287) );
  OAI21_X1 U608 ( .B1(n2), .B2(n180), .A(n181), .ZN(n179) );
  OAI21_X1 U609 ( .B1(n2), .B2(n213), .A(n214), .ZN(n212) );
  OAI21_X1 U610 ( .B1(n2), .B2(n204), .A(n205), .ZN(n203) );
  OAI21_X1 U611 ( .B1(n2), .B2(n340), .A(n341), .ZN(n339) );
  OAI21_X1 U612 ( .B1(n2), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U613 ( .B1(n2), .B2(n349), .A(n350), .ZN(n348) );
  OAI21_X1 U614 ( .B1(n2), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U615 ( .B1(n2), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U616 ( .B1(n2), .B2(n139), .A(n140), .ZN(n138) );
  OAI21_X1 U617 ( .B1(n2), .B2(n76), .A(n77), .ZN(n75) );
  OAI21_X1 U618 ( .B1(n2), .B2(n59), .A(n60), .ZN(n58) );
  OAI21_X1 U619 ( .B1(n2), .B2(n85), .A(n86), .ZN(n84) );
  OAI21_X1 U620 ( .B1(n2), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X1 U621 ( .B1(n2), .B2(n161), .A(n162), .ZN(n160) );
  OAI21_X1 U622 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  NAND2_X1 U623 ( .A1(A[30]), .A2(n418), .ZN(n48) );
  NOR2_X1 U624 ( .A1(A[30]), .A2(n418), .ZN(n47) );
  OAI21_X1 U625 ( .B1(n577), .B2(n123), .A(n124), .ZN(n579) );
  OAI21_X1 U626 ( .B1(n578), .B2(n123), .A(n124), .ZN(n116) );
  INV_X1 U627 ( .A(n224), .ZN(n222) );
  OAI21_X1 U628 ( .B1(n166), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U629 ( .B1(n306), .B2(n281), .A(n282), .ZN(n280) );
  CLKBUF_X1 U630 ( .A(n166), .Z(n580) );
  INV_X1 U631 ( .A(n170), .ZN(n168) );
  NAND2_X2 U632 ( .A1(n587), .A2(A[1]), .ZN(n384) );
  NOR2_X1 U633 ( .A1(n379), .A2(n376), .ZN(n374) );
  OAI21_X2 U634 ( .B1(n383), .B2(n385), .A(n384), .ZN(n382) );
  INV_X1 U635 ( .A(n580), .ZN(n164) );
  INV_X1 U636 ( .A(B[11]), .ZN(n437) );
  INV_X1 U637 ( .A(B[5]), .ZN(n443) );
  CLKBUF_X1 U638 ( .A(n577), .Z(n581) );
  CLKBUF_X1 U639 ( .A(n554), .Z(n582) );
  INV_X1 U640 ( .A(n250), .ZN(n248) );
  OAI21_X2 U641 ( .B1(n250), .B2(n225), .A(n226), .ZN(n224) );
  INV_X1 U642 ( .A(B[9]), .ZN(n439) );
  INV_X1 U643 ( .A(B[10]), .ZN(n438) );
  INV_X1 U644 ( .A(B[16]), .ZN(n432) );
  NAND2_X2 U645 ( .A1(n406), .A2(n405), .ZN(n281) );
  AOI21_X2 U646 ( .B1(n300), .B2(n406), .A(n293), .ZN(n289) );
  NAND2_X2 U647 ( .A1(n299), .A2(n406), .ZN(n288) );
  NAND2_X1 U648 ( .A1(n406), .A2(n295), .ZN(n25) );
  NAND2_X1 U649 ( .A1(n402), .A2(n239), .ZN(n21) );
  INV_X1 U650 ( .A(n239), .ZN(n237) );
  INV_X1 U651 ( .A(B[15]), .ZN(n433) );
  NAND2_X1 U652 ( .A1(n401), .A2(n230), .ZN(n20) );
  INV_X1 U653 ( .A(n561), .ZN(n274) );
  NAND2_X1 U654 ( .A1(n575), .A2(n247), .ZN(n245) );
  INV_X1 U655 ( .A(n575), .ZN(n273) );
  INV_X1 U656 ( .A(n115), .ZN(n113) );
  NAND2_X1 U657 ( .A1(n115), .A2(n67), .ZN(n63) );
  NAND2_X2 U658 ( .A1(n271), .A2(n167), .ZN(n165) );
  NAND2_X1 U659 ( .A1(A[28]), .A2(n420), .ZN(n74) );
  NOR2_X1 U660 ( .A1(A[28]), .A2(n420), .ZN(n73) );
  INV_X1 U661 ( .A(B[19]), .ZN(n429) );
  AOI21_X1 U662 ( .B1(n579), .B2(n67), .A(n68), .ZN(n583) );
  INV_X1 U663 ( .A(B[20]), .ZN(n428) );
  NAND2_X2 U664 ( .A1(n585), .A2(A[3]), .ZN(n377) );
  AOI21_X2 U665 ( .B1(n55), .B2(n45), .A(n46), .ZN(n44) );
  NAND2_X1 U666 ( .A1(A[26]), .A2(n422), .ZN(n98) );
  NOR2_X1 U667 ( .A1(A[26]), .A2(n422), .ZN(n97) );
  INV_X1 U668 ( .A(B[13]), .ZN(n435) );
  NOR2_X1 U669 ( .A1(A[27]), .A2(n421), .ZN(n82) );
  NAND2_X1 U670 ( .A1(A[27]), .A2(n421), .ZN(n83) );
  NAND2_X1 U671 ( .A1(n410), .A2(n409), .ZN(n333) );
  OAI21_X1 U672 ( .B1(n368), .B2(n43), .A(n44), .ZN(n42) );
  INV_X1 U673 ( .A(B[17]), .ZN(n431) );
  INV_X1 U674 ( .A(B[14]), .ZN(n434) );
  OAI21_X1 U675 ( .B1(n368), .B2(n143), .A(n581), .ZN(n142) );
  INV_X1 U676 ( .A(B[18]), .ZN(n430) );
  INV_X1 U677 ( .A(B[7]), .ZN(n441) );
  OAI21_X1 U678 ( .B1(n64), .B2(n56), .A(n57), .ZN(n55) );
  INV_X1 U679 ( .A(n583), .ZN(n62) );
  INV_X1 U680 ( .A(n42), .ZN(n40) );
  INV_X1 U681 ( .A(B[8]), .ZN(n440) );
  AOI21_X1 U682 ( .B1(n370), .B2(n154), .A(n582), .ZN(n153) );
  INV_X1 U683 ( .A(n564), .ZN(n411) );
  INV_X1 U684 ( .A(n579), .ZN(n114) );
  OAI21_X2 U685 ( .B1(n357), .B2(n365), .A(n358), .ZN(n356) );
  NOR2_X1 U686 ( .A1(n364), .A2(n564), .ZN(n355) );
  INV_X1 U687 ( .A(B[12]), .ZN(n436) );
  NAND2_X1 U688 ( .A1(A[23]), .A2(n425), .ZN(n137) );
  NOR2_X1 U689 ( .A1(A[23]), .A2(n425), .ZN(n136) );
  NAND2_X1 U690 ( .A1(A[22]), .A2(n426), .ZN(n150) );
  NOR2_X1 U691 ( .A1(A[22]), .A2(n426), .ZN(n149) );
  NAND2_X1 U692 ( .A1(A[24]), .A2(n424), .ZN(n128) );
  NOR2_X1 U693 ( .A1(A[24]), .A2(n424), .ZN(n127) );
  NOR2_X1 U694 ( .A1(A[25]), .A2(n423), .ZN(n106) );
  NAND2_X1 U695 ( .A1(A[25]), .A2(n423), .ZN(n107) );
  NAND2_X1 U696 ( .A1(A[31]), .A2(n417), .ZN(n37) );
  NOR2_X1 U697 ( .A1(A[31]), .A2(n417), .ZN(n36) );
  XNOR2_X1 U698 ( .A(n49), .B(n6), .ZN(DIFF[30]) );
  OAI21_X1 U699 ( .B1(n2), .B2(n50), .A(n51), .ZN(n49) );
  NAND2_X2 U700 ( .A1(A[19]), .A2(n429), .ZN(n187) );
  NAND2_X1 U701 ( .A1(n52), .A2(n45), .ZN(n43) );
  AOI21_X1 U702 ( .B1(n370), .B2(n52), .A(n55), .ZN(n51) );
  NAND2_X1 U703 ( .A1(n413), .A2(n52), .ZN(n50) );
  NOR2_X1 U704 ( .A1(n4), .A2(n43), .ZN(n41) );
  INV_X1 U705 ( .A(n41), .ZN(n39) );
  INV_X1 U706 ( .A(n158), .ZN(n396) );
  NAND2_X1 U707 ( .A1(A[21]), .A2(n427), .ZN(n159) );
  NOR2_X1 U708 ( .A1(A[21]), .A2(n427), .ZN(n158) );
  XNOR2_X1 U709 ( .A(n38), .B(n5), .ZN(DIFF[31]) );
  NAND2_X1 U710 ( .A1(A[18]), .A2(n565), .ZN(n202) );
  NOR2_X1 U711 ( .A1(n430), .A2(A[18]), .ZN(n201) );
  NOR2_X2 U712 ( .A1(n429), .A2(A[19]), .ZN(n186) );
  NAND2_X1 U713 ( .A1(A[15]), .A2(n433), .ZN(n239) );
  NOR2_X1 U714 ( .A1(A[15]), .A2(n433), .ZN(n238) );
  NOR2_X1 U715 ( .A1(A[17]), .A2(n431), .ZN(n210) );
  NAND2_X1 U716 ( .A1(A[17]), .A2(n431), .ZN(n211) );
  NOR2_X1 U717 ( .A1(A[13]), .A2(n435), .ZN(n262) );
  NAND2_X1 U718 ( .A1(A[13]), .A2(n435), .ZN(n263) );
  NOR2_X1 U719 ( .A1(n441), .A2(A[7]), .ZN(n346) );
  NAND2_X1 U720 ( .A1(A[7]), .A2(n441), .ZN(n347) );
  NAND2_X1 U721 ( .A1(A[11]), .A2(n437), .ZN(n295) );
  NOR2_X1 U722 ( .A1(A[11]), .A2(n437), .ZN(n294) );
  NAND2_X1 U723 ( .A1(A[20]), .A2(n428), .ZN(n178) );
  NOR2_X1 U724 ( .A1(A[20]), .A2(n428), .ZN(n177) );
  NAND2_X1 U725 ( .A1(A[16]), .A2(n432), .ZN(n230) );
  NOR2_X1 U726 ( .A1(A[16]), .A2(n432), .ZN(n229) );
  NOR2_X1 U727 ( .A1(A[9]), .A2(n439), .ZN(n318) );
  NAND2_X1 U728 ( .A1(A[9]), .A2(n439), .ZN(n319) );
  NAND2_X1 U729 ( .A1(A[12]), .A2(n436), .ZN(n286) );
  NOR2_X1 U730 ( .A1(A[12]), .A2(n436), .ZN(n285) );
  NAND2_X1 U731 ( .A1(A[6]), .A2(n442), .ZN(n358) );
  NOR2_X1 U732 ( .A1(A[6]), .A2(n442), .ZN(n357) );
  NAND2_X1 U733 ( .A1(A[14]), .A2(n434), .ZN(n254) );
  NOR2_X1 U734 ( .A1(A[14]), .A2(n434), .ZN(n253) );
  NAND2_X1 U735 ( .A1(A[8]), .A2(n440), .ZN(n338) );
  NAND2_X1 U736 ( .A1(A[10]), .A2(n438), .ZN(n310) );
  NOR2_X1 U737 ( .A1(A[10]), .A2(n438), .ZN(n309) );
  NOR2_X1 U738 ( .A1(A[5]), .A2(n443), .ZN(n364) );
  NAND2_X1 U739 ( .A1(A[5]), .A2(n443), .ZN(n365) );
  INV_X1 U740 ( .A(B[4]), .ZN(n584) );
  INV_X1 U741 ( .A(B[3]), .ZN(n585) );
  INV_X1 U742 ( .A(B[2]), .ZN(n586) );
  INV_X1 U743 ( .A(B[1]), .ZN(n587) );
  INV_X1 U744 ( .A(B[0]), .ZN(n588) );
  INV_X2 U745 ( .A(n98), .ZN(n96) );
  INV_X2 U746 ( .A(n94), .ZN(n92) );
  INV_X2 U747 ( .A(n93), .ZN(n91) );
  INV_X2 U748 ( .A(n87), .ZN(n85) );
  INV_X2 U749 ( .A(n83), .ZN(n81) );
  INV_X2 U750 ( .A(n74), .ZN(n72) );
  INV_X2 U751 ( .A(n48), .ZN(n46) );
  INV_X2 U752 ( .A(B[21]), .ZN(n427) );
  INV_X2 U753 ( .A(B[22]), .ZN(n426) );
  INV_X2 U754 ( .A(B[23]), .ZN(n425) );
  INV_X2 U755 ( .A(B[24]), .ZN(n424) );
  INV_X2 U756 ( .A(B[25]), .ZN(n423) );
  INV_X2 U757 ( .A(B[26]), .ZN(n422) );
  INV_X2 U758 ( .A(B[27]), .ZN(n421) );
  INV_X2 U759 ( .A(B[28]), .ZN(n420) );
  INV_X2 U760 ( .A(B[29]), .ZN(n419) );
  INV_X2 U761 ( .A(B[30]), .ZN(n418) );
  INV_X2 U762 ( .A(n383), .ZN(n416) );
  INV_X2 U763 ( .A(n379), .ZN(n415) );
  INV_X2 U764 ( .A(n376), .ZN(n414) );
  INV_X2 U765 ( .A(n97), .ZN(n95) );
  INV_X2 U766 ( .A(n82), .ZN(n80) );
  INV_X2 U767 ( .A(n73), .ZN(n71) );
  INV_X2 U768 ( .A(n56), .ZN(n388) );
  INV_X2 U769 ( .A(n47), .ZN(n45) );
  INV_X2 U770 ( .A(n36), .ZN(n386) );
  INV_X2 U771 ( .A(n382), .ZN(n381) );
  INV_X2 U772 ( .A(n368), .ZN(n370) );
  INV_X2 U773 ( .A(n4), .ZN(n413) );
  INV_X2 U774 ( .A(n364), .ZN(n412) );
  INV_X2 U775 ( .A(n352), .ZN(n350) );
  INV_X2 U776 ( .A(n351), .ZN(n349) );
  INV_X2 U777 ( .A(n324), .ZN(n322) );
  INV_X2 U778 ( .A(n323), .ZN(n321) );
  INV_X2 U779 ( .A(n319), .ZN(n317) );
  INV_X2 U780 ( .A(n318), .ZN(n408) );
  INV_X2 U781 ( .A(n309), .ZN(n407) );
  INV_X2 U782 ( .A(n306), .ZN(n304) );
  INV_X2 U783 ( .A(n305), .ZN(n303) );
  INV_X2 U784 ( .A(n300), .ZN(n298) );
  INV_X2 U785 ( .A(n299), .ZN(n297) );
  INV_X2 U786 ( .A(n295), .ZN(n293) );
  INV_X2 U787 ( .A(n294), .ZN(n406) );
  INV_X2 U788 ( .A(n285), .ZN(n405) );
  INV_X2 U789 ( .A(n268), .ZN(n266) );
  INV_X2 U790 ( .A(n267), .ZN(n265) );
  INV_X2 U791 ( .A(n263), .ZN(n261) );
  INV_X2 U792 ( .A(n262), .ZN(n404) );
  INV_X2 U793 ( .A(n253), .ZN(n403) );
  INV_X2 U794 ( .A(n249), .ZN(n247) );
  INV_X2 U795 ( .A(n244), .ZN(n242) );
  INV_X2 U796 ( .A(n243), .ZN(n241) );
  INV_X2 U797 ( .A(n238), .ZN(n402) );
  INV_X2 U798 ( .A(n230), .ZN(n228) );
  INV_X2 U799 ( .A(n229), .ZN(n401) );
  INV_X2 U800 ( .A(n223), .ZN(n221) );
  INV_X2 U801 ( .A(n220), .ZN(n218) );
  INV_X2 U802 ( .A(n219), .ZN(n217) );
  INV_X2 U803 ( .A(n216), .ZN(n214) );
  INV_X2 U804 ( .A(n215), .ZN(n213) );
  INV_X2 U805 ( .A(n211), .ZN(n209) );
  INV_X2 U806 ( .A(n210), .ZN(n400) );
  INV_X2 U807 ( .A(n198), .ZN(n196) );
  INV_X2 U808 ( .A(n197), .ZN(n195) );
  INV_X2 U809 ( .A(n192), .ZN(n190) );
  INV_X2 U810 ( .A(n191), .ZN(n189) );
  INV_X2 U811 ( .A(n187), .ZN(n185) );
  INV_X2 U812 ( .A(n177), .ZN(n397) );
  INV_X2 U813 ( .A(n169), .ZN(n167) );
  INV_X2 U814 ( .A(n165), .ZN(n163) );
  INV_X2 U815 ( .A(n150), .ZN(n148) );
  INV_X2 U816 ( .A(n149), .ZN(n395) );
  INV_X2 U817 ( .A(n142), .ZN(n140) );
  INV_X2 U818 ( .A(n141), .ZN(n139) );
  INV_X2 U819 ( .A(n137), .ZN(n135) );
  INV_X2 U820 ( .A(n136), .ZN(n394) );
  INV_X2 U821 ( .A(n128), .ZN(n126) );
  INV_X2 U822 ( .A(n127), .ZN(n393) );
  INV_X2 U823 ( .A(n112), .ZN(n110) );
  INV_X2 U824 ( .A(n111), .ZN(n109) );
  INV_X2 U825 ( .A(n107), .ZN(n105) );
  INV_X2 U826 ( .A(n106), .ZN(n392) );
endmodule


module up_island_DW01_add_2 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] ;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U1 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  AND2_X1 U2 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  XOR2_X1 U3 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  AND2_X1 U4 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  XOR2_X1 U5 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  AND2_X1 U6 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  XOR2_X1 U7 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  AND2_X1 U8 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  XOR2_X1 U9 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  AND2_X1 U10 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  XOR2_X1 U11 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  AND2_X1 U12 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  XOR2_X1 U13 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  AND2_X1 U14 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  XOR2_X1 U15 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  AND2_X1 U16 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  XOR2_X1 U17 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  AND2_X1 U18 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  XOR2_X1 U19 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  AND2_X1 U20 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  XOR2_X1 U21 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  XOR2_X1 U23 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  AND2_X1 U24 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  XOR2_X1 U25 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  AND2_X1 U26 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  XOR2_X1 U27 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  AND2_X1 U28 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  XOR2_X1 U29 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  AND2_X1 U30 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  XOR2_X1 U31 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  AND2_X1 U32 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  XOR2_X1 U33 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  AND2_X1 U34 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  XOR2_X1 U35 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  AND2_X1 U36 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  XOR2_X1 U37 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  AND2_X1 U38 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  XOR2_X1 U39 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  AND2_X1 U40 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  XOR2_X1 U41 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  INV_X1 U42 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module up_island_DW01_add_1 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \carry[21] , \carry[19] , \carry[18] , \carry[17] , \carry[16] ,
         \carry[15] , \carry[14] , \carry[13] , \carry[12] , \carry[11] ,
         \carry[10] , \carry[9] , \carry[8] , \carry[7] , \carry[6] ,
         \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[1] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130;

  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  INV_X1 U1 ( .A(n114), .ZN(n105) );
  NAND2_X1 U2 ( .A1(\carry[21] ), .A2(A[21]), .ZN(n1) );
  NAND3_X2 U3 ( .A1(n76), .A2(n77), .A3(n78), .ZN(\carry[21] ) );
  AND2_X1 U4 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n121), .A2(n122), .A3(n120), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n121), .A2(n122), .A3(n120), .ZN(\carry[6] ) );
  NAND3_X1 U7 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n4) );
  NAND3_X1 U8 ( .A1(n8), .A2(n10), .A3(n9), .ZN(\carry[7] ) );
  NAND2_X1 U9 ( .A1(n2), .A2(A[1]), .ZN(n5) );
  NAND2_X1 U10 ( .A1(\carry[1] ), .A2(A[1]), .ZN(n84) );
  NAND2_X1 U11 ( .A1(\carry[18] ), .A2(A[18]), .ZN(n65) );
  CLKBUF_X1 U12 ( .A(n3), .Z(n6) );
  XOR2_X1 U13 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR2_X1 U14 ( .A(n6), .B(n7), .Z(SUM[6]) );
  NAND2_X1 U15 ( .A1(n3), .A2(B[6]), .ZN(n8) );
  NAND2_X1 U16 ( .A1(\carry[6] ), .A2(A[6]), .ZN(n9) );
  NAND2_X1 U17 ( .A1(B[6]), .A2(A[6]), .ZN(n10) );
  CLKBUF_X1 U18 ( .A(\carry[17] ), .Z(n11) );
  NAND2_X1 U19 ( .A1(n24), .A2(A[16]), .ZN(n12) );
  NAND3_X1 U20 ( .A1(n43), .A2(n42), .A3(n41), .ZN(n13) );
  NAND3_X1 U21 ( .A1(n109), .A2(n107), .A3(n108), .ZN(n14) );
  NAND3_X1 U22 ( .A1(n70), .A2(n71), .A3(n72), .ZN(n15) );
  CLKBUF_X1 U23 ( .A(\carry[11] ), .Z(n16) );
  CLKBUF_X1 U24 ( .A(n4), .Z(n17) );
  CLKBUF_X1 U25 ( .A(n2), .Z(n18) );
  NAND3_X1 U26 ( .A1(n47), .A2(n46), .A3(n45), .ZN(n19) );
  NAND3_X1 U27 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n47), .A2(n46), .A3(n45), .ZN(\carry[9] ) );
  NAND2_X1 U29 ( .A1(n74), .A2(A[4]), .ZN(n21) );
  NAND2_X1 U30 ( .A1(n87), .A2(A[14]), .ZN(n22) );
  CLKBUF_X1 U31 ( .A(n20), .Z(n23) );
  NAND3_X1 U32 ( .A1(n61), .A2(n60), .A3(n59), .ZN(\carry[13] ) );
  NAND3_X1 U33 ( .A1(n31), .A2(n33), .A3(n32), .ZN(n24) );
  NAND3_X1 U34 ( .A1(n31), .A2(n32), .A3(n33), .ZN(\carry[16] ) );
  NAND3_X1 U35 ( .A1(n22), .A2(n99), .A3(n100), .ZN(n25) );
  CLKBUF_X1 U36 ( .A(n56), .Z(n26) );
  CLKBUF_X1 U37 ( .A(n25), .Z(n27) );
  NAND3_X1 U38 ( .A1(n22), .A2(n99), .A3(n100), .ZN(\carry[15] ) );
  CLKBUF_X1 U39 ( .A(n87), .Z(n28) );
  CLKBUF_X1 U40 ( .A(n57), .Z(n29) );
  AND3_X1 U41 ( .A1(n1), .A2(n91), .A3(n89), .ZN(n35) );
  NAND2_X1 U42 ( .A1(\carry[21] ), .A2(A[21]), .ZN(n90) );
  XOR2_X1 U43 ( .A(B[15]), .B(A[15]), .Z(n30) );
  XOR2_X1 U44 ( .A(n27), .B(n30), .Z(SUM[15]) );
  NAND2_X1 U45 ( .A1(n25), .A2(B[15]), .ZN(n31) );
  NAND2_X1 U46 ( .A1(\carry[15] ), .A2(A[15]), .ZN(n32) );
  NAND2_X1 U47 ( .A1(B[15]), .A2(A[15]), .ZN(n33) );
  NAND2_X1 U48 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n71) );
  CLKBUF_X1 U49 ( .A(n24), .Z(n34) );
  XNOR2_X1 U50 ( .A(n35), .B(n101), .ZN(SUM[22]) );
  XOR2_X2 U51 ( .A(n67), .B(n75), .Z(SUM[20]) );
  NAND3_X1 U52 ( .A1(n90), .A2(n91), .A3(n89), .ZN(n36) );
  CLKBUF_X1 U53 ( .A(n13), .Z(n37) );
  NAND3_X1 U54 ( .A1(n43), .A2(n42), .A3(n41), .ZN(\carry[8] ) );
  CLKBUF_X1 U55 ( .A(n19), .Z(n38) );
  NAND3_X1 U56 ( .A1(n83), .A2(n85), .A3(n84), .ZN(n39) );
  XOR2_X1 U57 ( .A(A[7]), .B(B[7]), .Z(n40) );
  XOR2_X1 U58 ( .A(n40), .B(n17), .Z(SUM[7]) );
  NAND2_X2 U59 ( .A1(A[7]), .A2(B[7]), .ZN(n41) );
  NAND2_X1 U60 ( .A1(n4), .A2(A[7]), .ZN(n42) );
  NAND2_X1 U61 ( .A1(B[7]), .A2(\carry[7] ), .ZN(n43) );
  XOR2_X1 U62 ( .A(A[8]), .B(B[8]), .Z(n44) );
  XOR2_X1 U63 ( .A(n44), .B(n37), .Z(SUM[8]) );
  NAND2_X1 U64 ( .A1(A[8]), .A2(B[8]), .ZN(n45) );
  NAND2_X1 U65 ( .A1(\carry[8] ), .A2(A[8]), .ZN(n46) );
  NAND2_X1 U66 ( .A1(n13), .A2(B[8]), .ZN(n47) );
  XOR2_X1 U67 ( .A(B[9]), .B(A[9]), .Z(n48) );
  XOR2_X1 U68 ( .A(n38), .B(n48), .Z(SUM[9]) );
  NAND2_X1 U69 ( .A1(\carry[9] ), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U70 ( .A1(n19), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U71 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NAND3_X1 U72 ( .A1(n50), .A2(n49), .A3(n51), .ZN(\carry[10] ) );
  NAND3_X1 U73 ( .A1(n55), .A2(n26), .A3(n29), .ZN(n52) );
  NAND3_X1 U74 ( .A1(n57), .A2(n56), .A3(n55), .ZN(\carry[12] ) );
  CLKBUF_X1 U75 ( .A(n39), .Z(n53) );
  NAND3_X1 U76 ( .A1(n83), .A2(n5), .A3(n85), .ZN(\carry[2] ) );
  XOR2_X1 U77 ( .A(A[11]), .B(B[11]), .Z(n54) );
  XOR2_X1 U78 ( .A(n54), .B(n16), .Z(SUM[11]) );
  NAND2_X2 U79 ( .A1(A[11]), .A2(B[11]), .ZN(n55) );
  NAND2_X1 U80 ( .A1(A[11]), .A2(\carry[11] ), .ZN(n56) );
  NAND2_X1 U81 ( .A1(\carry[11] ), .A2(B[11]), .ZN(n57) );
  XOR2_X1 U82 ( .A(A[12]), .B(B[12]), .Z(n58) );
  XOR2_X1 U83 ( .A(n58), .B(n52), .Z(SUM[12]) );
  NAND2_X1 U84 ( .A1(A[12]), .A2(B[12]), .ZN(n59) );
  NAND2_X1 U85 ( .A1(\carry[12] ), .A2(A[12]), .ZN(n60) );
  NAND2_X1 U86 ( .A1(\carry[12] ), .A2(B[12]), .ZN(n61) );
  NAND3_X1 U87 ( .A1(n70), .A2(n72), .A3(n71), .ZN(n62) );
  XOR2_X1 U88 ( .A(B[18]), .B(A[18]), .Z(n63) );
  XOR2_X1 U89 ( .A(\carry[18] ), .B(n63), .Z(SUM[18]) );
  NAND2_X1 U90 ( .A1(\carry[18] ), .A2(B[18]), .ZN(n64) );
  NAND2_X1 U91 ( .A1(B[18]), .A2(A[18]), .ZN(n66) );
  NAND3_X2 U92 ( .A1(n65), .A2(n64), .A3(n66), .ZN(\carry[19] ) );
  NAND3_X2 U93 ( .A1(n130), .A2(n129), .A3(n128), .ZN(\carry[18] ) );
  CLKBUF_X1 U94 ( .A(n15), .Z(n67) );
  NAND3_X1 U95 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n68) );
  XOR2_X1 U96 ( .A(B[19]), .B(A[19]), .Z(n69) );
  XOR2_X1 U97 ( .A(\carry[19] ), .B(n69), .Z(SUM[19]) );
  NAND2_X1 U98 ( .A1(\carry[19] ), .A2(B[19]), .ZN(n70) );
  NAND2_X1 U99 ( .A1(B[19]), .A2(A[19]), .ZN(n72) );
  CLKBUF_X1 U100 ( .A(B[2]), .Z(n73) );
  NAND3_X1 U101 ( .A1(n113), .A2(n112), .A3(n111), .ZN(n74) );
  XOR2_X1 U102 ( .A(B[20]), .B(A[20]), .Z(n75) );
  NAND2_X1 U103 ( .A1(n15), .A2(B[20]), .ZN(n76) );
  NAND2_X1 U104 ( .A1(n62), .A2(A[20]), .ZN(n77) );
  NAND2_X1 U105 ( .A1(B[20]), .A2(A[20]), .ZN(n78) );
  XNOR2_X1 U106 ( .A(n80), .B(n79), .ZN(SUM[23]) );
  INV_X32 U107 ( .A(n105), .ZN(n79) );
  AND3_X2 U108 ( .A1(n103), .A2(n102), .A3(n104), .ZN(n80) );
  CLKBUF_X1 U109 ( .A(n74), .Z(n81) );
  XOR2_X1 U110 ( .A(B[1]), .B(A[1]), .Z(n82) );
  XOR2_X1 U111 ( .A(n18), .B(n82), .Z(SUM[1]) );
  NAND2_X1 U112 ( .A1(\carry[1] ), .A2(B[1]), .ZN(n83) );
  NAND2_X1 U113 ( .A1(B[1]), .A2(A[1]), .ZN(n85) );
  NAND3_X1 U114 ( .A1(n113), .A2(n112), .A3(n111), .ZN(\carry[4] ) );
  CLKBUF_X1 U115 ( .A(n14), .Z(n86) );
  NAND3_X1 U116 ( .A1(n96), .A2(n95), .A3(n97), .ZN(n87) );
  XOR2_X1 U117 ( .A(B[21]), .B(A[21]), .Z(n88) );
  XOR2_X1 U118 ( .A(\carry[21] ), .B(n88), .Z(SUM[21]) );
  NAND2_X1 U119 ( .A1(n68), .A2(B[21]), .ZN(n89) );
  NAND2_X1 U120 ( .A1(B[21]), .A2(A[21]), .ZN(n91) );
  NAND3_X1 U121 ( .A1(n21), .A2(n118), .A3(n117), .ZN(n92) );
  CLKBUF_X1 U122 ( .A(B[0]), .Z(n93) );
  NAND3_X1 U123 ( .A1(n109), .A2(n107), .A3(n108), .ZN(\carry[3] ) );
  NAND3_X1 U124 ( .A1(n96), .A2(n95), .A3(n97), .ZN(\carry[14] ) );
  XOR2_X1 U125 ( .A(A[13]), .B(B[13]), .Z(n94) );
  XOR2_X1 U126 ( .A(n94), .B(n23), .Z(SUM[13]) );
  NAND2_X2 U127 ( .A1(A[13]), .A2(B[13]), .ZN(n95) );
  NAND2_X1 U128 ( .A1(n20), .A2(A[13]), .ZN(n96) );
  NAND2_X1 U129 ( .A1(\carry[13] ), .A2(B[13]), .ZN(n97) );
  XOR2_X1 U130 ( .A(A[14]), .B(B[14]), .Z(n98) );
  XOR2_X1 U131 ( .A(n98), .B(n28), .Z(SUM[14]) );
  NAND2_X1 U132 ( .A1(A[14]), .A2(B[14]), .ZN(n99) );
  NAND2_X1 U133 ( .A1(\carry[14] ), .A2(B[14]), .ZN(n100) );
  XOR2_X1 U134 ( .A(B[22]), .B(A[22]), .Z(n101) );
  NAND2_X1 U135 ( .A1(n36), .A2(B[22]), .ZN(n102) );
  NAND2_X1 U136 ( .A1(n36), .A2(A[22]), .ZN(n103) );
  NAND2_X1 U137 ( .A1(B[22]), .A2(A[22]), .ZN(n104) );
  XOR2_X1 U138 ( .A(A[2]), .B(n73), .Z(n106) );
  XOR2_X1 U139 ( .A(n106), .B(n53), .Z(SUM[2]) );
  NAND2_X1 U140 ( .A1(B[2]), .A2(A[2]), .ZN(n107) );
  NAND2_X1 U141 ( .A1(\carry[2] ), .A2(A[2]), .ZN(n108) );
  NAND2_X1 U142 ( .A1(n39), .A2(B[2]), .ZN(n109) );
  XOR2_X1 U143 ( .A(A[3]), .B(B[3]), .Z(n110) );
  XOR2_X1 U144 ( .A(n110), .B(n86), .Z(SUM[3]) );
  NAND2_X1 U145 ( .A1(A[3]), .A2(B[3]), .ZN(n111) );
  NAND2_X1 U146 ( .A1(\carry[3] ), .A2(A[3]), .ZN(n112) );
  NAND2_X1 U147 ( .A1(n14), .A2(B[3]), .ZN(n113) );
  XOR2_X1 U148 ( .A(B[23]), .B(A[23]), .Z(n114) );
  CLKBUF_X1 U149 ( .A(n92), .Z(n115) );
  NAND3_X1 U150 ( .A1(n21), .A2(n117), .A3(n118), .ZN(\carry[5] ) );
  XOR2_X1 U151 ( .A(A[4]), .B(B[4]), .Z(n116) );
  XOR2_X1 U152 ( .A(n116), .B(n81), .Z(SUM[4]) );
  NAND2_X1 U153 ( .A1(A[4]), .A2(B[4]), .ZN(n117) );
  NAND2_X1 U154 ( .A1(B[4]), .A2(\carry[4] ), .ZN(n118) );
  XOR2_X1 U155 ( .A(A[5]), .B(B[5]), .Z(n119) );
  XOR2_X1 U156 ( .A(n119), .B(n115), .Z(SUM[5]) );
  NAND2_X1 U157 ( .A1(A[5]), .A2(B[5]), .ZN(n120) );
  NAND2_X1 U158 ( .A1(n92), .A2(A[5]), .ZN(n121) );
  NAND2_X1 U159 ( .A1(\carry[5] ), .A2(B[5]), .ZN(n122) );
  NAND3_X1 U160 ( .A1(n12), .A2(n126), .A3(n125), .ZN(n123) );
  NAND3_X1 U161 ( .A1(n12), .A2(n126), .A3(n125), .ZN(\carry[17] ) );
  XOR2_X1 U162 ( .A(A[16]), .B(B[16]), .Z(n124) );
  XOR2_X1 U163 ( .A(n124), .B(n34), .Z(SUM[16]) );
  NAND2_X2 U164 ( .A1(A[16]), .A2(B[16]), .ZN(n125) );
  NAND2_X1 U165 ( .A1(\carry[16] ), .A2(B[16]), .ZN(n126) );
  XOR2_X1 U166 ( .A(A[17]), .B(B[17]), .Z(n127) );
  XOR2_X1 U167 ( .A(n127), .B(n11), .Z(SUM[17]) );
  NAND2_X1 U168 ( .A1(A[17]), .A2(B[17]), .ZN(n128) );
  NAND2_X1 U169 ( .A1(A[17]), .A2(n123), .ZN(n129) );
  NAND2_X1 U170 ( .A1(\carry[17] ), .A2(B[17]), .ZN(n130) );
  AND2_X2 U171 ( .A1(B[0]), .A2(A[0]), .ZN(\carry[1] ) );
  XOR2_X1 U172 ( .A(n93), .B(A[0]), .Z(SUM[0]) );
endmodule


module up_island ( CLK, reset, BUS_NREADY, BUS_BUSY, BUS_MR, BUS_MW, 
        BUS_ADDR_OUTBUS, BUS_DATA_INBUS, BUS_DATA_OUTBUS );
  output [31:0] BUS_ADDR_OUTBUS;
  input [31:0] BUS_DATA_INBUS;
  output [31:0] BUS_DATA_OUTBUS;
  input CLK, reset, BUS_NREADY;
  output BUS_BUSY, BUS_MR, BUS_MW;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, I_BUSY,
         dmem_read, dmem_write, dmem_isbyte, dmem_ishalf, iram_rd, N19, N20,
         N21, N22, N24, N25, N26, N27, N29, N30, N31, N33, N34, N35, N37, N38,
         N40, N41, N42, N43, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, \UUT/N77 , \UUT/N76 ,
         \UUT/m_mem_command[SIGN] , \UUT/m_mem_command[MR] , \UUT/m_we ,
         \UUT/x_we , \UUT/Alu_command[OP][0] , \UUT/Alu_command[OP][1] ,
         \UUT/Alu_command[OP][2] , \UUT/Alu_command[OP][3] ,
         \UUT/Alu_command[OP][4] , \UUT/Alu_command[OP][5] ,
         \UUT/byp_controlB[0] , \UUT/byp_controlB[2] , \UUT/byp_controlA[0] ,
         \UUT/byp_controlA[2] , \UUT/break_code[0] , \UUT/break_code[1] ,
         \UUT/break_code[4] , \UUT/break_code[5] , \UUT/break_code[6] ,
         \UUT/break_code[7] , \UUT/break_code[8] , \UUT/break_code[9] ,
         \UUT/break_code[10] , \UUT/break_code[11] , \UUT/break_code[12] ,
         \UUT/break_code[13] , \UUT/break_code[14] , \UUT/break_code[15] ,
         \UUT/break_code[16] , \UUT/break_code[17] , \UUT/break_code[18] ,
         \UUT/break_code[19] , \UUT/break_code[20] , \UUT/break_code[21] ,
         \UUT/break_code[22] , \UUT/break_code[23] , \UUT/N3 ,
         \UUT/regfile/N457 , \UUT/regfile/N456 , \UUT/regfile/N455 ,
         \UUT/regfile/N451 , \UUT/regfile/N450 , \UUT/regfile/N445 ,
         \UUT/regfile/N444 , \UUT/regfile/N439 , \UUT/regfile/N438 ,
         \UUT/regfile/N433 , \UUT/regfile/N432 , \UUT/regfile/N427 ,
         \UUT/regfile/N426 , \UUT/regfile/N421 , \UUT/regfile/N420 ,
         \UUT/regfile/N415 , \UUT/regfile/N414 , \UUT/regfile/N409 ,
         \UUT/regfile/N408 , \UUT/regfile/N403 , \UUT/regfile/N402 ,
         \UUT/regfile/N397 , \UUT/regfile/N396 , \UUT/regfile/N391 ,
         \UUT/regfile/N390 , \UUT/regfile/N385 , \UUT/regfile/N384 ,
         \UUT/regfile/N379 , \UUT/regfile/N378 , \UUT/regfile/N373 ,
         \UUT/regfile/N372 , \UUT/regfile/N367 , \UUT/regfile/N366 ,
         \UUT/regfile/N360 , \UUT/regfile/N359 , \UUT/regfile/N358 ,
         \UUT/regfile/N354 , \UUT/regfile/N353 , \UUT/regfile/N348 ,
         \UUT/regfile/N347 , \UUT/regfile/N342 , \UUT/regfile/N341 ,
         \UUT/regfile/N336 , \UUT/regfile/N335 , \UUT/regfile/N330 ,
         \UUT/regfile/N329 , \UUT/regfile/N324 , \UUT/regfile/N323 ,
         \UUT/regfile/N318 , \UUT/regfile/N317 , \UUT/regfile/N315 ,
         \UUT/regfile/N311 , \UUT/regfile/N310 , \UUT/regfile/N305 ,
         \UUT/regfile/N304 , \UUT/regfile/N299 , \UUT/regfile/N298 ,
         \UUT/regfile/N293 , \UUT/regfile/N292 , \UUT/regfile/N290 ,
         \UUT/regfile/N286 , \UUT/regfile/N285 , \UUT/regfile/N280 ,
         \UUT/regfile/N279 , \UUT/regfile/N273 , \UUT/regfile/N272 ,
         \UUT/regfile/N269 , \UUT/regfile/N267 , \UUT/regfile/N266 ,
         \UUT/regfile/N265 , \UUT/regfile/N262 , \UUT/regfile/N261 ,
         \UUT/regfile/N260 , \UUT/regfile/reg_out[18][0] ,
         \UUT/regfile/reg_out[18][1] , \UUT/regfile/reg_out[18][2] ,
         \UUT/regfile/reg_out[18][3] , \UUT/regfile/reg_out[18][4] ,
         \UUT/regfile/reg_out[18][5] , \UUT/regfile/reg_out[18][6] ,
         \UUT/regfile/reg_out[18][7] , \UUT/regfile/reg_out[18][8] ,
         \UUT/regfile/reg_out[18][9] , \UUT/regfile/reg_out[18][10] ,
         \UUT/regfile/reg_out[18][11] , \UUT/regfile/reg_out[18][12] ,
         \UUT/regfile/reg_out[18][13] , \UUT/regfile/reg_out[18][14] ,
         \UUT/regfile/reg_out[18][15] , \UUT/regfile/reg_out[18][16] ,
         \UUT/regfile/reg_out[18][17] , \UUT/regfile/reg_out[18][18] ,
         \UUT/regfile/reg_out[18][19] , \UUT/regfile/reg_out[18][20] ,
         \UUT/regfile/reg_out[18][21] , \UUT/regfile/reg_out[18][22] ,
         \UUT/regfile/reg_out[18][23] , \UUT/regfile/reg_out[18][24] ,
         \UUT/regfile/reg_out[18][25] , \UUT/regfile/reg_out[18][26] ,
         \UUT/regfile/reg_out[18][27] , \UUT/regfile/reg_out[18][28] ,
         \UUT/regfile/reg_out[18][29] , \UUT/regfile/reg_out[18][30] ,
         \UUT/regfile/reg_out[18][31] , \UUT/regfile/reg_out[19][0] ,
         \UUT/regfile/reg_out[19][1] , \UUT/regfile/reg_out[19][2] ,
         \UUT/regfile/reg_out[19][3] , \UUT/regfile/reg_out[19][4] ,
         \UUT/regfile/reg_out[19][5] , \UUT/regfile/reg_out[19][6] ,
         \UUT/regfile/reg_out[19][7] , \UUT/regfile/reg_out[19][8] ,
         \UUT/regfile/reg_out[19][9] , \UUT/regfile/reg_out[19][10] ,
         \UUT/regfile/reg_out[19][11] , \UUT/regfile/reg_out[19][12] ,
         \UUT/regfile/reg_out[19][13] , \UUT/regfile/reg_out[19][14] ,
         \UUT/regfile/reg_out[19][15] , \UUT/regfile/reg_out[19][16] ,
         \UUT/regfile/reg_out[19][17] , \UUT/regfile/reg_out[19][18] ,
         \UUT/regfile/reg_out[19][19] , \UUT/regfile/reg_out[19][20] ,
         \UUT/regfile/reg_out[19][21] , \UUT/regfile/reg_out[19][22] ,
         \UUT/regfile/reg_out[19][23] , \UUT/regfile/reg_out[19][24] ,
         \UUT/regfile/reg_out[19][25] , \UUT/regfile/reg_out[19][26] ,
         \UUT/regfile/reg_out[19][27] , \UUT/regfile/reg_out[19][28] ,
         \UUT/regfile/reg_out[19][29] , \UUT/regfile/reg_out[19][30] ,
         \UUT/regfile/reg_out[19][31] , \UUT/regfile/reg_out[20][0] ,
         \UUT/regfile/reg_out[20][1] , \UUT/regfile/reg_out[20][2] ,
         \UUT/regfile/reg_out[20][3] , \UUT/regfile/reg_out[20][4] ,
         \UUT/regfile/reg_out[20][5] , \UUT/regfile/reg_out[20][6] ,
         \UUT/regfile/reg_out[20][7] , \UUT/regfile/reg_out[20][8] ,
         \UUT/regfile/reg_out[20][9] , \UUT/regfile/reg_out[20][10] ,
         \UUT/regfile/reg_out[20][11] , \UUT/regfile/reg_out[20][12] ,
         \UUT/regfile/reg_out[20][13] , \UUT/regfile/reg_out[20][14] ,
         \UUT/regfile/reg_out[20][15] , \UUT/regfile/reg_out[20][16] ,
         \UUT/regfile/reg_out[20][17] , \UUT/regfile/reg_out[20][18] ,
         \UUT/regfile/reg_out[20][19] , \UUT/regfile/reg_out[20][20] ,
         \UUT/regfile/reg_out[20][21] , \UUT/regfile/reg_out[20][22] ,
         \UUT/regfile/reg_out[20][23] , \UUT/regfile/reg_out[20][24] ,
         \UUT/regfile/reg_out[20][25] , \UUT/regfile/reg_out[20][26] ,
         \UUT/regfile/reg_out[20][27] , \UUT/regfile/reg_out[20][28] ,
         \UUT/regfile/reg_out[20][29] , \UUT/regfile/reg_out[20][30] ,
         \UUT/regfile/reg_out[20][31] , \UUT/regfile/reg_out[21][0] ,
         \UUT/regfile/reg_out[21][1] , \UUT/regfile/reg_out[21][2] ,
         \UUT/regfile/reg_out[21][3] , \UUT/regfile/reg_out[21][4] ,
         \UUT/regfile/reg_out[21][5] , \UUT/regfile/reg_out[21][6] ,
         \UUT/regfile/reg_out[21][7] , \UUT/regfile/reg_out[21][8] ,
         \UUT/regfile/reg_out[21][9] , \UUT/regfile/reg_out[21][10] ,
         \UUT/regfile/reg_out[21][11] , \UUT/regfile/reg_out[21][12] ,
         \UUT/regfile/reg_out[21][13] , \UUT/regfile/reg_out[21][14] ,
         \UUT/regfile/reg_out[21][15] , \UUT/regfile/reg_out[21][16] ,
         \UUT/regfile/reg_out[21][17] , \UUT/regfile/reg_out[21][18] ,
         \UUT/regfile/reg_out[21][19] , \UUT/regfile/reg_out[21][20] ,
         \UUT/regfile/reg_out[21][21] , \UUT/regfile/reg_out[21][22] ,
         \UUT/regfile/reg_out[21][23] , \UUT/regfile/reg_out[21][24] ,
         \UUT/regfile/reg_out[21][25] , \UUT/regfile/reg_out[21][26] ,
         \UUT/regfile/reg_out[21][27] , \UUT/regfile/reg_out[21][28] ,
         \UUT/regfile/reg_out[21][29] , \UUT/regfile/reg_out[21][30] ,
         \UUT/regfile/reg_out[21][31] , \UUT/regfile/reg_out[24][0] ,
         \UUT/regfile/reg_out[24][1] , \UUT/regfile/reg_out[24][2] ,
         \UUT/regfile/reg_out[24][3] , \UUT/regfile/reg_out[24][4] ,
         \UUT/regfile/reg_out[24][5] , \UUT/regfile/reg_out[24][6] ,
         \UUT/regfile/reg_out[24][7] , \UUT/regfile/reg_out[24][8] ,
         \UUT/regfile/reg_out[24][9] , \UUT/regfile/reg_out[24][10] ,
         \UUT/regfile/reg_out[24][11] , \UUT/regfile/reg_out[24][12] ,
         \UUT/regfile/reg_out[24][13] , \UUT/regfile/reg_out[24][14] ,
         \UUT/regfile/reg_out[24][15] , \UUT/regfile/reg_out[24][16] ,
         \UUT/regfile/reg_out[24][17] , \UUT/regfile/reg_out[24][18] ,
         \UUT/regfile/reg_out[24][19] , \UUT/regfile/reg_out[24][20] ,
         \UUT/regfile/reg_out[24][21] , \UUT/regfile/reg_out[24][22] ,
         \UUT/regfile/reg_out[24][23] , \UUT/regfile/reg_out[24][24] ,
         \UUT/regfile/reg_out[24][25] , \UUT/regfile/reg_out[24][26] ,
         \UUT/regfile/reg_out[24][27] , \UUT/regfile/reg_out[24][28] ,
         \UUT/regfile/reg_out[24][29] , \UUT/regfile/reg_out[24][30] ,
         \UUT/regfile/reg_out[24][31] , \UUT/regfile/reg_out[25][0] ,
         \UUT/regfile/reg_out[25][1] , \UUT/regfile/reg_out[25][2] ,
         \UUT/regfile/reg_out[25][3] , \UUT/regfile/reg_out[25][4] ,
         \UUT/regfile/reg_out[25][5] , \UUT/regfile/reg_out[25][6] ,
         \UUT/regfile/reg_out[25][7] , \UUT/regfile/reg_out[25][8] ,
         \UUT/regfile/reg_out[25][9] , \UUT/regfile/reg_out[25][10] ,
         \UUT/regfile/reg_out[25][11] , \UUT/regfile/reg_out[25][12] ,
         \UUT/regfile/reg_out[25][13] , \UUT/regfile/reg_out[25][14] ,
         \UUT/regfile/reg_out[25][15] , \UUT/regfile/reg_out[25][16] ,
         \UUT/regfile/reg_out[25][17] , \UUT/regfile/reg_out[25][18] ,
         \UUT/regfile/reg_out[25][19] , \UUT/regfile/reg_out[25][20] ,
         \UUT/regfile/reg_out[25][21] , \UUT/regfile/reg_out[25][22] ,
         \UUT/regfile/reg_out[25][23] , \UUT/regfile/reg_out[25][24] ,
         \UUT/regfile/reg_out[25][25] , \UUT/regfile/reg_out[25][26] ,
         \UUT/regfile/reg_out[25][27] , \UUT/regfile/reg_out[25][28] ,
         \UUT/regfile/reg_out[25][29] , \UUT/regfile/reg_out[25][30] ,
         \UUT/regfile/reg_out[25][31] , \UUT/regfile/reg_out[28][0] ,
         \UUT/regfile/reg_out[28][1] , \UUT/regfile/reg_out[28][2] ,
         \UUT/regfile/reg_out[28][3] , \UUT/regfile/reg_out[28][4] ,
         \UUT/regfile/reg_out[28][5] , \UUT/regfile/reg_out[28][6] ,
         \UUT/regfile/reg_out[28][7] , \UUT/regfile/reg_out[28][8] ,
         \UUT/regfile/reg_out[28][9] , \UUT/regfile/reg_out[28][10] ,
         \UUT/regfile/reg_out[28][11] , \UUT/regfile/reg_out[28][12] ,
         \UUT/regfile/reg_out[28][13] , \UUT/regfile/reg_out[28][14] ,
         \UUT/regfile/reg_out[28][15] , \UUT/regfile/reg_out[28][16] ,
         \UUT/regfile/reg_out[28][17] , \UUT/regfile/reg_out[28][18] ,
         \UUT/regfile/reg_out[28][19] , \UUT/regfile/reg_out[28][20] ,
         \UUT/regfile/reg_out[28][21] , \UUT/regfile/reg_out[28][22] ,
         \UUT/regfile/reg_out[28][23] , \UUT/regfile/reg_out[28][24] ,
         \UUT/regfile/reg_out[28][25] , \UUT/regfile/reg_out[28][26] ,
         \UUT/regfile/reg_out[28][27] , \UUT/regfile/reg_out[28][28] ,
         \UUT/regfile/reg_out[28][29] , \UUT/regfile/reg_out[28][30] ,
         \UUT/regfile/reg_out[28][31] , \UUT/regfile/reg_out[29][0] ,
         \UUT/regfile/reg_out[29][1] , \UUT/regfile/reg_out[29][2] ,
         \UUT/regfile/reg_out[29][3] , \UUT/regfile/reg_out[29][4] ,
         \UUT/regfile/reg_out[29][5] , \UUT/regfile/reg_out[29][6] ,
         \UUT/regfile/reg_out[29][7] , \UUT/regfile/reg_out[29][8] ,
         \UUT/regfile/reg_out[29][9] , \UUT/regfile/reg_out[29][10] ,
         \UUT/regfile/reg_out[29][11] , \UUT/regfile/reg_out[29][12] ,
         \UUT/regfile/reg_out[29][13] , \UUT/regfile/reg_out[29][14] ,
         \UUT/regfile/reg_out[29][15] , \UUT/regfile/reg_out[29][16] ,
         \UUT/regfile/reg_out[29][17] , \UUT/regfile/reg_out[29][18] ,
         \UUT/regfile/reg_out[29][19] , \UUT/regfile/reg_out[29][20] ,
         \UUT/regfile/reg_out[29][21] , \UUT/regfile/reg_out[29][22] ,
         \UUT/regfile/reg_out[29][23] , \UUT/regfile/reg_out[29][24] ,
         \UUT/regfile/reg_out[29][25] , \UUT/regfile/reg_out[29][26] ,
         \UUT/regfile/reg_out[29][27] , \UUT/regfile/reg_out[29][28] ,
         \UUT/regfile/reg_out[29][29] , \UUT/regfile/reg_out[29][30] ,
         \UUT/regfile/reg_out[29][31] , \UUT/regfile/reg_out[4][0] ,
         \UUT/regfile/reg_out[4][1] , \UUT/regfile/reg_out[4][2] ,
         \UUT/regfile/reg_out[4][3] , \UUT/regfile/reg_out[4][4] ,
         \UUT/regfile/reg_out[4][5] , \UUT/regfile/reg_out[4][6] ,
         \UUT/regfile/reg_out[4][7] , \UUT/regfile/reg_out[4][8] ,
         \UUT/regfile/reg_out[4][9] , \UUT/regfile/reg_out[4][10] ,
         \UUT/regfile/reg_out[4][11] , \UUT/regfile/reg_out[4][12] ,
         \UUT/regfile/reg_out[4][13] , \UUT/regfile/reg_out[4][14] ,
         \UUT/regfile/reg_out[4][15] , \UUT/regfile/reg_out[4][16] ,
         \UUT/regfile/reg_out[4][17] , \UUT/regfile/reg_out[4][18] ,
         \UUT/regfile/reg_out[4][19] , \UUT/regfile/reg_out[4][20] ,
         \UUT/regfile/reg_out[4][21] , \UUT/regfile/reg_out[4][22] ,
         \UUT/regfile/reg_out[4][23] , \UUT/regfile/reg_out[4][24] ,
         \UUT/regfile/reg_out[4][25] , \UUT/regfile/reg_out[4][26] ,
         \UUT/regfile/reg_out[4][27] , \UUT/regfile/reg_out[4][28] ,
         \UUT/regfile/reg_out[4][29] , \UUT/regfile/reg_out[4][30] ,
         \UUT/regfile/reg_out[4][31] , \UUT/regfile/reg_out[5][0] ,
         \UUT/regfile/reg_out[5][1] , \UUT/regfile/reg_out[5][2] ,
         \UUT/regfile/reg_out[5][3] , \UUT/regfile/reg_out[5][4] ,
         \UUT/regfile/reg_out[5][5] , \UUT/regfile/reg_out[5][6] ,
         \UUT/regfile/reg_out[5][7] , \UUT/regfile/reg_out[5][8] ,
         \UUT/regfile/reg_out[5][9] , \UUT/regfile/reg_out[5][10] ,
         \UUT/regfile/reg_out[5][11] , \UUT/regfile/reg_out[5][12] ,
         \UUT/regfile/reg_out[5][13] , \UUT/regfile/reg_out[5][14] ,
         \UUT/regfile/reg_out[5][15] , \UUT/regfile/reg_out[5][16] ,
         \UUT/regfile/reg_out[5][17] , \UUT/regfile/reg_out[5][18] ,
         \UUT/regfile/reg_out[5][19] , \UUT/regfile/reg_out[5][20] ,
         \UUT/regfile/reg_out[5][21] , \UUT/regfile/reg_out[5][22] ,
         \UUT/regfile/reg_out[5][23] , \UUT/regfile/reg_out[5][24] ,
         \UUT/regfile/reg_out[5][25] , \UUT/regfile/reg_out[5][26] ,
         \UUT/regfile/reg_out[5][27] , \UUT/regfile/reg_out[5][28] ,
         \UUT/regfile/reg_out[5][29] , \UUT/regfile/reg_out[5][30] ,
         \UUT/regfile/reg_out[5][31] , \UUT/BYP_BRANCH_MUXB/N39 ,
         \UUT/BYP_BRANCH_MUXB/N4 , \UUT/Mcontrol/N22 , \UUT/Mcontrol/N19 ,
         \UUT/Mcontrol/x_sampled_dmem_command[SIGN] ,
         \UUT/Mcontrol/x_sampled_dmem_command[MW] ,
         \UUT/Mcontrol/m_sampled_xrd[0] , \UUT/Mcontrol/m_sampled_xrd[1] ,
         \UUT/Mcontrol/m_sampled_xrd[2] , \UUT/Mcontrol/m_sampled_xrd[3] ,
         \UUT/Mcontrol/m_sampled_xrd[4] , \UUT/Mcontrol/x_rd[0] ,
         \UUT/Mcontrol/x_rd[1] , \UUT/Mcontrol/x_rd[2] ,
         \UUT/Mcontrol/x_rd[3] , \UUT/Mcontrol/x_rd[4] ,
         \UUT/Mcontrol/d_jump_type[0] , \UUT/Mcontrol/d_jump_type[1] ,
         \UUT/Mcontrol/d_jump_type[2] , \UUT/Mcontrol/d_jump_type[3] ,
         \UUT/Mcontrol/int_reset , \UUT/Mcontrol/Program_counter/N28 ,
         \UUT/Mcontrol/Program_counter/N26 ,
         \UUT/Mcontrol/Program_counter/N24 ,
         \UUT/Mcontrol/Program_counter/N22 ,
         \UUT/Mcontrol/Program_counter/N20 ,
         \UUT/Mcontrol/Program_counter/N18 ,
         \UUT/Mcontrol/Program_counter/N16 ,
         \UUT/Mcontrol/Program_counter/N14 ,
         \UUT/Mcontrol/Program_counter/N12 ,
         \UUT/Mcontrol/Program_counter/N10 , \UUT/Mcontrol/Program_counter/N8 ,
         \UUT/Mcontrol/Operation_decoding32/N2088 ,
         \UUT/Mcontrol/Operation_decoding32/N2085 ,
         \UUT/Mcontrol/Operation_decoding32/N2084 ,
         \UUT/Mcontrol/Operation_decoding32/N2083 ,
         \UUT/Mcontrol/Operation_decoding32/N2082 ,
         \UUT/Mcontrol/Operation_decoding32/N2081 ,
         \UUT/Mcontrol/Operation_decoding32/N2079 ,
         \UUT/Mcontrol/Operation_decoding32/N2071 ,
         \UUT/Mcontrol/Operation_decoding32/N2066 ,
         \UUT/Mcontrol/Operation_decoding32/N2060 ,
         \UUT/Mcontrol/Operation_decoding32/N2057 ,
         \UUT/Mcontrol/Operation_decoding32/N2056 ,
         \UUT/Mcontrol/Operation_decoding32/N2054 ,
         \UUT/Mcontrol/Operation_decoding32/N2050 ,
         \UUT/Mcontrol/Operation_decoding32/N2047 ,
         \UUT/Mcontrol/Operation_decoding32/N2043 ,
         \UUT/Mcontrol/Operation_decoding32/N2027 ,
         \UUT/Mcontrol/Operation_decoding32/N2025 ,
         \UUT/Mcontrol/Operation_decoding32/N2023 ,
         \UUT/Mcontrol/Operation_decoding32/N2017 ,
         \UUT/Mcontrol/Operation_decoding32/N2016 ,
         \UUT/Mcontrol/Operation_decoding32/N2015 ,
         \UUT/Mcontrol/Operation_decoding32/N2009 ,
         \UUT/Mcontrol/Operation_decoding32/N2008 ,
         \UUT/Mcontrol/Operation_decoding32/N2007 ,
         \UUT/Mcontrol/Operation_decoding32/N2005 ,
         \UUT/Mcontrol/Operation_decoding32/N2002 ,
         \UUT/Mcontrol/Operation_decoding32/N2001 ,
         \UUT/Mcontrol/Operation_decoding32/N1999 ,
         \UUT/Mcontrol/Operation_decoding32/N1995 ,
         \UUT/Mcontrol/Operation_decoding32/N1994 ,
         \UUT/Mcontrol/Operation_decoding32/N1989 ,
         \UUT/Mcontrol/Operation_decoding32/N1987 ,
         \UUT/Mcontrol/Operation_decoding32/N1985 ,
         \UUT/Mcontrol/Operation_decoding32/N1984 ,
         \UUT/Mcontrol/Operation_decoding32/N1981 ,
         \UUT/Mcontrol/Operation_decoding32/N1979 ,
         \UUT/Mcontrol/Operation_decoding32/N1978 ,
         \UUT/Mcontrol/Operation_decoding32/N1977 ,
         \UUT/Mcontrol/Operation_decoding32/N1973 ,
         \UUT/Mcontrol/Operation_decoding32/N1965 ,
         \UUT/Mcontrol/Operation_decoding32/N1962 ,
         \UUT/Mcontrol/Operation_decoding32/N1958 ,
         \UUT/Mcontrol/Operation_decoding32/N1957 ,
         \UUT/Mcontrol/Operation_decoding32/N1956 ,
         \UUT/Mcontrol/Operation_decoding32/N1955 ,
         \UUT/Mcontrol/Operation_decoding32/N1952 ,
         \UUT/Mcontrol/Operation_decoding32/N1951 ,
         \UUT/Mcontrol/Operation_decoding32/N1950 ,
         \UUT/Mcontrol/Operation_decoding32/N1947 ,
         \UUT/Mcontrol/Operation_decoding32/N1946 ,
         \UUT/Mcontrol/Operation_decoding32/N1945 ,
         \UUT/Mcontrol/Operation_decoding32/N1940 ,
         \UUT/Mcontrol/Operation_decoding32/N1934 ,
         \UUT/Mcontrol/Operation_decoding32/N1933 ,
         \UUT/Mcontrol/Operation_decoding32/N1932 ,
         \UUT/Mcontrol/Operation_decoding32/N1928 ,
         \UUT/Mcontrol/Operation_decoding32/N1927 ,
         \UUT/Mcontrol/Operation_decoding32/N1924 ,
         \UUT/Mcontrol/Operation_decoding32/N1923 ,
         \UUT/Mcontrol/Operation_decoding32/N1922 ,
         \UUT/Mcontrol/Operation_decoding32/N1921 ,
         \UUT/Mcontrol/Operation_decoding32/N1919 ,
         \UUT/Mcontrol/Operation_decoding32/N1918 ,
         \UUT/Mcontrol/Operation_decoding32/N1917 ,
         \UUT/Mcontrol/Operation_decoding32/N1916 ,
         \UUT/Mcontrol/Operation_decoding32/N1915 ,
         \UUT/Mcontrol/Operation_decoding32/N1914 ,
         \UUT/Mcontrol/Operation_decoding32/N1913 ,
         \UUT/Mcontrol/Operation_decoding32/N1912 ,
         \UUT/Mcontrol/Operation_decoding32/N1911 ,
         \UUT/Mcontrol/Operation_decoding32/N1910 ,
         \UUT/Mcontrol/Operation_decoding32/N1909 ,
         \UUT/Mcontrol/Operation_decoding32/N1908 ,
         \UUT/Mcontrol/Operation_decoding32/N1907 ,
         \UUT/Mcontrol/Operation_decoding32/N1906 ,
         \UUT/Mcontrol/Operation_decoding32/N1905 ,
         \UUT/Mcontrol/Operation_decoding32/N1904 ,
         \UUT/Mcontrol/Operation_decoding32/N1903 ,
         \UUT/Mcontrol/Operation_decoding32/N1902 ,
         \UUT/Mcontrol/Operation_decoding32/N1901 ,
         \UUT/Mcontrol/Operation_decoding32/N1900 ,
         \UUT/Mcontrol/Operation_decoding32/N1899 ,
         \UUT/Mcontrol/Operation_decoding32/N1898 ,
         \UUT/Mcontrol/Operation_decoding32/N1897 ,
         \UUT/Mcontrol/Operation_decoding32/N1896 ,
         \UUT/Mcontrol/Operation_decoding32/N1895 ,
         \UUT/Mcontrol/Operation_decoding32/N1894 ,
         \UUT/Mcontrol/Operation_decoding32/N1893 ,
         \UUT/Mcontrol/Operation_decoding32/N1892 ,
         \UUT/Mcontrol/Operation_decoding32/N1891 ,
         \UUT/Mcontrol/Operation_decoding32/N1890 ,
         \UUT/Mcontrol/Operation_decoding32/N1889 ,
         \UUT/Mcontrol/Operation_decoding32/N1884 ,
         \UUT/Mcontrol/Operation_decoding32/N1883 ,
         \UUT/Mcontrol/Operation_decoding32/N1882 ,
         \UUT/Mcontrol/Operation_decoding32/N1877 ,
         \UUT/Mcontrol/Operation_decoding32/N1873 ,
         \UUT/Mcontrol/Operation_decoding32/N1871 ,
         \UUT/Mcontrol/Operation_decoding32/N62 ,
         \UUT/Mcontrol/Nextpc_decoding/N266 ,
         \UUT/Mcontrol/Nextpc_decoding/N265 ,
         \UUT/Mcontrol/Nextpc_decoding/N264 ,
         \UUT/Mcontrol/Nextpc_decoding/N263 ,
         \UUT/Mcontrol/Nextpc_decoding/N262 ,
         \UUT/Mcontrol/Nextpc_decoding/N260 ,
         \UUT/Mcontrol/Nextpc_decoding/N259 ,
         \UUT/Mcontrol/Nextpc_decoding/N258 ,
         \UUT/Mcontrol/Nextpc_decoding/N257 ,
         \UUT/Mcontrol/Nextpc_decoding/N256 ,
         \UUT/Mcontrol/Nextpc_decoding/N254 ,
         \UUT/Mcontrol/Nextpc_decoding/N253 ,
         \UUT/Mcontrol/Nextpc_decoding/N252 ,
         \UUT/Mcontrol/Nextpc_decoding/N251 ,
         \UUT/Mcontrol/Nextpc_decoding/N250 ,
         \UUT/Mcontrol/Nextpc_decoding/N248 ,
         \UUT/Mcontrol/Nextpc_decoding/N247 ,
         \UUT/Mcontrol/Nextpc_decoding/N246 ,
         \UUT/Mcontrol/Nextpc_decoding/N245 ,
         \UUT/Mcontrol/Nextpc_decoding/N244 ,
         \UUT/Mcontrol/Nextpc_decoding/N242 ,
         \UUT/Mcontrol/Nextpc_decoding/N241 ,
         \UUT/Mcontrol/Nextpc_decoding/N240 ,
         \UUT/Mcontrol/Nextpc_decoding/N239 ,
         \UUT/Mcontrol/Nextpc_decoding/N238 ,
         \UUT/Mcontrol/Nextpc_decoding/N236 ,
         \UUT/Mcontrol/Nextpc_decoding/N235 ,
         \UUT/Mcontrol/Nextpc_decoding/N234 ,
         \UUT/Mcontrol/Nextpc_decoding/N233 ,
         \UUT/Mcontrol/Nextpc_decoding/N232 ,
         \UUT/Mcontrol/Nextpc_decoding/N230 ,
         \UUT/Mcontrol/Nextpc_decoding/N229 ,
         \UUT/Mcontrol/Nextpc_decoding/N228 ,
         \UUT/Mcontrol/Nextpc_decoding/N227 ,
         \UUT/Mcontrol/Nextpc_decoding/N226 ,
         \UUT/Mcontrol/Nextpc_decoding/N224 ,
         \UUT/Mcontrol/Nextpc_decoding/N223 ,
         \UUT/Mcontrol/Nextpc_decoding/N205 ,
         \UUT/Mcontrol/Nextpc_decoding/N200 ,
         \UUT/Mcontrol/Nextpc_decoding/N194 ,
         \UUT/Mcontrol/Nextpc_decoding/N159 ,
         \UUT/Mcontrol/Nextpc_decoding/N142 ,
         \UUT/Mcontrol/Nextpc_decoding/N141 ,
         \UUT/Mcontrol/Nextpc_decoding/N140 ,
         \UUT/Mcontrol/Nextpc_decoding/N139 ,
         \UUT/Mcontrol/Nextpc_decoding/N138 ,
         \UUT/Mcontrol/Nextpc_decoding/N137 ,
         \UUT/Mcontrol/Nextpc_decoding/N134 ,
         \UUT/Mcontrol/Nextpc_decoding/N127 ,
         \UUT/Mcontrol/Nextpc_decoding/N125 ,
         \UUT/Mcontrol/Nextpc_decoding/N124 ,
         \UUT/Mcontrol/Nextpc_decoding/N123 ,
         \UUT/Mcontrol/Nextpc_decoding/N122 ,
         \UUT/Mcontrol/Nextpc_decoding/N120 ,
         \UUT/Mcontrol/Nextpc_decoding/N116 ,
         \UUT/Mcontrol/Nextpc_decoding/N115 ,
         \UUT/Mcontrol/Nextpc_decoding/N114 ,
         \UUT/Mcontrol/Nextpc_decoding/N32 ,
         \UUT/Mcontrol/Nextpc_decoding/N27 ,
         \UUT/Mcontrol/Nextpc_decoding/N25 ,
         \UUT/Mcontrol/Nextpc_decoding/condition ,
         \UUT/Mcontrol/Nextpc_decoding/N22 , \UUT/Mcontrol/bp_logicA/N16 ,
         \UUT/Mcontrol/bp_logicA/N15 , \UUT/Mcontrol/bp_logicA/N14 ,
         \UUT/Mcontrol/bp_logicA/N13 , \UUT/Mcontrol/bp_logicA/N12 ,
         \UUT/Mcontrol/bp_logicA/N11 , \UUT/Mcontrol/bp_logicA/N10 ,
         \UUT/Mcontrol/bp_logicA/N9 , \UUT/Mcontrol/bp_logicA/N8 ,
         \UUT/Mcontrol/bp_logicA/N7 , \UUT/Mcontrol/bp_logicA/N6 ,
         \UUT/Mcontrol/bp_logicA/N5 , \UUT/Mcontrol/bp_logicA/memory_main ,
         \UUT/Mcontrol/bp_logicA/N3 , \UUT/Mcontrol/bp_logicA/exec_main ,
         \UUT/Mcontrol/bp_logicA/N2 , \UUT/Mcontrol/bp_logicB/N16 ,
         \UUT/Mcontrol/bp_logicB/N15 , \UUT/Mcontrol/bp_logicB/N14 ,
         \UUT/Mcontrol/bp_logicB/N13 , \UUT/Mcontrol/bp_logicB/N12 ,
         \UUT/Mcontrol/bp_logicB/N11 , \UUT/Mcontrol/bp_logicB/N10 ,
         \UUT/Mcontrol/bp_logicB/N9 , \UUT/Mcontrol/bp_logicB/N8 ,
         \UUT/Mcontrol/bp_logicB/N7 , \UUT/Mcontrol/bp_logicB/N6 ,
         \UUT/Mcontrol/bp_logicB/N5 , \UUT/Mcontrol/bp_logicB/memory_main ,
         \UUT/Mcontrol/bp_logicB/N3 , \UUT/Mcontrol/bp_logicB/exec_main ,
         \UUT/Mcontrol/bp_logicB/N2 , \UUT/Mcontrol/st_logic/N120 ,
         \UUT/Mcontrol/st_logic/N119 , \UUT/Mcontrol/st_logic/N118 ,
         \UUT/Mcontrol/st_logic/N117 , \UUT/Mcontrol/st_logic/N112 ,
         \UUT/Mcontrol/st_logic/N111 , \UUT/Mcontrol/st_logic/N110 ,
         \UUT/Mcontrol/st_logic/N108 , \UUT/Mcontrol/st_logic/N107 ,
         \UUT/Mcontrol/st_logic/N106 , \UUT/Mcontrol/st_logic/N105 ,
         \UUT/Mcontrol/st_logic/N104 , \UUT/Mcontrol/st_logic/N103 ,
         \UUT/Mcontrol/st_logic/N101 , \UUT/Mcontrol/st_logic/N100 ,
         \UUT/Mcontrol/st_logic/N99 , \UUT/Mcontrol/st_logic/N98 ,
         \UUT/Mcontrol/st_logic/N96 , \UUT/Mcontrol/st_logic/N95 ,
         \UUT/Mcontrol/st_logic/N94 , \UUT/Mcontrol/st_logic/N93 ,
         \UUT/Mcontrol/st_logic/N92 , \UUT/Mcontrol/st_logic/N90 ,
         \UUT/Mcontrol/st_logic/N89 , \UUT/Mcontrol/st_logic/N88 ,
         \UUT/Mcontrol/st_logic/N87 , \UUT/Mcontrol/st_logic/N86 ,
         \UUT/Mcontrol/st_logic/N85 , \UUT/Mcontrol/st_logic/N83 ,
         \UUT/Mcontrol/st_logic/N82 , \UUT/Mcontrol/st_logic/N81 ,
         \UUT/Mcontrol/st_logic/N80 , \UUT/Mcontrol/st_logic/N79 ,
         \UUT/Mcontrol/st_logic/N77 , \UUT/Mcontrol/st_logic/N76 ,
         \UUT/Mcontrol/st_logic/N75 , \UUT/Mcontrol/st_logic/N74 ,
         \UUT/Mcontrol/st_logic/N73 , \UUT/Mcontrol/st_logic/N71 ,
         \UUT/Mcontrol/st_logic/N70 , \UUT/Mcontrol/st_logic/N69 ,
         \UUT/Mcontrol/st_logic/N68 , \UUT/Mcontrol/st_logic/N67 ,
         \UUT/Mcontrol/st_logic/N65 , \UUT/Mcontrol/st_logic/N64 ,
         \UUT/Mcontrol/st_logic/N63 , \UUT/Mcontrol/st_logic/N62 ,
         \UUT/Mcontrol/st_logic/N61 , \UUT/Mcontrol/st_logic/N60 ,
         \UUT/Mcontrol/st_logic/N58 , \UUT/Mcontrol/st_logic/N57 ,
         \UUT/Mcontrol/st_logic/N56 , \UUT/Mcontrol/st_logic/N55 ,
         \UUT/Mcontrol/st_logic/N54 , \UUT/Mcontrol/st_logic/N53 ,
         \UUT/Mcontrol/st_logic/N52 , \UUT/Mcontrol/st_logic/N51 ,
         \UUT/Mcontrol/st_logic/N50 , \UUT/Mcontrol/st_logic/N49 ,
         \UUT/Mcontrol/st_logic/N47 , \UUT/Mcontrol/st_logic/N46 ,
         \UUT/Mcontrol/st_logic/N45 , \UUT/Mcontrol/st_logic/N44 ,
         \UUT/Mcontrol/st_logic/N42 , \UUT/Mcontrol/st_logic/N41 ,
         \UUT/Mcontrol/st_logic/N40 , \UUT/Mcontrol/st_logic/N39 ,
         \UUT/Mcontrol/st_logic/N38 , \UUT/Mcontrol/st_logic/N37 ,
         \UUT/Mcontrol/st_logic/N36 , \UUT/Mcontrol/st_logic/N35 ,
         \UUT/Mcontrol/st_logic/N34 , \UUT/Mcontrol/st_logic/N33 ,
         \UUT/Mcontrol/st_logic/N32 , \UUT/Mcontrol/st_logic/N31 ,
         \UUT/Mcontrol/st_logic/N30 , \UUT/Mcontrol/st_logic/N29 ,
         \UUT/Mcontrol/st_logic/N28 , \UUT/Mcontrol/st_logic/N27 ,
         \UUT/Mcontrol/st_logic/N26 , \UUT/Mcontrol/st_logic/N25 ,
         \UUT/Mcontrol/st_logic/N24 , \UUT/Mcontrol/st_logic/N23 ,
         \UUT/Mcontrol/st_logic/N22 , \UUT/Mcontrol/st_logic/N19 ,
         \UUT/Mcontrol/st_logic/N18 , \UUT/Mcontrol/st_logic/N15 ,
         \UUT/Mcontrol/st_logic/N14 , \UUT/Mcontrol/st_logic/N13 ,
         \UUT/Mcontrol/st_logic/N12 , \UUT/Mcontrol/st_logic/N10 ,
         \UUT/Mcontrol/st_logic/branchmul_stall , \UUT/Mcontrol/st_logic/N8 ,
         \UUT/Mcontrol/st_logic/branch_uses_main_exe_result ,
         \UUT/Mcontrol/st_logic/N7 , \UUT/Mcontrol/st_logic/branchlw_stall ,
         \UUT/Mcontrol/st_logic/N6 , \UUT/Mcontrol/st_logic/branch_uses_regb ,
         \UUT/Mcontrol/st_logic/N4 , \UUT/Mcontrol/st_logic/load_stall ,
         \UUT/Mcontrol/st_logic/N2 , \UUT/Mpath/N128 , \UUT/Mpath/N127 ,
         \UUT/Mpath/N125 , \UUT/Mpath/N124 , \UUT/Mpath/N121 ,
         \UUT/Mpath/N119 , \UUT/Mpath/N118 , \UUT/Mpath/N117 ,
         \UUT/Mpath/N116 , \UUT/Mpath/N115 , \UUT/Mpath/N114 ,
         \UUT/Mpath/N113 , \UUT/Mpath/N112 , \UUT/Mpath/N111 ,
         \UUT/Mpath/out_regB[0] , \UUT/Mpath/out_regB[1] ,
         \UUT/Mpath/out_regB[2] , \UUT/Mpath/out_regB[3] ,
         \UUT/Mpath/out_regB[4] , \UUT/Mpath/out_regB[5] ,
         \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[7] ,
         \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[9] ,
         \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[11] ,
         \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[13] ,
         \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[15] ,
         \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[17] ,
         \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[19] ,
         \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[21] ,
         \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[23] ,
         \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[25] ,
         \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[27] ,
         \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[29] ,
         \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[31] ,
         \UUT/Mpath/out_regA[0] , \UUT/Mpath/out_regA[1] ,
         \UUT/Mpath/out_regA[2] , \UUT/Mpath/out_regA[3] ,
         \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[5] ,
         \UUT/Mpath/out_regA[6] , \UUT/Mpath/out_regA[7] ,
         \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[9] ,
         \UUT/Mpath/out_regA[10] , \UUT/Mpath/out_regA[11] ,
         \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[13] ,
         \UUT/Mpath/out_regA[14] , \UUT/Mpath/out_regA[15] ,
         \UUT/Mpath/out_regA[16] , \UUT/Mpath/out_regA[17] ,
         \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[19] ,
         \UUT/Mpath/out_regA[20] , \UUT/Mpath/out_regA[21] ,
         \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[23] ,
         \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[25] ,
         \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[27] ,
         \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[29] ,
         \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[31] ,
         \UUT/Mpath/the_alu/N526 , \UUT/Mpath/the_alu/N525 ,
         \UUT/Mpath/the_alu/N524 , \UUT/Mpath/the_alu/N523 ,
         \UUT/Mpath/the_alu/N520 , \UUT/Mpath/the_alu/N519 ,
         \UUT/Mpath/the_alu/N518 , \UUT/Mpath/the_alu/N517 ,
         \UUT/Mpath/the_alu/N515 , \UUT/Mpath/the_alu/N514 ,
         \UUT/Mpath/the_alu/N513 , \UUT/Mpath/the_alu/N512 ,
         \UUT/Mpath/the_alu/N511 , \UUT/Mpath/the_alu/N509 ,
         \UUT/Mpath/the_alu/N508 , \UUT/Mpath/the_alu/N507 ,
         \UUT/Mpath/the_alu/N506 , \UUT/Mpath/the_alu/N505 ,
         \UUT/Mpath/the_alu/N503 , \UUT/Mpath/the_alu/N502 ,
         \UUT/Mpath/the_alu/N501 , \UUT/Mpath/the_alu/N500 ,
         \UUT/Mpath/the_alu/N499 , \UUT/Mpath/the_alu/N498 ,
         \UUT/Mpath/the_alu/N497 , \UUT/Mpath/the_alu/N496 ,
         \UUT/Mpath/the_alu/N495 , \UUT/Mpath/the_alu/N494 ,
         \UUT/Mpath/the_alu/N493 , \UUT/Mpath/the_alu/N492 ,
         \UUT/Mpath/the_alu/N491 , \UUT/Mpath/the_alu/N490 ,
         \UUT/Mpath/the_alu/N489 , \UUT/Mpath/the_alu/N488 ,
         \UUT/Mpath/the_alu/N487 , \UUT/Mpath/the_alu/N486 ,
         \UUT/Mpath/the_alu/N485 , \UUT/Mpath/the_alu/N484 ,
         \UUT/Mpath/the_alu/N483 , \UUT/Mpath/the_alu/N482 ,
         \UUT/Mpath/the_alu/N481 , \UUT/Mpath/the_alu/N480 ,
         \UUT/Mpath/the_alu/N479 , \UUT/Mpath/the_alu/N478 ,
         \UUT/Mpath/the_alu/N477 , \UUT/Mpath/the_alu/N476 ,
         \UUT/Mpath/the_alu/N475 , \UUT/Mpath/the_alu/N474 ,
         \UUT/Mpath/the_alu/N473 , \UUT/Mpath/the_alu/N472 ,
         \UUT/Mpath/the_alu/N471 , \UUT/Mpath/the_alu/N470 ,
         \UUT/Mpath/the_alu/N469 , \UUT/Mpath/the_alu/N468 ,
         \UUT/Mpath/the_alu/N467 , \UUT/Mpath/the_alu/N466 ,
         \UUT/Mpath/the_alu/N453 , \UUT/Mpath/the_alu/N221 ,
         \UUT/Mpath/the_alu/N219 , \UUT/Mpath/the_alu/N218 ,
         \UUT/Mpath/the_alu/N217 , \UUT/Mpath/the_alu/N216 ,
         \UUT/Mpath/the_alu/N215 , \UUT/Mpath/the_alu/N214 ,
         \UUT/Mpath/the_alu/N213 , \UUT/Mpath/the_alu/N212 ,
         \UUT/Mpath/the_alu/N211 , \UUT/Mpath/the_alu/N210 ,
         \UUT/Mpath/the_alu/N209 , \UUT/Mpath/the_alu/N208 ,
         \UUT/Mpath/the_alu/N207 , \UUT/Mpath/the_alu/N206 ,
         \UUT/Mpath/the_alu/N205 , \UUT/Mpath/the_alu/N204 ,
         \UUT/Mpath/the_alu/N203 , \UUT/Mpath/the_alu/N202 ,
         \UUT/Mpath/the_alu/N201 , \UUT/Mpath/the_alu/N200 ,
         \UUT/Mpath/the_alu/N199 , \UUT/Mpath/the_alu/N198 ,
         \UUT/Mpath/the_alu/N189 , \UUT/Mpath/the_alu/N187 ,
         \UUT/Mpath/the_alu/N186 , \UUT/Mpath/the_alu/N185 ,
         \UUT/Mpath/the_alu/N184 , \UUT/Mpath/the_alu/N183 ,
         \UUT/Mpath/the_alu/N182 , \UUT/Mpath/the_alu/N181 ,
         \UUT/Mpath/the_alu/N180 , \UUT/Mpath/the_alu/N179 ,
         \UUT/Mpath/the_alu/N178 , \UUT/Mpath/the_alu/N177 ,
         \UUT/Mpath/the_alu/N176 , \UUT/Mpath/the_alu/N175 ,
         \UUT/Mpath/the_alu/N174 , \UUT/Mpath/the_alu/N173 ,
         \UUT/Mpath/the_alu/N172 , \UUT/Mpath/the_alu/N171 ,
         \UUT/Mpath/the_alu/N170 , \UUT/Mpath/the_alu/N169 ,
         \UUT/Mpath/the_alu/N168 , \UUT/Mpath/the_alu/N167 ,
         \UUT/Mpath/the_alu/N166 , \UUT/Mpath/the_alu/N157 ,
         \UUT/Mpath/the_alu/N155 , \UUT/Mpath/the_alu/N154 ,
         \UUT/Mpath/the_alu/N153 , \UUT/Mpath/the_alu/N152 ,
         \UUT/Mpath/the_alu/N151 , \UUT/Mpath/the_alu/N150 ,
         \UUT/Mpath/the_alu/N149 , \UUT/Mpath/the_alu/N148 ,
         \UUT/Mpath/the_alu/N147 , \UUT/Mpath/the_alu/N146 ,
         \UUT/Mpath/the_alu/N145 , \UUT/Mpath/the_alu/N144 ,
         \UUT/Mpath/the_alu/N143 , \UUT/Mpath/the_alu/N142 ,
         \UUT/Mpath/the_alu/N141 , \UUT/Mpath/the_alu/N140 ,
         \UUT/Mpath/the_alu/N139 , \UUT/Mpath/the_alu/N138 ,
         \UUT/Mpath/the_alu/N137 , \UUT/Mpath/the_alu/N136 ,
         \UUT/Mpath/the_alu/N135 , \UUT/Mpath/the_alu/N134 ,
         \UUT/Mpath/the_alu/N125 , \UUT/Mpath/the_alu/N123 ,
         \UUT/Mpath/the_alu/N122 , \UUT/Mpath/the_alu/N121 ,
         \UUT/Mpath/the_alu/N120 , \UUT/Mpath/the_alu/N119 ,
         \UUT/Mpath/the_alu/N118 , \UUT/Mpath/the_alu/N117 ,
         \UUT/Mpath/the_alu/N116 , \UUT/Mpath/the_alu/N115 ,
         \UUT/Mpath/the_alu/N114 , \UUT/Mpath/the_alu/N113 ,
         \UUT/Mpath/the_alu/N112 , \UUT/Mpath/the_alu/N111 ,
         \UUT/Mpath/the_alu/N110 , \UUT/Mpath/the_alu/N109 ,
         \UUT/Mpath/the_alu/N108 , \UUT/Mpath/the_alu/N107 ,
         \UUT/Mpath/the_alu/N106 , \UUT/Mpath/the_alu/N105 ,
         \UUT/Mpath/the_alu/N104 , \UUT/Mpath/the_alu/N103 ,
         \UUT/Mpath/the_alu/N102 , \UUT/Mpath/the_alu/N93 ,
         \UUT/Mpath/the_alu/N91 , \UUT/Mpath/the_alu/diff[0] ,
         \UUT/Mpath/the_alu/diff[1] , \UUT/Mpath/the_alu/diff[2] ,
         \UUT/Mpath/the_alu/diff[3] , \UUT/Mpath/the_alu/diff[4] ,
         \UUT/Mpath/the_alu/diff[5] , \UUT/Mpath/the_alu/diff[6] ,
         \UUT/Mpath/the_alu/diff[7] , \UUT/Mpath/the_alu/diff[8] ,
         \UUT/Mpath/the_alu/diff[9] , \UUT/Mpath/the_alu/diff[10] ,
         \UUT/Mpath/the_alu/diff[11] , \UUT/Mpath/the_alu/diff[12] ,
         \UUT/Mpath/the_alu/diff[13] , \UUT/Mpath/the_alu/diff[14] ,
         \UUT/Mpath/the_alu/diff[15] , \UUT/Mpath/the_alu/diff[16] ,
         \UUT/Mpath/the_alu/diff[17] , \UUT/Mpath/the_alu/diff[18] ,
         \UUT/Mpath/the_alu/diff[19] , \UUT/Mpath/the_alu/diff[20] ,
         \UUT/Mpath/the_alu/diff[21] , \UUT/Mpath/the_alu/diff[22] ,
         \UUT/Mpath/the_alu/diff[23] , \UUT/Mpath/the_alu/diff[24] ,
         \UUT/Mpath/the_alu/diff[25] , \UUT/Mpath/the_alu/diff[26] ,
         \UUT/Mpath/the_alu/diff[27] , \UUT/Mpath/the_alu/diff[28] ,
         \UUT/Mpath/the_alu/diff[29] , \UUT/Mpath/the_alu/diff[30] ,
         \UUT/Mpath/the_alu/diff[31] , \UUT/Mpath/the_alu/sum[0] ,
         \UUT/Mpath/the_alu/sum[1] , \UUT/Mpath/the_alu/sum[2] ,
         \UUT/Mpath/the_alu/sum[3] , \UUT/Mpath/the_alu/sum[4] ,
         \UUT/Mpath/the_alu/sum[5] , \UUT/Mpath/the_alu/sum[6] ,
         \UUT/Mpath/the_alu/sum[7] , \UUT/Mpath/the_alu/sum[8] ,
         \UUT/Mpath/the_alu/sum[9] , \UUT/Mpath/the_alu/sum[10] ,
         \UUT/Mpath/the_alu/sum[11] , \UUT/Mpath/the_alu/sum[12] ,
         \UUT/Mpath/the_alu/sum[13] , \UUT/Mpath/the_alu/sum[14] ,
         \UUT/Mpath/the_alu/sum[15] , \UUT/Mpath/the_alu/sum[16] ,
         \UUT/Mpath/the_alu/sum[17] , \UUT/Mpath/the_alu/sum[18] ,
         \UUT/Mpath/the_alu/sum[19] , \UUT/Mpath/the_alu/sum[20] ,
         \UUT/Mpath/the_alu/sum[21] , \UUT/Mpath/the_alu/sum[22] ,
         \UUT/Mpath/the_alu/sum[23] , \UUT/Mpath/the_alu/sum[24] ,
         \UUT/Mpath/the_alu/sum[25] , \UUT/Mpath/the_alu/sum[26] ,
         \UUT/Mpath/the_alu/sum[27] , \UUT/Mpath/the_alu/sum[28] ,
         \UUT/Mpath/the_alu/sum[29] , \UUT/Mpath/the_alu/sum[30] ,
         \UUT/Mpath/the_alu/sum[31] , \UUT/Mpath/the_alu/N84 ,
         \UUT/Mpath/the_alu/N83 , \UUT/Mpath/the_alu/N82 ,
         \UUT/Mpath/the_alu/N81 , \UUT/Mpath/the_alu/N80 ,
         \UUT/Mpath/the_alu/N79 , \UUT/Mpath/the_alu/N78 ,
         \UUT/Mpath/the_alu/N77 , \UUT/Mpath/the_alu/N76 ,
         \UUT/Mpath/the_alu/N75 , \UUT/Mpath/the_alu/N74 ,
         \UUT/Mpath/the_alu/N73 , \UUT/Mpath/the_alu/N72 ,
         \UUT/Mpath/the_alu/N71 , \UUT/Mpath/the_alu/N70 ,
         \UUT/Mpath/the_alu/N69 , \UUT/Mpath/the_alu/N68 ,
         \UUT/Mpath/the_alu/N67 , \UUT/Mpath/the_alu/N66 ,
         \UUT/Mpath/the_alu/N65 , \UUT/Mpath/the_alu/N64 ,
         \UUT/Mpath/the_alu/N63 , \UUT/Mpath/the_alu/N62 ,
         \UUT/Mpath/the_alu/N61 , \UUT/Mpath/the_alu/N60 ,
         \UUT/Mpath/the_alu/N59 , \UUT/Mpath/the_alu/N58 ,
         \UUT/Mpath/the_alu/N57 , \UUT/Mpath/the_alu/N56 ,
         \UUT/Mpath/the_alu/N55 , \UUT/Mpath/the_alu/N54 ,
         \UUT/Mpath/the_alu/N53 , \UUT/Mpath/the_alu/N52 ,
         \UUT/Mpath/the_alu/N51 , \UUT/Mpath/the_alu/N50 ,
         \UUT/Mpath/the_alu/N49 , \UUT/Mpath/the_alu/N48 ,
         \UUT/Mpath/the_alu/N47 , \UUT/Mpath/the_alu/N46 ,
         \UUT/Mpath/the_alu/N45 , \UUT/Mpath/the_alu/N44 ,
         \UUT/Mpath/the_alu/N43 , \UUT/Mpath/the_alu/N42 ,
         \UUT/Mpath/the_alu/N41 , \UUT/Mpath/the_alu/N40 ,
         \UUT/Mpath/the_alu/N39 , \UUT/Mpath/the_alu/N38 ,
         \UUT/Mpath/the_alu/N37 , \UUT/Mpath/the_alu/N36 ,
         \UUT/Mpath/the_alu/N35 , \UUT/Mpath/the_alu/N34 ,
         \UUT/Mpath/the_alu/N33 , \UUT/Mpath/the_alu/N32 ,
         \UUT/Mpath/the_alu/N31 , \UUT/Mpath/the_alu/N30 ,
         \UUT/Mpath/the_alu/N29 , \UUT/Mpath/the_alu/N28 ,
         \UUT/Mpath/the_alu/N27 , \UUT/Mpath/the_alu/N26 ,
         \UUT/Mpath/the_alu/N25 , \UUT/Mpath/the_alu/N24 ,
         \UUT/Mpath/the_alu/N23 , \UUT/Mpath/the_alu/N22 ,
         \UUT/Mpath/the_alu/N21 , \UUT/Mpath/the_shift/N118 ,
         \UUT/Mpath/the_shift/N117 , \UUT/Mpath/the_shift/N116 ,
         \UUT/Mpath/the_shift/N115 , \UUT/Mpath/the_shift/N114 ,
         \UUT/Mpath/the_shift/N113 , \UUT/Mpath/the_shift/N112 ,
         \UUT/Mpath/the_shift/N111 , \UUT/Mpath/the_shift/N110 ,
         \UUT/Mpath/the_shift/N109 , \UUT/Mpath/the_shift/N107 ,
         \UUT/Mpath/the_shift/N106 , \UUT/Mpath/the_shift/N105 ,
         \UUT/Mpath/the_shift/N104 , \UUT/Mpath/the_mult/N314 ,
         \UUT/Mpath/the_mult/N313 , \UUT/Mpath/the_mult/N312 ,
         \UUT/Mpath/the_mult/N311 , \UUT/Mpath/the_mult/N310 ,
         \UUT/Mpath/the_mult/N309 , \UUT/Mpath/the_mult/N308 ,
         \UUT/Mpath/the_mult/N307 , \UUT/Mpath/the_mult/N306 ,
         \UUT/Mpath/the_mult/N305 , \UUT/Mpath/the_mult/N304 ,
         \UUT/Mpath/the_mult/N303 , \UUT/Mpath/the_mult/N302 ,
         \UUT/Mpath/the_mult/N301 , \UUT/Mpath/the_mult/N300 ,
         \UUT/Mpath/the_mult/N299 , \UUT/Mpath/the_mult/N298 ,
         \UUT/Mpath/the_mult/N297 , \UUT/Mpath/the_mult/N296 ,
         \UUT/Mpath/the_mult/N295 , \UUT/Mpath/the_mult/N294 ,
         \UUT/Mpath/the_mult/N293 , \UUT/Mpath/the_mult/N292 ,
         \UUT/Mpath/the_mult/N291 , \UUT/Mpath/the_mult/N290 ,
         \UUT/Mpath/the_mult/N289 , \UUT/Mpath/the_mult/N288 ,
         \UUT/Mpath/the_mult/N287 , \UUT/Mpath/the_mult/N285 ,
         \UUT/Mpath/the_mult/N284 , \UUT/Mpath/the_mult/N283 ,
         \UUT/Mpath/the_mult/N282 , \UUT/Mpath/the_mult/N281 ,
         \UUT/Mpath/the_mult/N280 , \UUT/Mpath/the_mult/N279 ,
         \UUT/Mpath/the_mult/N278 , \UUT/Mpath/the_mult/N277 ,
         \UUT/Mpath/the_mult/N276 , \UUT/Mpath/the_mult/N275 ,
         \UUT/Mpath/the_mult/N274 , \UUT/Mpath/the_mult/N273 ,
         \UUT/Mpath/the_mult/N272 , \UUT/Mpath/the_mult/N271 ,
         \UUT/Mpath/the_mult/N270 , \UUT/Mpath/the_mult/N269 ,
         \UUT/Mpath/the_mult/N268 , \UUT/Mpath/the_mult/N267 ,
         \UUT/Mpath/the_mult/N266 , \UUT/Mpath/the_mult/N265 ,
         \UUT/Mpath/the_mult/N264 , \UUT/Mpath/the_mult/N263 ,
         \UUT/Mpath/the_mult/N262 , \UUT/Mpath/the_mult/N261 ,
         \UUT/Mpath/the_mult/N260 , \UUT/Mpath/the_mult/N259 ,
         \UUT/Mpath/the_mult/N258 , \UUT/Mpath/the_mult/N257 ,
         \UUT/Mpath/the_mult/N255 , \UUT/Mpath/the_mult/N254 ,
         \UUT/Mpath/the_mult/N253 , \UUT/Mpath/the_mult/N252 ,
         \UUT/Mpath/the_mult/N251 , \UUT/Mpath/the_mult/N244 ,
         \UUT/Mpath/the_mult/N231 , \UUT/Mpath/the_mult/N230 ,
         \UUT/Mpath/the_mult/N229 , \UUT/Mpath/the_mult/N227 ,
         \UUT/Mpath/the_mult/N226 , \UUT/Mpath/the_mult/N225 ,
         \UUT/Mpath/the_mult/N224 , \UUT/Mpath/the_mult/N223 ,
         \UUT/Mpath/the_mult/N222 , \UUT/Mpath/the_mult/N221 ,
         \UUT/Mpath/the_mult/N220 , \UUT/Mpath/the_mult/N216 ,
         \UUT/Mpath/the_mult/N215 , \UUT/Mpath/the_mult/N214 ,
         \UUT/Mpath/the_mult/N213 , \UUT/Mpath/the_mult/N212 ,
         \UUT/Mpath/the_mult/N198 , \UUT/Mpath/the_mult/N197 ,
         \UUT/Mpath/the_mult/N196 , \UUT/Mpath/the_mult/N195 ,
         \UUT/Mpath/the_mult/N194 , \UUT/Mpath/the_mult/N193 ,
         \UUT/Mpath/the_mult/N192 , \UUT/Mpath/the_mult/acc_out[0] ,
         \UUT/Mpath/the_mult/acc_out[1] , \UUT/Mpath/the_mult/acc_out[2] ,
         \UUT/Mpath/the_mult/acc_out[3] , \UUT/Mpath/the_mult/acc_out[4] ,
         \UUT/Mpath/the_mult/acc_out[5] , \UUT/Mpath/the_mult/acc_out[6] ,
         \UUT/Mpath/the_mult/acc_out[7] , \UUT/Mpath/the_mult/acc_out[8] ,
         \UUT/Mpath/the_mult/acc_out[9] , \UUT/Mpath/the_mult/acc_out[10] ,
         \UUT/Mpath/the_mult/acc_out[11] , \UUT/Mpath/the_mult/acc_out[12] ,
         \UUT/Mpath/the_mult/acc_out[13] , \UUT/Mpath/the_mult/acc_out[14] ,
         \UUT/Mpath/the_mult/acc_out[15] , \UUT/Mpath/the_mult/acc_out[16] ,
         \UUT/Mpath/the_mult/acc_out[17] , \UUT/Mpath/the_mult/acc_out[18] ,
         \UUT/Mpath/the_mult/acc_out[19] , \UUT/Mpath/the_mult/acc_out[20] ,
         \UUT/Mpath/the_mult/acc_out[21] , \UUT/Mpath/the_mult/acc_out[22] ,
         \UUT/Mpath/the_mult/acc_out[23] , \UUT/Mpath/the_mult/acc_out[24] ,
         \UUT/Mpath/the_mult/acc_out[25] , \UUT/Mpath/the_mult/acc_out[26] ,
         \UUT/Mpath/the_mult/acc_out[27] , \UUT/Mpath/the_mult/acc_out[28] ,
         \UUT/Mpath/the_mult/acc_out[29] , \UUT/Mpath/the_mult/acc_out[30] ,
         \UUT/Mpath/the_mult/acc_out[31] , \UUT/Mpath/the_mult/acc_out[32] ,
         \UUT/Mpath/the_mult/acc_out[33] , \UUT/Mpath/the_mult/acc_out[34] ,
         \UUT/Mpath/the_mult/acc_out[35] , \UUT/Mpath/the_mult/acc_out[36] ,
         \UUT/Mpath/the_mult/acc_out[37] , \UUT/Mpath/the_mult/acc_out[38] ,
         \UUT/Mpath/the_mult/acc_out[39] , \UUT/Mpath/the_mult/acc_out[40] ,
         \UUT/Mpath/the_mult/acc_out[41] , \UUT/Mpath/the_mult/acc_out[42] ,
         \UUT/Mpath/the_mult/acc_out[43] , \UUT/Mpath/the_mult/acc_out[44] ,
         \UUT/Mpath/the_mult/acc_out[45] , \UUT/Mpath/the_mult/acc_out[46] ,
         \UUT/Mpath/the_mult/acc_out[47] , \UUT/Mpath/the_mult/acc_out[48] ,
         \UUT/Mpath/the_mult/acc_out[49] , \UUT/Mpath/the_mult/acc_out[50] ,
         \UUT/Mpath/the_mult/acc_out[51] , \UUT/Mpath/the_mult/acc_out[52] ,
         \UUT/Mpath/the_mult/acc_out[53] , \UUT/Mpath/the_mult/acc_out[54] ,
         \UUT/Mpath/the_mult/acc_out[55] , \UUT/Mpath/the_mult/acc_out[56] ,
         \UUT/Mpath/the_mult/acc_out[57] , \UUT/Mpath/the_mult/acc_out[58] ,
         \UUT/Mpath/the_mult/acc_out[59] , \UUT/Mpath/the_mult/acc_out[60] ,
         \UUT/Mpath/the_mult/acc_out[61] , \UUT/Mpath/the_mult/acc_out[62] ,
         \UUT/Mpath/the_mult/acc_out[63] , \UUT/Mpath/the_mult/Mult_out[0] ,
         \UUT/Mpath/the_mult/Mult_out[1] , \UUT/Mpath/the_mult/Mult_out[2] ,
         \UUT/Mpath/the_mult/Mult_out[3] , \UUT/Mpath/the_mult/Mult_out[4] ,
         \UUT/Mpath/the_mult/Mult_out[5] , \UUT/Mpath/the_mult/Mult_out[6] ,
         \UUT/Mpath/the_mult/Mult_out[7] , \UUT/Mpath/the_mult/Mult_out[8] ,
         \UUT/Mpath/the_mult/Mult_out[9] , \UUT/Mpath/the_mult/Mult_out[10] ,
         \UUT/Mpath/the_mult/Mult_out[11] , \UUT/Mpath/the_mult/Mult_out[12] ,
         \UUT/Mpath/the_mult/Mult_out[13] , \UUT/Mpath/the_mult/Mult_out[14] ,
         \UUT/Mpath/the_mult/Mult_out[15] , \UUT/Mpath/the_mult/Mult_out[16] ,
         \UUT/Mpath/the_mult/Mult_out[17] , \UUT/Mpath/the_mult/Mult_out[18] ,
         \UUT/Mpath/the_mult/Mult_out[19] , \UUT/Mpath/the_mult/Mult_out[20] ,
         \UUT/Mpath/the_mult/Mult_out[21] , \UUT/Mpath/the_mult/Mult_out[22] ,
         \UUT/Mpath/the_mult/Mult_out[23] , \UUT/Mpath/the_mult/Mult_out[24] ,
         \UUT/Mpath/the_mult/Mult_out[25] , \UUT/Mpath/the_mult/Mult_out[26] ,
         \UUT/Mpath/the_mult/Mult_out[27] , \UUT/Mpath/the_mult/Mult_out[28] ,
         \UUT/Mpath/the_mult/Mult_out[29] , \UUT/Mpath/the_mult/Mult_out[30] ,
         \UUT/Mpath/the_mult/Mult_out[31] , \UUT/Mpath/the_mult/Mult_out[32] ,
         \UUT/Mpath/the_mult/Mult_out[33] , \UUT/Mpath/the_mult/Mult_out[34] ,
         \UUT/Mpath/the_mult/Mult_out[35] , \UUT/Mpath/the_mult/Mult_out[36] ,
         \UUT/Mpath/the_mult/Mult_out[37] , \UUT/Mpath/the_mult/Mult_out[38] ,
         \UUT/Mpath/the_mult/Mult_out[39] , \UUT/Mpath/the_mult/Mult_out[40] ,
         \UUT/Mpath/the_mult/Mult_out[41] , \UUT/Mpath/the_mult/Mult_out[42] ,
         \UUT/Mpath/the_mult/Mult_out[43] , \UUT/Mpath/the_mult/Mult_out[44] ,
         \UUT/Mpath/the_mult/Mult_out[45] , \UUT/Mpath/the_mult/Mult_out[46] ,
         \UUT/Mpath/the_mult/Mult_out[47] , \UUT/Mpath/the_mult/Mult_out[48] ,
         \UUT/Mpath/the_mult/Mult_out[49] , \UUT/Mpath/the_mult/Mult_out[50] ,
         \UUT/Mpath/the_mult/Mult_out[51] , \UUT/Mpath/the_mult/Mult_out[52] ,
         \UUT/Mpath/the_mult/Mult_out[53] , \UUT/Mpath/the_mult/Mult_out[54] ,
         \UUT/Mpath/the_mult/Mult_out[55] , \UUT/Mpath/the_mult/Mult_out[56] ,
         \UUT/Mpath/the_mult/Mult_out[57] , \UUT/Mpath/the_mult/Mult_out[58] ,
         \UUT/Mpath/the_mult/Mult_out[59] , \UUT/Mpath/the_mult/Mult_out[60] ,
         \UUT/Mpath/the_mult/Mult_out[61] , \UUT/Mpath/the_mult/Mult_out[62] ,
         \UUT/Mpath/the_mult/Mult_out[63] ,
         \UUT/Mpath/the_mult/m_mul_command[0] ,
         \UUT/Mpath/the_mult/m_mul_command[1] ,
         \UUT/Mpath/the_mult/m_mul_command[2] ,
         \UUT/Mpath/the_mult/m_mul_command[3] ,
         \UUT/Mpath/the_mult/m_mul_command[4] ,
         \UUT/Mpath/the_mult/m_mul_command[5] ,
         \UUT/Mpath/the_mult/x_mult_out[0] ,
         \UUT/Mpath/the_mult/x_mult_out[1] ,
         \UUT/Mpath/the_mult/x_mult_out[2] ,
         \UUT/Mpath/the_mult/x_mult_out[3] ,
         \UUT/Mpath/the_mult/x_mult_out[4] ,
         \UUT/Mpath/the_mult/x_mult_out[5] ,
         \UUT/Mpath/the_mult/x_mult_out[6] ,
         \UUT/Mpath/the_mult/x_mult_out[7] ,
         \UUT/Mpath/the_mult/x_mult_out[8] ,
         \UUT/Mpath/the_mult/x_mult_out[9] ,
         \UUT/Mpath/the_mult/x_mult_out[10] ,
         \UUT/Mpath/the_mult/x_mult_out[11] ,
         \UUT/Mpath/the_mult/x_mult_out[12] ,
         \UUT/Mpath/the_mult/x_mult_out[13] ,
         \UUT/Mpath/the_mult/x_mult_out[14] ,
         \UUT/Mpath/the_mult/x_mult_out[15] ,
         \UUT/Mpath/the_mult/x_mult_out[16] ,
         \UUT/Mpath/the_mult/x_mult_out[17] ,
         \UUT/Mpath/the_mult/x_mult_out[18] ,
         \UUT/Mpath/the_mult/x_mult_out[19] ,
         \UUT/Mpath/the_mult/x_mult_out[20] ,
         \UUT/Mpath/the_mult/x_mult_out[21] ,
         \UUT/Mpath/the_mult/x_mult_out[22] ,
         \UUT/Mpath/the_mult/x_mult_out[23] ,
         \UUT/Mpath/the_mult/x_mult_out[24] ,
         \UUT/Mpath/the_mult/x_mult_out[25] ,
         \UUT/Mpath/the_mult/x_mult_out[26] ,
         \UUT/Mpath/the_mult/x_mult_out[27] ,
         \UUT/Mpath/the_mult/x_mult_out[28] ,
         \UUT/Mpath/the_mult/x_mult_out[29] ,
         \UUT/Mpath/the_mult/x_mult_out[30] ,
         \UUT/Mpath/the_mult/x_mult_out[31] ,
         \UUT/Mpath/the_mult/x_mult_out[32] ,
         \UUT/Mpath/the_mult/x_mult_out[33] ,
         \UUT/Mpath/the_mult/x_mult_out[34] ,
         \UUT/Mpath/the_mult/x_mult_out[35] ,
         \UUT/Mpath/the_mult/x_mult_out[36] ,
         \UUT/Mpath/the_mult/x_mult_out[37] ,
         \UUT/Mpath/the_mult/x_mult_out[38] ,
         \UUT/Mpath/the_mult/x_mult_out[39] ,
         \UUT/Mpath/the_mult/x_mult_out[40] ,
         \UUT/Mpath/the_mult/x_mult_out[41] ,
         \UUT/Mpath/the_mult/x_mult_out[42] ,
         \UUT/Mpath/the_mult/x_mult_out[43] ,
         \UUT/Mpath/the_mult/x_mult_out[44] ,
         \UUT/Mpath/the_mult/x_mult_out[45] ,
         \UUT/Mpath/the_mult/x_mult_out[46] ,
         \UUT/Mpath/the_mult/x_mult_out[47] ,
         \UUT/Mpath/the_mult/x_mult_out[48] ,
         \UUT/Mpath/the_mult/x_mult_out[49] ,
         \UUT/Mpath/the_mult/x_mult_out[50] ,
         \UUT/Mpath/the_mult/x_mult_out[51] ,
         \UUT/Mpath/the_mult/x_mult_out[52] ,
         \UUT/Mpath/the_mult/x_mult_out[53] ,
         \UUT/Mpath/the_mult/x_mult_out[54] ,
         \UUT/Mpath/the_mult/x_mult_out[55] ,
         \UUT/Mpath/the_mult/x_mult_out[56] ,
         \UUT/Mpath/the_mult/x_mult_out[57] ,
         \UUT/Mpath/the_mult/x_mult_out[58] ,
         \UUT/Mpath/the_mult/x_mult_out[59] ,
         \UUT/Mpath/the_mult/x_mult_out[60] ,
         \UUT/Mpath/the_mult/x_mult_out[61] ,
         \UUT/Mpath/the_mult/x_mult_out[62] ,
         \UUT/Mpath/the_mult/x_mult_out[63] ,
         \UUT/Mpath/the_mult/x_mul_command[0] ,
         \UUT/Mpath/the_mult/x_mul_command[1] ,
         \UUT/Mpath/the_mult/x_mul_command[2] ,
         \UUT/Mpath/the_mult/x_mul_command[3] ,
         \UUT/Mpath/the_mult/x_mul_command[4] ,
         \UUT/Mpath/the_mult/x_mul_command[5] ,
         \UUT/Mpath/the_mult/x_operand1[0] ,
         \UUT/Mpath/the_mult/x_operand1[1] ,
         \UUT/Mpath/the_mult/x_operand1[2] ,
         \UUT/Mpath/the_mult/x_operand1[3] ,
         \UUT/Mpath/the_mult/x_operand1[4] ,
         \UUT/Mpath/the_mult/x_operand1[5] ,
         \UUT/Mpath/the_mult/x_operand1[6] ,
         \UUT/Mpath/the_mult/x_operand1[7] ,
         \UUT/Mpath/the_mult/x_operand1[8] ,
         \UUT/Mpath/the_mult/x_operand1[9] ,
         \UUT/Mpath/the_mult/x_operand1[10] ,
         \UUT/Mpath/the_mult/x_operand1[11] ,
         \UUT/Mpath/the_mult/x_operand1[12] ,
         \UUT/Mpath/the_mult/x_operand1[13] ,
         \UUT/Mpath/the_mult/x_operand1[14] ,
         \UUT/Mpath/the_mult/x_operand1[15] ,
         \UUT/Mpath/the_mult/x_operand1[16] ,
         \UUT/Mpath/the_mult/x_operand1[17] ,
         \UUT/Mpath/the_mult/x_operand1[18] ,
         \UUT/Mpath/the_mult/x_operand1[19] ,
         \UUT/Mpath/the_mult/x_operand1[20] ,
         \UUT/Mpath/the_mult/x_operand1[21] ,
         \UUT/Mpath/the_mult/x_operand1[22] ,
         \UUT/Mpath/the_mult/x_operand1[23] ,
         \UUT/Mpath/the_mult/x_operand1[24] ,
         \UUT/Mpath/the_mult/x_operand1[25] ,
         \UUT/Mpath/the_mult/x_operand1[26] ,
         \UUT/Mpath/the_mult/x_operand1[27] ,
         \UUT/Mpath/the_mult/x_operand1[28] ,
         \UUT/Mpath/the_mult/x_operand1[29] ,
         \UUT/Mpath/the_mult/x_operand1[30] ,
         \UUT/Mpath/the_mult/x_operand1[31] , \UUT/Mpath/the_memhandle/N244 ,
         \UUT/Mpath/the_memhandle/N243 , \UUT/Mpath/the_memhandle/N242 ,
         \UUT/Mpath/the_memhandle/N241 , \UUT/Mpath/the_memhandle/N240 ,
         \UUT/Mpath/the_memhandle/N239 , \UUT/Mpath/the_memhandle/N238 ,
         \UUT/Mpath/the_memhandle/N237 , \UUT/Mpath/the_memhandle/N236 ,
         \UUT/Mpath/the_memhandle/N235 , \UUT/Mpath/the_memhandle/N234 ,
         \UUT/Mpath/the_memhandle/N120 , \UUT/Mpath/the_memhandle/N86 ,
         \UUT/Mpath/the_memhandle/N77 , \UUT/Mpath/the_memhandle/N76 ,
         \UUT/Mpath/the_memhandle/N74 , \UUT/Mpath/the_memhandle/N72 ,
         \UUT/Mpath/the_memhandle/N39 , \UUT/Mpath/the_memhandle/N38 ,
         \UUT/Mpath/the_memhandle/N37 , \UUT/Mpath/the_memhandle/N36 ,
         \UUT/Mpath/the_memhandle/N34 , \UUT/Mpath/the_memhandle/smdr_out[16] ,
         \UUT/Mpath/the_memhandle/smdr_out[17] ,
         \UUT/Mpath/the_memhandle/smdr_out[18] ,
         \UUT/Mpath/the_memhandle/smdr_out[19] ,
         \UUT/Mpath/the_memhandle/smdr_out[20] ,
         \UUT/Mpath/the_memhandle/smdr_out[21] ,
         \UUT/Mpath/the_memhandle/smdr_out[22] ,
         \UUT/Mpath/the_memhandle/smdr_out[23] ,
         \UUT/Mpath/the_memhandle/smdr_out[24] ,
         \UUT/Mpath/the_memhandle/smdr_out[25] ,
         \UUT/Mpath/the_memhandle/smdr_out[26] ,
         \UUT/Mpath/the_memhandle/smdr_out[27] ,
         \UUT/Mpath/the_memhandle/smdr_out[28] ,
         \UUT/Mpath/the_memhandle/smdr_out[29] ,
         \UUT/Mpath/the_memhandle/smdr_out[30] ,
         \UUT/Mpath/the_memhandle/smdr_out[31] , n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n223, n224, n225, n227, n229,
         n230, n231, n232, n233, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n255, n256, n257, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2642, n2645, n2648, n2651, n2654, n2657,
         n2660, n2663, n2666, n2669, n2671, n2674, n2681, n2684, n2687, n2690,
         n2693, n2696, n2699, n2703, n2709, n2710, n2711, n2712, n2713, n2715,
         n2717, n2719, n2724, n2727, n2728, n2730, n2732, n2734, n2736, n2761,
         n2763, n2764, n2765, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5327, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5911, n5913, n5914, n5915, n5916, n5917, n5920, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5944, n5945, n5946, n5947, n5948, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6034, n6035, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6282, n6283, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, dram_mw, dram_mr,
         \dram_data_outbus[9] , \dram_data_outbus[8] , \dram_data_outbus[7] ,
         \dram_data_outbus[6] , \dram_data_outbus[5] , \dram_data_outbus[4] ,
         \dram_data_outbus[3] , \dram_data_outbus[31] , \dram_data_outbus[30] ,
         \dram_data_outbus[2] , \dram_data_outbus[29] , \dram_data_outbus[28] ,
         \dram_data_outbus[27] , \dram_data_outbus[26] ,
         \dram_data_outbus[25] , \dram_data_outbus[24] ,
         \dram_data_outbus[23] , \dram_data_outbus[22] ,
         \dram_data_outbus[21] , \dram_data_outbus[20] , \dram_data_outbus[1] ,
         \dram_data_outbus[19] , \dram_data_outbus[18] ,
         \dram_data_outbus[17] , \dram_data_outbus[16] ,
         \dram_data_outbus[15] , \dram_data_outbus[14] ,
         \dram_data_outbus[13] , \dram_data_outbus[12] ,
         \dram_data_outbus[11] , \dram_data_outbus[10] , \dram_data_outbus[0] ,
         \dram_data_inbus[9] , \dram_data_inbus[8] , \dram_data_inbus[7] ,
         \dram_data_inbus[6] , \dram_data_inbus[5] , \dram_data_inbus[4] ,
         \dram_data_inbus[3] , \dram_data_inbus[31] , \dram_data_inbus[30] ,
         \dram_data_inbus[2] , \dram_data_inbus[29] , \dram_data_inbus[28] ,
         \dram_data_inbus[27] , \dram_data_inbus[26] , \dram_data_inbus[25] ,
         \dram_data_inbus[24] , \dram_data_inbus[23] , \dram_data_inbus[22] ,
         \dram_data_inbus[21] , \dram_data_inbus[20] , \dram_data_inbus[1] ,
         \dram_data_inbus[19] , \dram_data_inbus[18] , \dram_data_inbus[17] ,
         \dram_data_inbus[16] , \dram_data_inbus[15] , \dram_data_inbus[14] ,
         \dram_data_inbus[13] , \dram_data_inbus[12] , \dram_data_inbus[11] ,
         \dram_data_inbus[10] , \dram_data_inbus[0] , \dram_addr_outbus[9] ,
         \dram_addr_outbus[8] , \dram_addr_outbus[7] , \dram_addr_outbus[6] ,
         \dram_addr_outbus[5] , \dram_addr_outbus[4] , \dram_addr_outbus[3] ,
         \dram_addr_outbus[2] , \dram_addr_outbus[12] , \dram_addr_outbus[11] ,
         \dram_addr_outbus[10] , n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432;
  wire   [31:0] I_DATA_INBUS;
  wire   [31:0] D_ADDR_OUTBUS;
  wire   [31:0] D_DATA_INBUS;
  wire   [31:0] D_DATA_OUTBUS;
  wire   [31:0] d_select;
  wire   [5:0] \UUT/d_mul_command ;
  wire   [2:0] \UUT/exe_outsel ;
  wire   [2:0] \UUT/shift_op ;
  wire   [23:0] \UUT/jar_in ;
  wire   [31:0] \UUT/branch_regb ;
  wire   [31:0] \UUT/branch_rega ;
  wire   [4:0] \UUT/rd_addr ;
  wire   [4:0] \UUT/rs2_addr ;
  wire   [4:0] \UUT/rs1_addr ;
  wire   [31:0] \UUT/daddr_out ;
  wire   [5:0] \UUT/Mcontrol/x_mul_command ;
  wire   [31:0] \UUT/Mcontrol/d_instr ;
  wire   [31:0] \UUT/Mcontrol/d_sampled_finstr ;
  wire   [23:0] \UUT/Mcontrol/f_currpc ;
  wire   [23:0] \UUT/Mcontrol/Nextpc_decoding/Bta ;
  wire   [1:0] \UUT/Mpath/mem_baddr ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_sll ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_srl ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_sra ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_ror ;
  wire   [31:0] \UUT/Mpath/the_shift/sh_rol ;
  wire   [63:0] \UUT/Mpath/the_mult/Mad_out ;
  wire   [31:0] \UUT/Mpath/the_mult/x_operand2 ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;
  assign \UUT/Mcontrol/int_reset  = reset;

  INV_X2 \UUT/Mpath/the_memhandle/I_0  ( .A(dmem_isbyte), .ZN(
        \UUT/Mpath/the_memhandle/N234 ) );
  INV_X2 \UUT/Mpath/the_memhandle/I_3  ( .A(dmem_ishalf), .ZN(
        \UUT/Mpath/the_memhandle/N237 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C342  ( .A1(\UUT/Mpath/the_memhandle/N235 ), 
        .A2(\UUT/Mpath/the_memhandle/N236 ), .ZN(\UUT/Mpath/the_memhandle/N34 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C344  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N36 ) );
  INV_X2 \UUT/Mpath/the_memhandle/I_8  ( .A(\UUT/Mpath/the_memhandle/N241 ), 
        .ZN(\UUT/Mpath/the_memhandle/N37 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C348  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N241 )
         );
  INV_X2 \UUT/Mpath/the_memhandle/I_9  ( .A(\UUT/Mpath/the_memhandle/N242 ), 
        .ZN(\UUT/Mpath/the_memhandle/N38 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C351  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N242 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C353  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N39 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C354  ( .A1(\UUT/m_mem_command[SIGN] ), 
        .A2(\UUT/Mpath/the_memhandle/N236 ), .ZN(\UUT/Mpath/the_memhandle/N72 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C356  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N74 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C360  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/the_memhandle/N240 ), .ZN(\UUT/Mpath/the_memhandle/N243 )
         );
  INV_X2 \UUT/Mpath/the_memhandle/I_12  ( .A(\UUT/Mpath/the_memhandle/N244 ), 
        .ZN(\UUT/Mpath/the_memhandle/N76 ) );
  OR2_X2 \UUT/Mpath/the_memhandle/C363  ( .A1(\UUT/Mpath/the_memhandle/N239 ), 
        .A2(\UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N244 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C365  ( .A1(\UUT/Mpath/mem_baddr [1]), .A2(
        \UUT/Mpath/mem_baddr [0]), .ZN(\UUT/Mpath/the_memhandle/N77 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C366  ( .A1(\UUT/Mpath/the_memhandle/N235 ), 
        .A2(\UUT/Mpath/the_memhandle/N238 ), .ZN(\UUT/Mpath/the_memhandle/N86 ) );
  AND2_X2 \UUT/Mpath/the_memhandle/C369  ( .A1(\UUT/m_mem_command[SIGN] ), 
        .A2(\UUT/Mpath/the_memhandle/N238 ), .ZN(
        \UUT/Mpath/the_memhandle/N120 ) );
  OR2_X2 \UUT/Mpath/the_mult/C331  ( .A1(\UUT/Mpath/the_mult/x_mul_command[4] ), .A2(\UUT/Mpath/the_mult/x_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N194 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C332  ( .A1(\UUT/Mpath/the_mult/N192 ), .A2(
        \UUT/Mpath/the_mult/N194 ), .ZN(\UUT/Mpath/the_mult/N195 ) );
  OR2_X2 \UUT/Mpath/the_mult/C333  ( .A1(\UUT/Mpath/the_mult/x_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N195 ), .ZN(\UUT/Mpath/the_mult/N196 ) );
  OR2_X2 \UUT/Mpath/the_mult/C334  ( .A1(\UUT/Mpath/the_mult/x_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N196 ), .ZN(\UUT/Mpath/the_mult/N197 ) );
  OR2_X2 \UUT/Mpath/the_mult/C335  ( .A1(\UUT/Mpath/the_mult/N193 ), .A2(
        \UUT/Mpath/the_mult/N197 ), .ZN(\UUT/Mpath/the_mult/N198 ) );
  OR2_X2 \UUT/Mpath/the_mult/C353  ( .A1(\UUT/Mpath/the_mult/x_mul_command[4] ), .A2(\UUT/Mpath/the_mult/x_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N212 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C354  ( .A1(\UUT/Mpath/the_mult/N192 ), .A2(
        \UUT/Mpath/the_mult/N212 ), .ZN(\UUT/Mpath/the_mult/N213 ) );
  OR2_X2 \UUT/Mpath/the_mult/C355  ( .A1(\UUT/Mpath/the_mult/x_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N213 ), .ZN(\UUT/Mpath/the_mult/N214 ) );
  OR2_X2 \UUT/Mpath/the_mult/C356  ( .A1(\UUT/Mpath/the_mult/x_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N214 ), .ZN(\UUT/Mpath/the_mult/N215 ) );
  OR2_X2 \UUT/Mpath/the_mult/C357  ( .A1(\UUT/Mpath/the_mult/x_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N215 ), .ZN(\UUT/Mpath/the_mult/N216 ) );
  INV_X2 \UUT/Mpath/the_mult/I_8  ( .A(\UUT/d_mul_command [3]), .ZN(
        \UUT/Mpath/the_mult/N220 ) );
  INV_X2 \UUT/Mpath/the_mult/I_9  ( .A(\UUT/d_mul_command [2]), .ZN(
        \UUT/Mpath/the_mult/N221 ) );
  INV_X2 \UUT/Mpath/the_mult/I_10  ( .A(\UUT/d_mul_command [1]), .ZN(
        \UUT/Mpath/the_mult/N222 ) );
  INV_X2 \UUT/Mpath/the_mult/I_11  ( .A(\UUT/d_mul_command [0]), .ZN(
        \UUT/Mpath/the_mult/N223 ) );
  OR2_X2 \UUT/Mpath/the_mult/C370  ( .A1(\UUT/d_mul_command [4]), .A2(
        \UUT/d_mul_command [5]), .ZN(\UUT/Mpath/the_mult/N224 ) );
  OR2_X2 \UUT/Mpath/the_mult/C371  ( .A1(\UUT/Mpath/the_mult/N220 ), .A2(
        \UUT/Mpath/the_mult/N224 ), .ZN(\UUT/Mpath/the_mult/N225 ) );
  OR2_X2 \UUT/Mpath/the_mult/C372  ( .A1(\UUT/Mpath/the_mult/N221 ), .A2(
        \UUT/Mpath/the_mult/N225 ), .ZN(\UUT/Mpath/the_mult/N226 ) );
  OR2_X2 \UUT/Mpath/the_mult/C373  ( .A1(\UUT/Mpath/the_mult/N222 ), .A2(
        \UUT/Mpath/the_mult/N226 ), .ZN(\UUT/Mpath/the_mult/N227 ) );
  OR2_X2 \UUT/Mpath/the_mult/C404  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N251 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C405  ( .A1(\UUT/Mpath/the_mult/N229 ), .A2(
        \UUT/Mpath/the_mult/N251 ), .ZN(\UUT/Mpath/the_mult/N252 ) );
  OR2_X2 \UUT/Mpath/the_mult/C406  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N252 ), .ZN(\UUT/Mpath/the_mult/N253 ) );
  OR2_X2 \UUT/Mpath/the_mult/C407  ( .A1(\UUT/Mpath/the_mult/N230 ), .A2(
        \UUT/Mpath/the_mult/N253 ), .ZN(\UUT/Mpath/the_mult/N254 ) );
  OR2_X2 \UUT/Mpath/the_mult/C410  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N257 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C411  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N257 ), .ZN(\UUT/Mpath/the_mult/N258 ) );
  OR2_X2 \UUT/Mpath/the_mult/C412  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N258 ), .ZN(\UUT/Mpath/the_mult/N259 ) );
  OR2_X2 \UUT/Mpath/the_mult/C413  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N259 ), .ZN(\UUT/Mpath/the_mult/N260 ) );
  OR2_X2 \UUT/Mpath/the_mult/C414  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N260 ), .ZN(\UUT/Mpath/the_mult/N261 ) );
  INV_X2 \UUT/Mpath/the_mult/I_21  ( .A(\UUT/Mpath/the_mult/N261 ), .ZN(
        \UUT/Mpath/the_mult/N262 ) );
  OR2_X2 \UUT/Mpath/the_mult/C417  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N263 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C418  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N263 ), .ZN(\UUT/Mpath/the_mult/N264 ) );
  OR2_X2 \UUT/Mpath/the_mult/C419  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N264 ), .ZN(\UUT/Mpath/the_mult/N265 ) );
  OR2_X2 \UUT/Mpath/the_mult/C420  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N265 ), .ZN(\UUT/Mpath/the_mult/N266 ) );
  OR2_X2 \UUT/Mpath/the_mult/C421  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N266 ), .ZN(\UUT/Mpath/the_mult/N267 ) );
  INV_X2 \UUT/Mpath/the_mult/I_22  ( .A(\UUT/Mpath/the_mult/N267 ), .ZN(
        \UUT/Mpath/the_mult/N268 ) );
  OR2_X2 \UUT/Mpath/the_mult/C424  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N269 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C425  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N269 ), .ZN(\UUT/Mpath/the_mult/N270 ) );
  OR2_X2 \UUT/Mpath/the_mult/C426  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N270 ), .ZN(\UUT/Mpath/the_mult/N271 ) );
  OR2_X2 \UUT/Mpath/the_mult/C427  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N271 ), .ZN(\UUT/Mpath/the_mult/N272 ) );
  OR2_X2 \UUT/Mpath/the_mult/C428  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N272 ), .ZN(\UUT/Mpath/the_mult/N273 ) );
  INV_X2 \UUT/Mpath/the_mult/I_23  ( .A(\UUT/Mpath/the_mult/N273 ), .ZN(
        \UUT/Mpath/the_mult/N274 ) );
  OR2_X2 \UUT/Mpath/the_mult/C432  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N275 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C433  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N275 ), .ZN(\UUT/Mpath/the_mult/N276 ) );
  OR2_X2 \UUT/Mpath/the_mult/C434  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N276 ), .ZN(\UUT/Mpath/the_mult/N277 ) );
  OR2_X2 \UUT/Mpath/the_mult/C435  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N277 ), .ZN(\UUT/Mpath/the_mult/N278 ) );
  OR2_X2 \UUT/Mpath/the_mult/C436  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N278 ), .ZN(\UUT/Mpath/the_mult/N279 ) );
  INV_X2 \UUT/Mpath/the_mult/I_24  ( .A(\UUT/Mpath/the_mult/N279 ), .ZN(
        \UUT/Mpath/the_mult/N280 ) );
  OR2_X2 \UUT/Mpath/the_mult/C440  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N281 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C441  ( .A1(\UUT/Mpath/the_mult/N229 ), .A2(
        \UUT/Mpath/the_mult/N281 ), .ZN(\UUT/Mpath/the_mult/N282 ) );
  OR2_X2 \UUT/Mpath/the_mult/C442  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N282 ), .ZN(\UUT/Mpath/the_mult/N283 ) );
  OR2_X2 \UUT/Mpath/the_mult/C443  ( .A1(\UUT/Mpath/the_mult/N230 ), .A2(
        \UUT/Mpath/the_mult/N283 ), .ZN(\UUT/Mpath/the_mult/N284 ) );
  OR2_X2 \UUT/Mpath/the_mult/C446  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N287 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C447  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N287 ), .ZN(\UUT/Mpath/the_mult/N288 ) );
  OR2_X2 \UUT/Mpath/the_mult/C448  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N288 ), .ZN(\UUT/Mpath/the_mult/N289 ) );
  OR2_X2 \UUT/Mpath/the_mult/C449  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N289 ), .ZN(\UUT/Mpath/the_mult/N290 ) );
  OR2_X2 \UUT/Mpath/the_mult/C450  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N290 ), .ZN(\UUT/Mpath/the_mult/N291 ) );
  INV_X2 \UUT/Mpath/the_mult/I_26  ( .A(\UUT/Mpath/the_mult/N291 ), .ZN(
        \UUT/Mpath/the_mult/N292 ) );
  OR2_X2 \UUT/Mpath/the_mult/C453  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N293 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C454  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N293 ), .ZN(\UUT/Mpath/the_mult/N294 ) );
  OR2_X2 \UUT/Mpath/the_mult/C455  ( .A1(\UUT/Mpath/the_mult/m_mul_command[2] ), .A2(\UUT/Mpath/the_mult/N294 ), .ZN(\UUT/Mpath/the_mult/N295 ) );
  OR2_X2 \UUT/Mpath/the_mult/C456  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N295 ), .ZN(\UUT/Mpath/the_mult/N296 ) );
  OR2_X2 \UUT/Mpath/the_mult/C457  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N296 ), .ZN(\UUT/Mpath/the_mult/N297 ) );
  INV_X2 \UUT/Mpath/the_mult/I_27  ( .A(\UUT/Mpath/the_mult/N297 ), .ZN(
        \UUT/Mpath/the_mult/N298 ) );
  OR2_X2 \UUT/Mpath/the_mult/C460  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N299 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C461  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N299 ), .ZN(\UUT/Mpath/the_mult/N300 ) );
  OR2_X2 \UUT/Mpath/the_mult/C462  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N300 ), .ZN(\UUT/Mpath/the_mult/N301 ) );
  OR2_X2 \UUT/Mpath/the_mult/C463  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N301 ), .ZN(\UUT/Mpath/the_mult/N302 ) );
  OR2_X2 \UUT/Mpath/the_mult/C464  ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(\UUT/Mpath/the_mult/N302 ), .ZN(\UUT/Mpath/the_mult/N303 ) );
  INV_X2 \UUT/Mpath/the_mult/I_28  ( .A(\UUT/Mpath/the_mult/N303 ), .ZN(
        \UUT/Mpath/the_mult/N304 ) );
  OR2_X2 \UUT/Mpath/the_mult/C468  ( .A1(\UUT/Mpath/the_mult/m_mul_command[4] ), .A2(\UUT/Mpath/the_mult/m_mul_command[5] ), .ZN(\UUT/Mpath/the_mult/N305 )
         );
  OR2_X2 \UUT/Mpath/the_mult/C469  ( .A1(\UUT/Mpath/the_mult/m_mul_command[3] ), .A2(\UUT/Mpath/the_mult/N305 ), .ZN(\UUT/Mpath/the_mult/N306 ) );
  OR2_X2 \UUT/Mpath/the_mult/C470  ( .A1(\UUT/Mpath/the_mult/N244 ), .A2(
        \UUT/Mpath/the_mult/N306 ), .ZN(\UUT/Mpath/the_mult/N307 ) );
  OR2_X2 \UUT/Mpath/the_mult/C471  ( .A1(\UUT/Mpath/the_mult/m_mul_command[1] ), .A2(\UUT/Mpath/the_mult/N307 ), .ZN(\UUT/Mpath/the_mult/N308 ) );
  OR2_X2 \UUT/Mpath/the_mult/C472  ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(
        \UUT/Mpath/the_mult/N308 ), .ZN(\UUT/Mpath/the_mult/N309 ) );
  INV_X2 \UUT/Mpath/the_mult/I_29  ( .A(\UUT/Mpath/the_mult/N309 ), .ZN(
        \UUT/Mpath/the_mult/N310 ) );
  OR2_X2 \UUT/Mpath/the_mult/C499  ( .A1(\UUT/Mpath/the_mult/N274 ), .A2(
        \UUT/Mpath/the_mult/N280 ), .ZN(\UUT/Mpath/the_mult/N312 ) );
  OR2_X2 \UUT/Mpath/the_mult/C507  ( .A1(\UUT/Mpath/the_mult/N304 ), .A2(
        \UUT/Mpath/the_mult/N310 ), .ZN(\UUT/Mpath/the_mult/N314 ) );
  OR2_X2 \UUT/Mpath/the_shift/C151  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/Mpath/the_shift/N104 ), .ZN(\UUT/Mpath/the_shift/N106 ) );
  OR2_X2 \UUT/Mpath/the_shift/C152  ( .A1(\UUT/Mpath/the_shift/N105 ), .A2(
        \UUT/Mpath/the_shift/N106 ), .ZN(\UUT/Mpath/the_shift/N107 ) );
  OR2_X2 \UUT/Mpath/the_shift/C155  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/Mpath/the_shift/N104 ), .ZN(\UUT/Mpath/the_shift/N109 ) );
  OR2_X2 \UUT/Mpath/the_shift/C156  ( .A1(\UUT/shift_op [0]), .A2(
        \UUT/Mpath/the_shift/N109 ), .ZN(\UUT/Mpath/the_shift/N110 ) );
  INV_X2 \UUT/Mpath/the_shift/I_3  ( .A(\UUT/Mpath/the_shift/N110 ), .ZN(
        \UUT/Mpath/the_shift/N111 ) );
  OR2_X2 \UUT/Mpath/the_shift/C159  ( .A1(\UUT/Mpath/the_shift/N112 ), .A2(
        \UUT/shift_op [2]), .ZN(\UUT/Mpath/the_shift/N113 ) );
  OR2_X2 \UUT/Mpath/the_shift/C160  ( .A1(\UUT/shift_op [0]), .A2(
        \UUT/Mpath/the_shift/N113 ), .ZN(\UUT/Mpath/the_shift/N114 ) );
  INV_X2 \UUT/Mpath/the_shift/I_5  ( .A(\UUT/Mpath/the_shift/N114 ), .ZN(
        \UUT/Mpath/the_shift/N115 ) );
  OR2_X2 \UUT/Mpath/the_shift/C163  ( .A1(\UUT/shift_op [1]), .A2(
        \UUT/shift_op [2]), .ZN(\UUT/Mpath/the_shift/N116 ) );
  OR2_X2 \UUT/Mpath/the_shift/C164  ( .A1(\UUT/Mpath/the_shift/N105 ), .A2(
        \UUT/Mpath/the_shift/N116 ), .ZN(\UUT/Mpath/the_shift/N117 ) );
  OR2_X2 \UUT/Mpath/the_alu/C476  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N469 ) );
  OR2_X2 \UUT/Mpath/the_alu/C477  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N469 ), .ZN(\UUT/Mpath/the_alu/N470 ) );
  OR2_X2 \UUT/Mpath/the_alu/C478  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N470 ), .ZN(\UUT/Mpath/the_alu/N471 ) );
  OR2_X2 \UUT/Mpath/the_alu/C479  ( .A1(\UUT/Mpath/the_alu/N467 ), .A2(
        \UUT/Mpath/the_alu/N471 ), .ZN(\UUT/Mpath/the_alu/N472 ) );
  OR2_X2 \UUT/Mpath/the_alu/C480  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N472 ), .ZN(\UUT/Mpath/the_alu/N473 ) );
  INV_X2 \UUT/Mpath/the_alu/I_9  ( .A(\UUT/Mpath/the_alu/N473 ), .ZN(
        \UUT/Mpath/the_alu/N474 ) );
  OR2_X2 \UUT/Mpath/the_alu/C485  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N475 ) );
  OR2_X2 \UUT/Mpath/the_alu/C486  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N475 ), .ZN(\UUT/Mpath/the_alu/N476 ) );
  OR2_X2 \UUT/Mpath/the_alu/C487  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N476 ), .ZN(\UUT/Mpath/the_alu/N477 ) );
  OR2_X2 \UUT/Mpath/the_alu/C488  ( .A1(\UUT/Mpath/the_alu/N467 ), .A2(
        \UUT/Mpath/the_alu/N477 ), .ZN(\UUT/Mpath/the_alu/N478 ) );
  OR2_X2 \UUT/Mpath/the_alu/C489  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N478 ), .ZN(\UUT/Mpath/the_alu/N479 ) );
  INV_X2 \UUT/Mpath/the_alu/I_10  ( .A(\UUT/Mpath/the_alu/N479 ), .ZN(
        \UUT/Mpath/the_alu/N480 ) );
  OR2_X2 \UUT/Mpath/the_alu/C494  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N481 ) );
  OR2_X2 \UUT/Mpath/the_alu/C495  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N481 ), .ZN(\UUT/Mpath/the_alu/N482 ) );
  OR2_X2 \UUT/Mpath/the_alu/C496  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N482 ), .ZN(\UUT/Mpath/the_alu/N483 ) );
  OR2_X2 \UUT/Mpath/the_alu/C497  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N483 ), .ZN(\UUT/Mpath/the_alu/N484 ) );
  OR2_X2 \UUT/Mpath/the_alu/C498  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N484 ), .ZN(\UUT/Mpath/the_alu/N485 ) );
  INV_X2 \UUT/Mpath/the_alu/I_11  ( .A(\UUT/Mpath/the_alu/N485 ), .ZN(
        \UUT/Mpath/the_alu/N486 ) );
  OR2_X2 \UUT/Mpath/the_alu/C502  ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N487 ) );
  OR2_X2 \UUT/Mpath/the_alu/C503  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N487 ), .ZN(\UUT/Mpath/the_alu/N488 ) );
  OR2_X2 \UUT/Mpath/the_alu/C504  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N488 ), .ZN(\UUT/Mpath/the_alu/N489 ) );
  OR2_X2 \UUT/Mpath/the_alu/C505  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N489 ), .ZN(\UUT/Mpath/the_alu/N490 ) );
  OR2_X2 \UUT/Mpath/the_alu/C506  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N490 ), .ZN(\UUT/Mpath/the_alu/N491 ) );
  OR2_X2 \UUT/Mpath/the_alu/C510  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N493 ) );
  OR2_X2 \UUT/Mpath/the_alu/C511  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N493 ), .ZN(\UUT/Mpath/the_alu/N494 ) );
  OR2_X2 \UUT/Mpath/the_alu/C512  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N494 ), .ZN(\UUT/Mpath/the_alu/N495 ) );
  OR2_X2 \UUT/Mpath/the_alu/C513  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N495 ), .ZN(\UUT/Mpath/the_alu/N496 ) );
  OR2_X2 \UUT/Mpath/the_alu/C514  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N496 ), .ZN(\UUT/Mpath/the_alu/N497 ) );
  INV_X2 \UUT/Mpath/the_alu/I_13  ( .A(\UUT/Mpath/the_alu/N497 ), .ZN(
        \UUT/Mpath/the_alu/N498 ) );
  OR2_X2 \UUT/Mpath/the_alu/C517  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Mpath/the_alu/N466 ), .ZN(\UUT/Mpath/the_alu/N499 ) );
  OR2_X2 \UUT/Mpath/the_alu/C518  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N499 ), .ZN(\UUT/Mpath/the_alu/N500 ) );
  OR2_X2 \UUT/Mpath/the_alu/C519  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N500 ), .ZN(\UUT/Mpath/the_alu/N501 ) );
  OR2_X2 \UUT/Mpath/the_alu/C520  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N501 ), .ZN(\UUT/Mpath/the_alu/N502 ) );
  OR2_X2 \UUT/Mpath/the_alu/C521  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N502 ), .ZN(\UUT/Mpath/the_alu/N503 ) );
  OR2_X2 \UUT/Mpath/the_alu/C525  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N505 ), .ZN(\UUT/Mpath/the_alu/N506 ) );
  OR2_X2 \UUT/Mpath/the_alu/C526  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N506 ), .ZN(\UUT/Mpath/the_alu/N507 ) );
  OR2_X2 \UUT/Mpath/the_alu/C527  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N507 ), .ZN(\UUT/Mpath/the_alu/N508 ) );
  OR2_X2 \UUT/Mpath/the_alu/C528  ( .A1(\UUT/Alu_command[OP][0] ), .A2(
        \UUT/Mpath/the_alu/N508 ), .ZN(\UUT/Mpath/the_alu/N509 ) );
  OR2_X2 \UUT/Mpath/the_alu/C533  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N511 ), .ZN(\UUT/Mpath/the_alu/N512 ) );
  OR2_X2 \UUT/Mpath/the_alu/C534  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N512 ), .ZN(\UUT/Mpath/the_alu/N513 ) );
  OR2_X2 \UUT/Mpath/the_alu/C535  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N513 ), .ZN(\UUT/Mpath/the_alu/N514 ) );
  OR2_X2 \UUT/Mpath/the_alu/C536  ( .A1(\UUT/Mpath/the_alu/N468 ), .A2(
        \UUT/Mpath/the_alu/N514 ), .ZN(\UUT/Mpath/the_alu/N515 ) );
  OR2_X2 \UUT/Mpath/the_alu/C539  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N517 ), .ZN(\UUT/Mpath/the_alu/N518 ) );
  OR2_X2 \UUT/Mpath/the_alu/C540  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N518 ), .ZN(\UUT/Mpath/the_alu/N519 ) );
  OR2_X2 \UUT/Mpath/the_alu/C541  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N519 ), .ZN(\UUT/Mpath/the_alu/N520 ) );
  OR2_X2 \UUT/Mpath/the_alu/C545  ( .A1(\UUT/Alu_command[OP][4] ), .A2(
        \UUT/Alu_command[OP][5] ), .ZN(\UUT/Mpath/the_alu/N523 ) );
  OR2_X2 \UUT/Mpath/the_alu/C546  ( .A1(\UUT/Alu_command[OP][3] ), .A2(
        \UUT/Mpath/the_alu/N523 ), .ZN(\UUT/Mpath/the_alu/N524 ) );
  OR2_X2 \UUT/Mpath/the_alu/C547  ( .A1(\UUT/Alu_command[OP][2] ), .A2(
        \UUT/Mpath/the_alu/N524 ), .ZN(\UUT/Mpath/the_alu/N525 ) );
  OR2_X2 \UUT/Mpath/the_alu/C548  ( .A1(\UUT/Alu_command[OP][1] ), .A2(
        \UUT/Mpath/the_alu/N525 ), .ZN(\UUT/Mpath/the_alu/N526 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C649  ( .A(\UUT/Mpath/out_regA[23] ), .B(
        \UUT/Mpath/out_regB[23] ), .Z(\UUT/Mpath/the_alu/N166 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C650  ( .A(\UUT/Mpath/out_regA[22] ), .B(
        \UUT/Mpath/out_regB[22] ), .Z(\UUT/Mpath/the_alu/N167 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C651  ( .A(\UUT/Mpath/out_regA[21] ), .B(
        \UUT/Mpath/out_regB[21] ), .Z(\UUT/Mpath/the_alu/N168 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C652  ( .A(n7138), .B(n7194), .Z(
        \UUT/Mpath/the_alu/N169 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C653  ( .A(n7167), .B(n7190), .Z(
        \UUT/Mpath/the_alu/N170 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C654  ( .A(\UUT/Mpath/out_regA[18] ), .B(n7135), 
        .Z(\UUT/Mpath/the_alu/N171 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C655  ( .A(\UUT/Mpath/out_regA[17] ), .B(n7197), 
        .Z(\UUT/Mpath/the_alu/N172 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C656  ( .A(n7129), .B(n7136), .Z(
        \UUT/Mpath/the_alu/N173 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C657  ( .A(n7112), .B(n7125), .Z(
        \UUT/Mpath/the_alu/N174 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C658  ( .A(n7113), .B(n7140), .Z(
        \UUT/Mpath/the_alu/N175 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C659  ( .A(n1245), .B(n7122), .Z(
        \UUT/Mpath/the_alu/N176 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C660  ( .A(n7193), .B(n7134), .Z(
        \UUT/Mpath/the_alu/N177 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C661  ( .A(n7198), .B(n7107), .Z(
        \UUT/Mpath/the_alu/N178 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C662  ( .A(\UUT/Mpath/out_regA[10] ), .B(n7137), 
        .Z(\UUT/Mpath/the_alu/N179 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C663  ( .A(n7132), .B(n7128), .Z(
        \UUT/Mpath/the_alu/N180 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C664  ( .A(n7189), .B(\UUT/Mpath/out_regB[8] ), 
        .Z(\UUT/Mpath/the_alu/N181 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C665  ( .A(\UUT/Mpath/out_regA[7] ), .B(
        \UUT/Mpath/out_regB[7] ), .Z(\UUT/Mpath/the_alu/N182 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C666  ( .A(n7106), .B(n7099), .Z(
        \UUT/Mpath/the_alu/N183 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C667  ( .A(n1321), .B(n7114), .Z(
        \UUT/Mpath/the_alu/N184 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C668  ( .A(\UUT/Mpath/out_regA[4] ), .B(n7400), 
        .Z(\UUT/Mpath/the_alu/N185 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C669  ( .A(\UUT/Mpath/out_regA[3] ), .B(n7401), 
        .Z(\UUT/Mpath/the_alu/N186 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C670  ( .A(\UUT/Mpath/out_regA[2] ), .B(n7404), 
        .Z(\UUT/Mpath/the_alu/N187 ) );
  XOR2_X1 \UUT/Mpath/the_alu/C672  ( .A(\UUT/Mpath/out_regA[0] ), .B(n7408), 
        .Z(\UUT/Mpath/the_alu/N189 ) );
  AND2_X2 \UUT/Mpath/the_alu/C682  ( .A1(\UUT/Mpath/the_alu/N37 ), .A2(
        \UUT/Mpath/the_alu/N38 ), .ZN(\UUT/Mpath/the_alu/N198 ) );
  AND2_X2 \UUT/Mpath/the_alu/C683  ( .A1(\UUT/Mpath/the_alu/N39 ), .A2(
        \UUT/Mpath/the_alu/N40 ), .ZN(\UUT/Mpath/the_alu/N199 ) );
  AND2_X2 \UUT/Mpath/the_alu/C684  ( .A1(\UUT/Mpath/the_alu/N41 ), .A2(
        \UUT/Mpath/the_alu/N42 ), .ZN(\UUT/Mpath/the_alu/N200 ) );
  AND2_X2 \UUT/Mpath/the_alu/C685  ( .A1(\UUT/Mpath/the_alu/N43 ), .A2(
        \UUT/Mpath/the_alu/N44 ), .ZN(\UUT/Mpath/the_alu/N201 ) );
  AND2_X2 \UUT/Mpath/the_alu/C686  ( .A1(\UUT/Mpath/the_alu/N45 ), .A2(
        \UUT/Mpath/the_alu/N46 ), .ZN(\UUT/Mpath/the_alu/N202 ) );
  AND2_X2 \UUT/Mpath/the_alu/C687  ( .A1(\UUT/Mpath/the_alu/N47 ), .A2(
        \UUT/Mpath/the_alu/N48 ), .ZN(\UUT/Mpath/the_alu/N203 ) );
  AND2_X2 \UUT/Mpath/the_alu/C688  ( .A1(\UUT/Mpath/the_alu/N49 ), .A2(
        \UUT/Mpath/the_alu/N50 ), .ZN(\UUT/Mpath/the_alu/N204 ) );
  AND2_X2 \UUT/Mpath/the_alu/C689  ( .A1(\UUT/Mpath/the_alu/N51 ), .A2(
        \UUT/Mpath/the_alu/N52 ), .ZN(\UUT/Mpath/the_alu/N205 ) );
  AND2_X2 \UUT/Mpath/the_alu/C690  ( .A1(\UUT/Mpath/the_alu/N53 ), .A2(
        \UUT/Mpath/the_alu/N54 ), .ZN(\UUT/Mpath/the_alu/N206 ) );
  AND2_X2 \UUT/Mpath/the_alu/C691  ( .A1(\UUT/Mpath/the_alu/N55 ), .A2(
        \UUT/Mpath/the_alu/N56 ), .ZN(\UUT/Mpath/the_alu/N207 ) );
  AND2_X2 \UUT/Mpath/the_alu/C692  ( .A1(\UUT/Mpath/the_alu/N57 ), .A2(
        \UUT/Mpath/the_alu/N58 ), .ZN(\UUT/Mpath/the_alu/N208 ) );
  AND2_X2 \UUT/Mpath/the_alu/C693  ( .A1(\UUT/Mpath/the_alu/N59 ), .A2(
        \UUT/Mpath/the_alu/N60 ), .ZN(\UUT/Mpath/the_alu/N209 ) );
  AND2_X2 \UUT/Mpath/the_alu/C694  ( .A1(\UUT/Mpath/the_alu/N61 ), .A2(
        \UUT/Mpath/the_alu/N62 ), .ZN(\UUT/Mpath/the_alu/N210 ) );
  AND2_X2 \UUT/Mpath/the_alu/C695  ( .A1(\UUT/Mpath/the_alu/N63 ), .A2(
        \UUT/Mpath/the_alu/N64 ), .ZN(\UUT/Mpath/the_alu/N211 ) );
  AND2_X2 \UUT/Mpath/the_alu/C696  ( .A1(\UUT/Mpath/the_alu/N65 ), .A2(
        \UUT/Mpath/the_alu/N66 ), .ZN(\UUT/Mpath/the_alu/N212 ) );
  AND2_X2 \UUT/Mpath/the_alu/C697  ( .A1(\UUT/Mpath/the_alu/N67 ), .A2(
        \UUT/Mpath/the_alu/N68 ), .ZN(\UUT/Mpath/the_alu/N213 ) );
  AND2_X2 \UUT/Mpath/the_alu/C698  ( .A1(\UUT/Mpath/the_alu/N69 ), .A2(
        \UUT/Mpath/the_alu/N70 ), .ZN(\UUT/Mpath/the_alu/N214 ) );
  AND2_X2 \UUT/Mpath/the_alu/C699  ( .A1(\UUT/Mpath/the_alu/N71 ), .A2(
        \UUT/Mpath/the_alu/N72 ), .ZN(\UUT/Mpath/the_alu/N215 ) );
  AND2_X2 \UUT/Mpath/the_alu/C700  ( .A1(\UUT/Mpath/the_alu/N73 ), .A2(
        \UUT/Mpath/the_alu/N74 ), .ZN(\UUT/Mpath/the_alu/N216 ) );
  AND2_X2 \UUT/Mpath/the_alu/C701  ( .A1(\UUT/Mpath/the_alu/N75 ), .A2(
        \UUT/Mpath/the_alu/N76 ), .ZN(\UUT/Mpath/the_alu/N217 ) );
  AND2_X2 \UUT/Mpath/the_alu/C702  ( .A1(\UUT/Mpath/the_alu/N77 ), .A2(
        \UUT/Mpath/the_alu/N78 ), .ZN(\UUT/Mpath/the_alu/N218 ) );
  AND2_X2 \UUT/Mpath/the_alu/C703  ( .A1(\UUT/Mpath/the_alu/N79 ), .A2(
        \UUT/Mpath/the_alu/N80 ), .ZN(\UUT/Mpath/the_alu/N219 ) );
  AND2_X2 \UUT/Mpath/the_alu/C705  ( .A1(\UUT/Mpath/the_alu/N83 ), .A2(
        \UUT/Mpath/the_alu/N84 ), .ZN(\UUT/Mpath/the_alu/N221 ) );
  OR2_X2 \UUT/Mpath/C262  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/Mpath/N111 ), 
        .ZN(\UUT/Mpath/N113 ) );
  OR2_X2 \UUT/Mpath/C263  ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N113 ), .ZN(
        \UUT/Mpath/N114 ) );
  INV_X2 \UUT/Mpath/I_3  ( .A(\UUT/Mpath/N114 ), .ZN(\UUT/Mpath/N115 ) );
  OR2_X2 \UUT/Mpath/C266  ( .A1(\UUT/Mpath/N116 ), .A2(\UUT/exe_outsel [2]), 
        .ZN(\UUT/Mpath/N117 ) );
  OR2_X2 \UUT/Mpath/C267  ( .A1(\UUT/exe_outsel [0]), .A2(\UUT/Mpath/N117 ), 
        .ZN(\UUT/Mpath/N118 ) );
  INV_X2 \UUT/Mpath/I_5  ( .A(\UUT/Mpath/N118 ), .ZN(\UUT/Mpath/N119 ) );
  OR2_X2 \UUT/Mpath/C271  ( .A1(\UUT/Mpath/N116 ), .A2(\UUT/exe_outsel [2]), 
        .ZN(\UUT/Mpath/N121 ) );
  OR2_X2 \UUT/Mpath/C275  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/exe_outsel [2]), 
        .ZN(\UUT/Mpath/N124 ) );
  OR2_X2 \UUT/Mpath/C276  ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N124 ), .ZN(
        \UUT/Mpath/N125 ) );
  OR2_X2 \UUT/Mpath/C280  ( .A1(\UUT/exe_outsel [1]), .A2(\UUT/Mpath/N111 ), 
        .ZN(\UUT/Mpath/N127 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_0  ( .A(\UUT/Mcontrol/st_logic/load_stall ), 
        .ZN(\UUT/Mcontrol/st_logic/N12 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_3  ( .A(dmem_read), .ZN(
        \UUT/Mcontrol/st_logic/N15 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_4  ( .A(\UUT/byp_controlA[2] ), .ZN(
        \UUT/Mcontrol/st_logic/N55 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C75  ( .A1(\UUT/byp_controlA[0] ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N18 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_5  ( .A(\UUT/Mcontrol/st_logic/N18 ), .ZN(
        \UUT/Mcontrol/st_logic/N19 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_6  ( .A(\UUT/byp_controlB[2] ), .ZN(
        \UUT/Mcontrol/st_logic/N52 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C79  ( .A1(\UUT/byp_controlB[0] ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N22 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_7  ( .A(\UUT/Mcontrol/st_logic/N22 ), .ZN(
        \UUT/Mcontrol/st_logic/N23 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_8  ( .A(\UUT/m_mem_command[MR] ), .ZN(
        \UUT/Mcontrol/st_logic/N24 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C85  ( .A1(\UUT/Mcontrol/x_mul_command [4]), 
        .A2(\UUT/Mcontrol/x_mul_command [5]), .ZN(\UUT/Mcontrol/st_logic/N28 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C86  ( .A1(\UUT/Mcontrol/x_mul_command [3]), 
        .A2(\UUT/Mcontrol/st_logic/N28 ), .ZN(\UUT/Mcontrol/st_logic/N29 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C87  ( .A1(\UUT/Mcontrol/st_logic/N26 ), .A2(
        \UUT/Mcontrol/st_logic/N29 ), .ZN(\UUT/Mcontrol/st_logic/N30 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C88  ( .A1(\UUT/Mcontrol/st_logic/N27 ), .A2(
        \UUT/Mcontrol/st_logic/N30 ), .ZN(\UUT/Mcontrol/st_logic/N31 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C89  ( .A1(\UUT/Mcontrol/x_mul_command [0]), 
        .A2(\UUT/Mcontrol/st_logic/N31 ), .ZN(\UUT/Mcontrol/st_logic/N32 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_12  ( .A(\UUT/Mcontrol/st_logic/N32 ), .ZN(
        \UUT/Mcontrol/st_logic/N33 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C94  ( .A1(\UUT/Mcontrol/x_mul_command [4]), 
        .A2(\UUT/Mcontrol/x_mul_command [5]), .ZN(\UUT/Mcontrol/st_logic/N35 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C95  ( .A1(\UUT/Mcontrol/x_mul_command [3]), 
        .A2(\UUT/Mcontrol/st_logic/N35 ), .ZN(\UUT/Mcontrol/st_logic/N36 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C96  ( .A1(\UUT/Mcontrol/st_logic/N26 ), .A2(
        \UUT/Mcontrol/st_logic/N36 ), .ZN(\UUT/Mcontrol/st_logic/N37 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C97  ( .A1(\UUT/Mcontrol/st_logic/N27 ), .A2(
        \UUT/Mcontrol/st_logic/N37 ), .ZN(\UUT/Mcontrol/st_logic/N38 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C98  ( .A1(\UUT/Mcontrol/st_logic/N34 ), .A2(
        \UUT/Mcontrol/st_logic/N38 ), .ZN(\UUT/Mcontrol/st_logic/N39 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_14  ( .A(\UUT/Mcontrol/st_logic/N39 ), .ZN(
        \UUT/Mcontrol/st_logic/N40 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C104  ( .A1(\UUT/Mcontrol/st_logic/N42 ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N44 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_17  ( .A(\UUT/Mcontrol/st_logic/N44 ), .ZN(
        \UUT/Mcontrol/st_logic/N45 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_18  ( .A(
        \UUT/Mcontrol/st_logic/branch_uses_regb ), .ZN(
        \UUT/Mcontrol/st_logic/N46 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C110  ( .A1(\UUT/Mcontrol/st_logic/N47 ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N49 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_20  ( .A(\UUT/Mcontrol/st_logic/N49 ), .ZN(
        \UUT/Mcontrol/st_logic/N50 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_21  ( .A(n6877), .ZN(
        \UUT/Mcontrol/st_logic/N51 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C115  ( .A1(\UUT/byp_controlB[0] ), .A2(
        \UUT/Mcontrol/st_logic/N52 ), .ZN(\UUT/Mcontrol/st_logic/N53 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_22  ( .A(\UUT/Mcontrol/st_logic/N53 ), .ZN(
        \UUT/Mcontrol/st_logic/N54 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C120  ( .A1(\UUT/byp_controlA[0] ), .A2(
        \UUT/Mcontrol/st_logic/N55 ), .ZN(\UUT/Mcontrol/st_logic/N56 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_23  ( .A(\UUT/Mcontrol/st_logic/N56 ), .ZN(
        \UUT/Mcontrol/st_logic/N57 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_24  ( .A(\UUT/Mcontrol/d_jump_type[2] ), 
        .ZN(\UUT/Mcontrol/st_logic/N58 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C126  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N60 ), .ZN(\UUT/Mcontrol/st_logic/N61 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C128  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N62 ), .ZN(\UUT/Mcontrol/st_logic/N63 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_25  ( .A(\UUT/Mcontrol/st_logic/N63 ), .ZN(
        \UUT/Mcontrol/st_logic/N64 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_26  ( .A(\UUT/Mcontrol/d_jump_type[0] ), 
        .ZN(\UUT/Mcontrol/st_logic/N65 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C134  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N67 ), .ZN(\UUT/Mcontrol/st_logic/N68 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C136  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N69 ), .ZN(\UUT/Mcontrol/st_logic/N70 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_27  ( .A(\UUT/Mcontrol/st_logic/N70 ), .ZN(
        \UUT/Mcontrol/st_logic/N71 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C141  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N73 ), .ZN(\UUT/Mcontrol/st_logic/N74 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C155  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N85 ), .ZN(\UUT/Mcontrol/st_logic/N86 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C157  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N87 ), .ZN(\UUT/Mcontrol/st_logic/N88 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_30  ( .A(\UUT/Mcontrol/st_logic/N88 ), .ZN(
        \UUT/Mcontrol/st_logic/N89 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C163  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N92 ), .ZN(\UUT/Mcontrol/st_logic/N93 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C164  ( .A1(\UUT/Mcontrol/st_logic/N90 ), .A2(
        \UUT/Mcontrol/st_logic/N93 ), .ZN(\UUT/Mcontrol/st_logic/N94 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C165  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N94 ), .ZN(\UUT/Mcontrol/st_logic/N95 ) );
  INV_X2 \UUT/Mcontrol/st_logic/I_32  ( .A(\UUT/Mcontrol/st_logic/N95 ), .ZN(
        \UUT/Mcontrol/st_logic/N96 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C171  ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N98 ), .ZN(\UUT/Mcontrol/st_logic/N99 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C172  ( .A1(\UUT/Mcontrol/st_logic/N90 ), .A2(
        \UUT/Mcontrol/st_logic/N99 ), .ZN(\UUT/Mcontrol/st_logic/N100 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C173  ( .A1(\UUT/Mcontrol/d_jump_type[0] ), 
        .A2(\UUT/Mcontrol/st_logic/N100 ), .ZN(\UUT/Mcontrol/st_logic/N101 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C179  ( .A1(\UUT/Mcontrol/d_jump_type[2] ), 
        .A2(\UUT/Mcontrol/st_logic/N105 ), .ZN(\UUT/Mcontrol/st_logic/N106 )
         );
  OR2_X2 \UUT/Mcontrol/st_logic/C181  ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N107 ), .ZN(\UUT/Mcontrol/st_logic/N108 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C193  ( .A1(\UUT/Mcontrol/st_logic/N15 ), 
        .A2(\UUT/Mcontrol/st_logic/N110 ), .ZN(\UUT/Mcontrol/st_logic/N2 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C194  ( .A1(\UUT/Mcontrol/st_logic/N19 ), .A2(
        \UUT/Mcontrol/st_logic/N23 ), .ZN(\UUT/Mcontrol/st_logic/N110 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C198  ( .A1(\UUT/Mcontrol/st_logic/N111 ), 
        .A2(\UUT/Mcontrol/st_logic/N89 ), .ZN(\UUT/Mcontrol/st_logic/N112 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C199  ( .A1(\UUT/Mcontrol/st_logic/N77 ), .A2(
        \UUT/Mcontrol/st_logic/N83 ), .ZN(\UUT/Mcontrol/st_logic/N111 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C200  ( .A1(\UUT/Mcontrol/st_logic/N64 ), .A2(
        \UUT/Mcontrol/st_logic/N71 ), .ZN(\UUT/Mcontrol/st_logic/N4 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C204  ( .A1(\UUT/Mcontrol/st_logic/N24 ), 
        .A2(\UUT/Mcontrol/st_logic/N25 ), .ZN(\UUT/Mcontrol/st_logic/N6 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C205  ( .A1(\UUT/Mcontrol/st_logic/N117 ), 
        .A2(\UUT/Mcontrol/st_logic/N118 ), .ZN(\UUT/Mcontrol/st_logic/N7 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C206  ( .A1(\UUT/Mcontrol/st_logic/N54 ), 
        .A2(\UUT/Mcontrol/st_logic/N46 ), .ZN(\UUT/Mcontrol/st_logic/N117 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C207  ( .A1(\UUT/Mcontrol/st_logic/N57 ), 
        .A2(\UUT/Mcontrol/st_logic/N51 ), .ZN(\UUT/Mcontrol/st_logic/N118 ) );
  AND2_X2 \UUT/Mcontrol/st_logic/C208  ( .A1(\UUT/Mcontrol/st_logic/N119 ), 
        .A2(\UUT/Mcontrol/st_logic/N41 ), .ZN(\UUT/Mcontrol/st_logic/N8 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C209  ( .A1(\UUT/Mcontrol/st_logic/N33 ), .A2(
        \UUT/Mcontrol/st_logic/N40 ), .ZN(\UUT/Mcontrol/st_logic/N119 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C211  ( .A1(\UUT/Mcontrol/st_logic/N120 ), 
        .A2(\UUT/Mcontrol/st_logic/N14 ), .ZN(\UUT/Mcontrol/st_logic/N10 ) );
  OR2_X2 \UUT/Mcontrol/st_logic/C212  ( .A1(\UUT/Mcontrol/st_logic/N12 ), .A2(
        \UUT/Mcontrol/st_logic/N13 ), .ZN(\UUT/Mcontrol/st_logic/N120 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C19  ( .A1(\UUT/Mcontrol/x_rd[3] ), .A2(
        \UUT/Mcontrol/x_rd[4] ), .ZN(\UUT/Mcontrol/bp_logicB/N5 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C20  ( .A1(\UUT/Mcontrol/x_rd[2] ), .A2(
        \UUT/Mcontrol/bp_logicB/N5 ), .ZN(\UUT/Mcontrol/bp_logicB/N6 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C21  ( .A1(\UUT/Mcontrol/x_rd[1] ), .A2(
        \UUT/Mcontrol/bp_logicB/N6 ), .ZN(\UUT/Mcontrol/bp_logicB/N7 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C22  ( .A1(\UUT/Mcontrol/x_rd[0] ), .A2(
        \UUT/Mcontrol/bp_logicB/N7 ), .ZN(\UUT/Mcontrol/bp_logicB/N8 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C26  ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), 
        .A2(\UUT/Mcontrol/m_sampled_xrd[4] ), .ZN(\UUT/Mcontrol/bp_logicB/N10 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C27  ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N10 ), .ZN(\UUT/Mcontrol/bp_logicB/N11 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C28  ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N11 ), .ZN(\UUT/Mcontrol/bp_logicB/N12 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicB/C29  ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), 
        .A2(\UUT/Mcontrol/bp_logicB/N12 ), .ZN(\UUT/Mcontrol/bp_logicB/N13 )
         );
  INV_X2 \UUT/Mcontrol/bp_logicB/I_3  ( .A(\UUT/m_we ), .ZN(
        \UUT/Mcontrol/bp_logicB/N14 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C36  ( .A1(\UUT/Mcontrol/bp_logicB/N15 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N9 ), .ZN(
        \UUT/Mcontrol/bp_logicB/exec_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C37  ( .A1(\UUT/Mcontrol/bp_logicB/N2 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N8 ), .ZN(\UUT/Mcontrol/bp_logicB/N15 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C38  ( .A1(\UUT/Mcontrol/bp_logicB/N16 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N14 ), .ZN(
        \UUT/Mcontrol/bp_logicB/memory_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicB/C39  ( .A1(\UUT/Mcontrol/bp_logicB/N3 ), 
        .A2(\UUT/Mcontrol/bp_logicB/N13 ), .ZN(\UUT/Mcontrol/bp_logicB/N16 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C19  ( .A1(\UUT/Mcontrol/x_rd[3] ), .A2(
        \UUT/Mcontrol/x_rd[4] ), .ZN(\UUT/Mcontrol/bp_logicA/N5 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C20  ( .A1(\UUT/Mcontrol/x_rd[2] ), .A2(
        \UUT/Mcontrol/bp_logicA/N5 ), .ZN(\UUT/Mcontrol/bp_logicA/N6 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C21  ( .A1(\UUT/Mcontrol/x_rd[1] ), .A2(
        \UUT/Mcontrol/bp_logicA/N6 ), .ZN(\UUT/Mcontrol/bp_logicA/N7 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C22  ( .A1(\UUT/Mcontrol/x_rd[0] ), .A2(
        \UUT/Mcontrol/bp_logicA/N7 ), .ZN(\UUT/Mcontrol/bp_logicA/N8 ) );
  INV_X2 \UUT/Mcontrol/bp_logicA/I_1  ( .A(\UUT/x_we ), .ZN(
        \UUT/Mcontrol/bp_logicA/N9 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C26  ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), 
        .A2(\UUT/Mcontrol/m_sampled_xrd[4] ), .ZN(\UUT/Mcontrol/bp_logicA/N10 ) );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C27  ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N10 ), .ZN(\UUT/Mcontrol/bp_logicA/N11 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C28  ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N11 ), .ZN(\UUT/Mcontrol/bp_logicA/N12 )
         );
  OR2_X2 \UUT/Mcontrol/bp_logicA/C29  ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), 
        .A2(\UUT/Mcontrol/bp_logicA/N12 ), .ZN(\UUT/Mcontrol/bp_logicA/N13 )
         );
  INV_X2 \UUT/Mcontrol/bp_logicA/I_3  ( .A(\UUT/m_we ), .ZN(
        \UUT/Mcontrol/bp_logicA/N14 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C36  ( .A1(\UUT/Mcontrol/bp_logicA/N15 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N9 ), .ZN(
        \UUT/Mcontrol/bp_logicA/exec_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C37  ( .A1(\UUT/Mcontrol/bp_logicA/N2 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N8 ), .ZN(\UUT/Mcontrol/bp_logicA/N15 ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C38  ( .A1(\UUT/Mcontrol/bp_logicA/N16 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N14 ), .ZN(
        \UUT/Mcontrol/bp_logicA/memory_main ) );
  AND2_X2 \UUT/Mcontrol/bp_logicA/C39  ( .A1(\UUT/Mcontrol/bp_logicA/N3 ), 
        .A2(\UUT/Mcontrol/bp_logicA/N13 ), .ZN(\UUT/Mcontrol/bp_logicA/N16 )
         );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_0  ( .A(\UUT/Mcontrol/d_jump_type[3] ), .ZN(\UUT/Mcontrol/st_logic/N103 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C198  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N114 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N115 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_3  ( .A(\UUT/Mcontrol/d_jump_type[0] ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N120 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C208  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N122 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N123 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C210  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N124 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N125 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C223  ( .A1(\UUT/branch_rega [19]), 
        .A2(\UUT/Mcontrol/Nextpc_decoding/N137 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N138 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C224  ( .A1(\UUT/branch_rega [18]), 
        .A2(\UUT/Mcontrol/Nextpc_decoding/N138 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N139 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C225  ( .A1(\UUT/branch_rega [17]), 
        .A2(\UUT/Mcontrol/Nextpc_decoding/N139 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N140 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C226  ( .A1(\UUT/branch_rega [16]), 
        .A2(\UUT/Mcontrol/Nextpc_decoding/N140 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N141 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C227  ( .A1(\UUT/branch_rega [15]), 
        .A2(\UUT/Mcontrol/Nextpc_decoding/N141 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N142 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C283  ( .A1(n7186), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N127 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N194 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_10  ( .A(
        \UUT/Mcontrol/d_jump_type[2] ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N223 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C318  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N226 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N227 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C319  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N227 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N228 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C320  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N228 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N229 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_12  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N229 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N230 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C326  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N232 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N233 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C327  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N233 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N234 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C328  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N234 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N235 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C333  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N238 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N239 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C334  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N224 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N239 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N240 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C335  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N240 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N241 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C340  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N244 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N245 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C342  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N246 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N247 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_15  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N247 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N248 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C346  ( .A1(
        \UUT/Mcontrol/d_jump_type[2] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N250 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N251 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C348  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N252 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N253 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_16  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N253 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N254 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C354  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N256 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N257 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C356  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N120 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N258 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N259 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_17  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N259 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N260 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C361  ( .A1(
        \UUT/Mcontrol/Nextpc_decoding/N223 ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N262 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N263 ) );
  OR2_X2 \UUT/Mcontrol/Nextpc_decoding/C363  ( .A1(
        \UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N264 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N265 ) );
  INV_X2 \UUT/Mcontrol/Nextpc_decoding/I_18  ( .A(
        \UUT/Mcontrol/Nextpc_decoding/N265 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N266 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2058  ( .A1(
        \UUT/Mcontrol/d_sampled_finstr [4]), .A2(\UUT/Mcontrol/d_instr [5]), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1883 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2059  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1883 ), .A2(n7200), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1884 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2070  ( .A1(n7044), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1891 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1892 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2071  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1892 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1893 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2077  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1896 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1897 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2078  ( .A1(
        \UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1897 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1898 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_6  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1898 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1899 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2085  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1904 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1905 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2086  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1901 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1905 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1906 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_9  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1906 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1907 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2091  ( .A1(
        \UUT/Mcontrol/d_instr [1]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1910 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1911 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2092  ( .A1(
        \UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1911 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1912 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_10  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1912 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1913 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2094  ( .A1(
        \UUT/Mcontrol/d_instr [6]), .A2(\UUT/Mcontrol/d_instr [7]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1914 ) );
  INV_X2 \UUT/Mcontrol/Operation_decoding32/I_11  ( .A(
        \UUT/Mcontrol/Operation_decoding32/N1914 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1915 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2120  ( .A1(
        \UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1932 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1933 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2326  ( .A1(n7044), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2082 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2083 ) );
  OR2_X2 \UUT/Mcontrol/Operation_decoding32/C2327  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2083 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2084 ) );
  AND2_X2 \UUT/Mcontrol/Operation_decoding32/C2606  ( .A1(
        \UUT/Mcontrol/Operation_decoding32/N1913 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1915 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N62 ) );
  AND2_X2 \UUT/Mcontrol/C112  ( .A1(\UUT/Mcontrol/N19 ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(I_BUSY) );
  INV_X2 \UUT/BYP_BRANCH_MUXB/I_0  ( .A(\UUT/BYP_BRANCH_MUXB/N39 ), .ZN(
        \UUT/BYP_BRANCH_MUXB/N4 ) );
  INV_X2 \UUT/BYP_BRANCH_MUXB/I_1  ( .A(\UUT/byp_controlB[2] ), .ZN(
        \UUT/BYP_BRANCH_MUXB/N39 ) );
  OR2_X2 \UUT/regfile/C1390  ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/regfile/N261 ), 
        .ZN(\UUT/regfile/N262 ) );
  OR2_X2 \UUT/regfile/C1394  ( .A1(\UUT/rs2_addr [3]), .A2(\UUT/rs2_addr [4]), 
        .ZN(\UUT/regfile/N265 ) );
  OR2_X2 \UUT/regfile/C1395  ( .A1(\UUT/rs2_addr [2]), .A2(\UUT/regfile/N265 ), 
        .ZN(\UUT/regfile/N266 ) );
  OR2_X2 \UUT/regfile/C1396  ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/regfile/N266 ), 
        .ZN(\UUT/regfile/N267 ) );
  OR2_X2 \UUT/regfile/C1401  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N272 ) );
  OR2_X2 \UUT/regfile/C1402  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N272 ), 
        .ZN(\UUT/regfile/N273 ) );
  OR2_X2 \UUT/regfile/C1408  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N279 ) );
  OR2_X2 \UUT/regfile/C1409  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N279 ), 
        .ZN(\UUT/regfile/N280 ) );
  OR2_X2 \UUT/regfile/C1416  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N285 ) );
  OR2_X2 \UUT/regfile/C1417  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N285 ), 
        .ZN(\UUT/regfile/N286 ) );
  INV_X2 \UUT/regfile/I_7  ( .A(\UUT/rd_addr [2]), .ZN(\UUT/regfile/N290 ) );
  OR2_X2 \UUT/regfile/C1423  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N292 ) );
  OR2_X2 \UUT/regfile/C1424  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N292 ), .ZN(\UUT/regfile/N293 ) );
  OR2_X2 \UUT/regfile/C1431  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N298 ) );
  OR2_X2 \UUT/regfile/C1432  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N298 ), .ZN(\UUT/regfile/N299 ) );
  OR2_X2 \UUT/regfile/C1439  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N304 ) );
  OR2_X2 \UUT/regfile/C1440  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N304 ), .ZN(\UUT/regfile/N305 ) );
  OR2_X2 \UUT/regfile/C1448  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N358 ), 
        .ZN(\UUT/regfile/N310 ) );
  OR2_X2 \UUT/regfile/C1449  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N310 ), .ZN(\UUT/regfile/N311 ) );
  INV_X2 \UUT/regfile/I_12  ( .A(\UUT/rd_addr [3]), .ZN(\UUT/regfile/N315 ) );
  OR2_X2 \UUT/regfile/C1455  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N317 ) );
  OR2_X2 \UUT/regfile/C1456  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N317 ), 
        .ZN(\UUT/regfile/N318 ) );
  OR2_X2 \UUT/regfile/C1463  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N323 ) );
  OR2_X2 \UUT/regfile/C1464  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N323 ), 
        .ZN(\UUT/regfile/N324 ) );
  OR2_X2 \UUT/regfile/C1471  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N329 ) );
  OR2_X2 \UUT/regfile/C1472  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N329 ), 
        .ZN(\UUT/regfile/N330 ) );
  OR2_X2 \UUT/regfile/C1480  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N335 ) );
  OR2_X2 \UUT/regfile/C1481  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N335 ), 
        .ZN(\UUT/regfile/N336 ) );
  OR2_X2 \UUT/regfile/C1488  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N341 ) );
  OR2_X2 \UUT/regfile/C1489  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N341 ), .ZN(\UUT/regfile/N342 ) );
  OR2_X2 \UUT/regfile/C1497  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N347 ) );
  OR2_X2 \UUT/regfile/C1498  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N347 ), .ZN(\UUT/regfile/N348 ) );
  OR2_X2 \UUT/regfile/C1506  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N353 ) );
  OR2_X2 \UUT/regfile/C1507  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N353 ), .ZN(\UUT/regfile/N354 ) );
  OR2_X2 \UUT/regfile/C1516  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N359 ) );
  OR2_X2 \UUT/regfile/C1517  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N359 ), .ZN(\UUT/regfile/N360 ) );
  INV_X2 \UUT/regfile/I_21  ( .A(\UUT/regfile/N358 ), .ZN(\UUT/regfile/N455 )
         );
  OR2_X2 \UUT/regfile/C1523  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N366 ) );
  OR2_X2 \UUT/regfile/C1524  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N366 ), 
        .ZN(\UUT/regfile/N367 ) );
  OR2_X2 \UUT/regfile/C1531  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N372 ) );
  OR2_X2 \UUT/regfile/C1532  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N372 ), 
        .ZN(\UUT/regfile/N373 ) );
  OR2_X2 \UUT/regfile/C1539  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N378 ) );
  OR2_X2 \UUT/regfile/C1540  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N378 ), 
        .ZN(\UUT/regfile/N379 ) );
  OR2_X2 \UUT/regfile/C1548  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N384 ) );
  OR2_X2 \UUT/regfile/C1549  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N384 ), 
        .ZN(\UUT/regfile/N385 ) );
  OR2_X2 \UUT/regfile/C1556  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N390 ) );
  OR2_X2 \UUT/regfile/C1557  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N390 ), .ZN(\UUT/regfile/N391 ) );
  OR2_X2 \UUT/regfile/C1565  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N396 ) );
  OR2_X2 \UUT/regfile/C1566  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N396 ), .ZN(\UUT/regfile/N397 ) );
  OR2_X2 \UUT/regfile/C1574  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N402 ) );
  OR2_X2 \UUT/regfile/C1575  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N402 ), .ZN(\UUT/regfile/N403 ) );
  OR2_X2 \UUT/regfile/C1584  ( .A1(\UUT/rd_addr [3]), .A2(\UUT/regfile/N455 ), 
        .ZN(\UUT/regfile/N408 ) );
  OR2_X2 \UUT/regfile/C1585  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N408 ), .ZN(\UUT/regfile/N409 ) );
  OR2_X2 \UUT/regfile/C1592  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N414 ) );
  OR2_X2 \UUT/regfile/C1593  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N414 ), 
        .ZN(\UUT/regfile/N415 ) );
  OR2_X2 \UUT/regfile/C1601  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N420 ) );
  OR2_X2 \UUT/regfile/C1602  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N420 ), 
        .ZN(\UUT/regfile/N421 ) );
  OR2_X2 \UUT/regfile/C1610  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N426 ) );
  OR2_X2 \UUT/regfile/C1611  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N426 ), 
        .ZN(\UUT/regfile/N427 ) );
  OR2_X2 \UUT/regfile/C1620  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N432 ) );
  OR2_X2 \UUT/regfile/C1621  ( .A1(\UUT/rd_addr [2]), .A2(\UUT/regfile/N432 ), 
        .ZN(\UUT/regfile/N433 ) );
  OR2_X2 \UUT/regfile/C1629  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N438 ) );
  OR2_X2 \UUT/regfile/C1630  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N438 ), .ZN(\UUT/regfile/N439 ) );
  OR2_X2 \UUT/regfile/C1639  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N444 ) );
  OR2_X2 \UUT/regfile/C1640  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N444 ), .ZN(\UUT/regfile/N445 ) );
  OR2_X2 \UUT/regfile/C1649  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N450 ) );
  OR2_X2 \UUT/regfile/C1650  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N450 ), .ZN(\UUT/regfile/N451 ) );
  OR2_X2 \UUT/regfile/C1660  ( .A1(\UUT/regfile/N315 ), .A2(\UUT/regfile/N455 ), .ZN(\UUT/regfile/N456 ) );
  OR2_X2 \UUT/regfile/C1661  ( .A1(\UUT/regfile/N290 ), .A2(\UUT/regfile/N456 ), .ZN(\UUT/regfile/N457 ) );
  INV_X2 \UUT/I_2  ( .A(dmem_read), .ZN(\UUT/N76 ) );
  INV_X2 \UUT/I_3  ( .A(dmem_write), .ZN(\UUT/N77 ) );
  AND2_X2 C271 ( .A1(N40), .A2(N41), .ZN(N178) );
  AND2_X2 C270 ( .A1(N178), .A2(N172), .ZN(N42) );
  AND2_X2 C268 ( .A1(N37), .A2(N38), .ZN(N177) );
  AND2_X2 C267 ( .A1(N177), .A2(N171), .ZN(N43) );
  AND2_X2 C265 ( .A1(N33), .A2(N34), .ZN(N176) );
  AND2_X2 C264 ( .A1(N176), .A2(N168), .ZN(N35) );
  AND2_X2 C262 ( .A1(N29), .A2(N30), .ZN(N175) );
  AND2_X2 C261 ( .A1(N175), .A2(N165), .ZN(N31) );
  AND2_X2 C259 ( .A1(N24), .A2(N25), .ZN(N174) );
  AND2_X2 C258 ( .A1(N174), .A2(N26), .ZN(N27) );
  AND2_X2 C256 ( .A1(N19), .A2(N20), .ZN(N173) );
  AND2_X2 C255 ( .A1(N173), .A2(N21), .ZN(N22) );
  INV_X2 I_19 ( .A(I_BUSY), .ZN(iram_rd) );
  AND2_X2 C246 ( .A1(D_ADDR_OUTBUS[0]), .A2(D_ADDR_OUTBUS[1]), .ZN(N172) );
  INV_X2 I_18 ( .A(N170), .ZN(N171) );
  OR2_X2 C244 ( .A1(D_ADDR_OUTBUS[0]), .A2(N169), .ZN(N170) );
  INV_X2 I_17 ( .A(D_ADDR_OUTBUS[1]), .ZN(N169) );
  INV_X2 I_16 ( .A(N167), .ZN(N168) );
  OR2_X2 C241 ( .A1(N166), .A2(D_ADDR_OUTBUS[1]), .ZN(N167) );
  INV_X2 I_15 ( .A(D_ADDR_OUTBUS[0]), .ZN(N166) );
  INV_X2 I_14 ( .A(N164), .ZN(N165) );
  OR2_X2 C238 ( .A1(D_ADDR_OUTBUS[0]), .A2(D_ADDR_OUTBUS[1]), .ZN(N164) );
  INV_X2 I_13 ( .A(N13), .ZN(N41) );
  INV_X2 I_12 ( .A(N12), .ZN(N40) );
  INV_X2 I_11 ( .A(N11), .ZN(N38) );
  INV_X2 I_10 ( .A(N10), .ZN(N37) );
  INV_X2 I_9 ( .A(N9), .ZN(N34) );
  INV_X2 I_8 ( .A(N8), .ZN(N33) );
  INV_X2 I_7 ( .A(N7), .ZN(N30) );
  INV_X2 I_6 ( .A(N6), .ZN(N29) );
  INV_X2 I_5 ( .A(N5), .ZN(N26) );
  INV_X2 I_4 ( .A(N4), .ZN(N25) );
  INV_X2 I_3 ( .A(N3), .ZN(N24) );
  INV_X2 I_2 ( .A(N2), .ZN(N21) );
  INV_X2 I_1 ( .A(N1), .ZN(N20) );
  INV_X2 I_0 ( .A(N0), .ZN(N19) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[31]  ( .D(n4312), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[31] ), 
        .QN(n2835) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[63]  ( .D(n4311), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[63] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[62]  ( .D(n4310), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[62] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[61]  ( .D(n4309), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[61] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[60]  ( .D(n4308), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[60] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[59]  ( .D(n4307), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[59] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[58]  ( .D(n4306), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[58] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[56]  ( .D(n4304), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[56] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[55]  ( .D(n4303), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[55] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[54]  ( .D(n4302), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[54] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[53]  ( .D(n4301), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[53] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[52]  ( .D(n4300), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[52] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[51]  ( .D(n4299), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[51] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[50]  ( .D(n4298), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[50] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[49]  ( .D(n4297), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[49] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[48]  ( .D(n4296), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[48] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[47]  ( .D(n4295), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[47] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[46]  ( .D(n4294), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[46] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[45]  ( .D(n4293), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[45] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[44]  ( .D(n4292), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[44] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[43]  ( .D(n4291), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[43] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[42]  ( .D(n4290), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[42] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[41]  ( .D(n4289), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[41] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[40]  ( .D(n4288), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[40] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[39]  ( .D(n4287), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[39] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[38]  ( .D(n4286), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[38] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[37]  ( .D(n4285), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[37] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[36]  ( .D(n4284), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[36] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[35]  ( .D(n4283), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[35] ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[34]  ( .D(n4282), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[34] ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][0]  ( .D(n4247), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][0] ), .QN(
        \UUT/Mpath/the_alu/N468 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[31]  ( .D(n4246), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [31]), 
        .QN(n7228) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[30]  ( .D(n4243), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [30]), 
        .QN(n7237) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[29]  ( .D(n4242), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [29]), 
        .QN(n7216) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[1]  ( .D(n4238), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [1]), .QN(
        \UUT/Mpath/N116 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[0]  ( .D(n4237), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [0]), .QN(
        \UUT/Mpath/N112 ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MW]  ( .D(n4235), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[MW] ), .QN(n2761) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[5]  ( .D(n4211), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [5]), 
        .QN(n7217) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[5]  ( .D(n4210), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [5]), 
        .QN(n2736) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[5]  ( .D(n4208), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[5] ), .QN(n2734) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][5]  ( .D(n4207), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][5] ), .QN(
        \UUT/Mpath/the_alu/N466 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[4]  ( .D(n4206), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [4]), 
        .QN(n7221) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[4]  ( .D(n4205), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [4]), 
        .QN(n2732) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[4]  ( .D(n4203), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[4] ), .QN(n2730) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][4]  ( .D(n4202), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][4] ), .QN(
        \UUT/Mpath/the_alu/N453 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[3]  ( .D(n4201), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [3]), 
        .QN(n7199) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[3]  ( .D(n4200), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [3]), 
        .QN(n2728) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[3]  ( .D(n4199), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[3] ), .QN(\UUT/Mpath/the_mult/N192 )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[3]  ( .D(n4198), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[3] ), .QN(\UUT/Mpath/the_mult/N229 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][3]  ( .D(n4197), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][3] ), .QN(n2727) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[2]  ( .D(n4196), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [2]), 
        .QN(n7210) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[2]  ( .D(n4195), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mcontrol/st_logic/N26 ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[2]  ( .D(n4193), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[2] ), .QN(\UUT/Mpath/the_mult/N244 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[2]  ( .D(n4192), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [2]), .QN(
        \UUT/Mpath/the_shift/N104 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][2]  ( .D(n4191), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][2] ), .QN(n2724) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[1]  ( .D(n4190), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [1]), 
        .QN(n7188) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[1]  ( .D(n4189), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mcontrol/st_logic/N27 ) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[1]  ( .D(n4187), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[1] ), .QN(\UUT/Mpath/the_mult/N230 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[1]  ( .D(n4186), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [1]), .QN(
        \UUT/Mpath/the_shift/N112 ) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[0]  ( .D(n4185), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [0]), 
        .QN(n7139) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[0]  ( .D(n4184), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_mul_command [0]), 
        .QN(\UUT/Mcontrol/st_logic/N34 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[0]  ( .D(n4183), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[0] ), .QN(\UUT/Mpath/the_mult/N193 )
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[0]  ( .D(n4182), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/m_mul_command[0] ), .QN(\UUT/Mpath/the_mult/N231 )
         );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[0]  ( .D(n4181), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/shift_op [0]), .QN(
        \UUT/Mpath/the_shift/N105 ) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[4]  ( .D(n4179), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[4] ), .QN(
        n2719) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[3]  ( .D(n4177), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[3] ), .QN(
        n2717) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[2]  ( .D(n4175), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[2] ), .QN(
        n2715) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[1]  ( .D(n4173), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[1] ), .QN(
        n2713) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_rf_we_reg  ( .D(n4172), .CK(CLK), .SN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/x_we ), .QN(
        \UUT/Mcontrol/bp_logicB/N9 ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_rf_we_reg  ( .D(n4171), .CK(CLK), .SN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/m_we ), .QN(n5315) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[SIGN]  ( .D(n4170), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/m_mem_command[SIGN] ), .QN(
        \UUT/Mpath/the_memhandle/N235 ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MH]  ( .D(n4168), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mpath/the_memhandle/N238 ) );
  DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MB]  ( .D(n4167), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(\UUT/Mpath/the_memhandle/N236 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][1]  ( .D(n4165), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Alu_command[OP][1] ), .QN(
        \UUT/Mpath/the_alu/N467 ) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[2]  ( .D(n4164), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/exe_outsel [2]), .QN(
        \UUT/Mpath/N111 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[0]  ( .D(n4162), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[0] ), .QN(
        \UUT/Mpath/the_alu/N84 ) );
  DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[0]  ( .D(n4161), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/mem_baddr [0]), .QN(
        \UUT/Mpath/the_memhandle/N240 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[10]  ( .D(n4160), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [10]), .QN(
        n2711) );
  DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[0]  ( .D(n4157), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [0]), .QN(
        n2709) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[23]  ( .D(n4132), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[23] ), .QN(
        \UUT/Mpath/the_alu/N38 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[31]  ( .D(n4130), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[31] ), .QN(
        \UUT/Mpath/the_alu/N22 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[30]  ( .D(n4128), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[30] ), .QN(
        \UUT/Mpath/the_alu/N23 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[30]  ( .D(n4127), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[30] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[30]  ( .D(n4125), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[62] ), .QN(
        n5599) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[30]  ( .D(n4124), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[30] ), .QN(
        n5543) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[29]  ( .D(n4123), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[61] ), .QN(
        n5601) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[28]  ( .D(n4119), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[28] ), .QN(
        \UUT/Mpath/the_alu/N27 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[27]  ( .D(n4117), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[27] ), .QN(
        \UUT/Mpath/the_alu/N29 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[26]  ( .D(n4115), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[26] ), .QN(
        \UUT/Mpath/the_alu/N31 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[25]  ( .D(n4113), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[25] ), .QN(
        \UUT/Mpath/the_alu/N33 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[1]  ( .D(n4111), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[1] ), .QN(
        \UUT/Mpath/the_alu/N82 ) );
  DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[1]  ( .D(n4110), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/mem_baddr [1]), .QN(
        \UUT/Mpath/the_memhandle/N239 ) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[31]  ( .D(n4105), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][31] ), .QN(n4458) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[31]  ( .D(n4104), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][31] ), .QN(n4490) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[31]  ( .D(n4099), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][31] ), .QN(
        n4650) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[31]  ( .D(n4098), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][31] ), .QN(
        n4682) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[31]  ( .D(n4095), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][31] ), .QN(
        n4778) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[31]  ( .D(n4094), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][31] ), .QN(
        n4810) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[31]  ( .D(n4091), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][31] ), .QN(
        n4906) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[31]  ( .D(n4090), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][31] ), .QN(
        n4938) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[31]  ( .D(n4088), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][31] ), .QN(
        n5002) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[31]  ( .D(n4087), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][31] ), .QN(
        n5034) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[31]  ( .D(n4078), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[31] ), .QN(
        \UUT/Mpath/the_alu/N21 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[31]  ( .D(n4077), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[31] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[31]  ( .D(n4075), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[31] ), .QN(
        n5541) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[30]  ( .D(n4070), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][30] ), .QN(n4459) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[30]  ( .D(n4069), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][30] ), .QN(n4491) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[30]  ( .D(n4064), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][30] ), .QN(
        n4651) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[30]  ( .D(n4063), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][30] ), .QN(
        n4683) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[30]  ( .D(n4060), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][30] ), .QN(
        n4779) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[30]  ( .D(n4059), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][30] ), .QN(
        n4811) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[30]  ( .D(n4056), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][30] ), .QN(
        n4907) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[30]  ( .D(n4055), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][30] ), .QN(
        n4939) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[30]  ( .D(n4053), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][30] ), .QN(
        n5003) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[30]  ( .D(n4052), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][30] ), .QN(
        n5035) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[29]  ( .D(n4039), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][29] ), .QN(n4461) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[29]  ( .D(n4038), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][29] ), .QN(n4493) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[29]  ( .D(n4033), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][29] ), .QN(
        n4653) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[29]  ( .D(n4032), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][29] ), .QN(
        n4685) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[29]  ( .D(n4029), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][29] ), .QN(
        n4781) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[29]  ( .D(n4028), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][29] ), .QN(
        n4813) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[29]  ( .D(n4025), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][29] ), .QN(
        n4909) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[29]  ( .D(n4024), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][29] ), .QN(
        n4941) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[29]  ( .D(n4022), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][29] ), .QN(
        n5005) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[29]  ( .D(n4021), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][29] ), .QN(
        n5037) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[28]  ( .D(n4008), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][28] ), .QN(n4462) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[28]  ( .D(n4007), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][28] ), .QN(n4494) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[28]  ( .D(n4002), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][28] ), .QN(
        n4654) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[28]  ( .D(n4001), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][28] ), .QN(
        n4686) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[28]  ( .D(n3998), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][28] ), .QN(
        n4782) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[28]  ( .D(n3997), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][28] ), .QN(
        n4814) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[28]  ( .D(n3994), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][28] ), .QN(
        n4910) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[28]  ( .D(n3993), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][28] ), .QN(
        n4942) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[28]  ( .D(n3991), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][28] ), .QN(
        n5006) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[28]  ( .D(n3990), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][28] ), .QN(
        n5038) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[27]  ( .D(n3977), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][27] ), .QN(n4463) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[27]  ( .D(n3976), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][27] ), .QN(n4495) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[27]  ( .D(n3971), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][27] ), .QN(
        n4655) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[27]  ( .D(n3970), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][27] ), .QN(
        n4687) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[27]  ( .D(n3967), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][27] ), .QN(
        n4783) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[27]  ( .D(n3966), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][27] ), .QN(
        n4815) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[27]  ( .D(n3963), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][27] ), .QN(
        n4911) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[27]  ( .D(n3962), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][27] ), .QN(
        n4943) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[27]  ( .D(n3960), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][27] ), .QN(
        n5007) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[27]  ( .D(n3959), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][27] ), .QN(
        n5039) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[26]  ( .D(n3946), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][26] ), .QN(n4464) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[26]  ( .D(n3945), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][26] ), .QN(n4496) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[26]  ( .D(n3940), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][26] ), .QN(
        n4656) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[26]  ( .D(n3939), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][26] ), .QN(
        n4688) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[26]  ( .D(n3936), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][26] ), .QN(
        n4784) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[26]  ( .D(n3935), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][26] ), .QN(
        n4816) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[26]  ( .D(n3932), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][26] ), .QN(
        n4912) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[26]  ( .D(n3931), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][26] ), .QN(
        n4944) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[26]  ( .D(n3929), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][26] ), .QN(
        n5008) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[26]  ( .D(n3928), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][26] ), .QN(
        n5040) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[25]  ( .D(n3915), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][25] ), .QN(n4465) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[25]  ( .D(n3914), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][25] ), .QN(n4497) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[25]  ( .D(n3909), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][25] ), .QN(
        n4657) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[25]  ( .D(n3908), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][25] ), .QN(
        n4689) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[25]  ( .D(n3905), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][25] ), .QN(
        n4785) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[25]  ( .D(n3904), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][25] ), .QN(
        n4817) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[25]  ( .D(n3901), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][25] ), .QN(
        n4913) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[25]  ( .D(n3900), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][25] ), .QN(
        n4945) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[25]  ( .D(n3898), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][25] ), .QN(
        n5009) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[25]  ( .D(n3897), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][25] ), .QN(
        n5041) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[23]  ( .D(n3884), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][23] ), .QN(n4467) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[23]  ( .D(n3883), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][23] ), .QN(n4499) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[23]  ( .D(n3878), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][23] ), .QN(
        n4659) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[23]  ( .D(n3877), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][23] ), .QN(
        n4691) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[23]  ( .D(n3874), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][23] ), .QN(
        n4787) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[23]  ( .D(n3873), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][23] ), .QN(
        n4819) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[23]  ( .D(n3870), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][23] ), .QN(
        n4915) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[23]  ( .D(n3869), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][23] ), .QN(
        n4947) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[23]  ( .D(n3867), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][23] ), .QN(
        n5011) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[23]  ( .D(n3866), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][23] ), .QN(
        n5043) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[23]  ( .D(n3857), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[23] ), .QN(
        \UUT/Mpath/the_alu/N37 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[23]  ( .D(n3856), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[23] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[23]  ( .D(n3854), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[23] ), .QN(
        n5559) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[23]  ( .D(n3853), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[55] ), .QN(
        n5607) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[1]  ( .D(n3848), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][1] ), .QN(n4471)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[1]  ( .D(n3847), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][1] ), .QN(n4503)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[1]  ( .D(n3842), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][1] ), .QN(n4663) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[1]  ( .D(n3841), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][1] ), .QN(n4695) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[1]  ( .D(n3838), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][1] ), .QN(n4791) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[1]  ( .D(n3837), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][1] ), .QN(n4823) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[1]  ( .D(n3834), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][1] ), .QN(n4919) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[1]  ( .D(n3833), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][1] ), .QN(n4951) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[1]  ( .D(n3831), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][1] ), .QN(n5015) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[1]  ( .D(n3830), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][1] ), .QN(n5047) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[1]  ( .D(n3821), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[1] ), .QN(
        \UUT/Mpath/the_alu/N81 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[1]  ( .D(n3820), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[1] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[1]  ( .D(n3818), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[1] ), 
        .QN(n5567) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[1]  ( .D(n3817), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[33] ), 
        .QN(n5611) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[0]  ( .D(n3812), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][0] ), .QN(n4482)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[0]  ( .D(n3811), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][0] ), .QN(n4514)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[0]  ( .D(n3806), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][0] ), .QN(n4674) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[0]  ( .D(n3805), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][0] ), .QN(n4706) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[0]  ( .D(n3802), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][0] ), .QN(n4802) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[0]  ( .D(n3801), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][0] ), .QN(n4834) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[0]  ( .D(n3798), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][0] ), .QN(n4930) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[0]  ( .D(n3797), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][0] ), .QN(n4962) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[0]  ( .D(n3795), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][0] ), .QN(n5026) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[0]  ( .D(n3794), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][0] ), .QN(n5058) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[0]  ( .D(n3782), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[0] ), 
        .QN(n5589) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[0]  ( .D(n3781), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[32] ), 
        .QN(n5622) );
  DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[1]  ( .D(n3780), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [1]), .QN(
        n2703) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[2]  ( .D(n3773), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][2] ), .QN(n4460)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[2]  ( .D(n3772), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][2] ), .QN(n4492)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[2]  ( .D(n3767), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][2] ), .QN(n4652) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[2]  ( .D(n3766), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][2] ), .QN(n4684) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[2]  ( .D(n3763), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][2] ), .QN(n4780) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[2]  ( .D(n3762), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][2] ), .QN(n4812) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[2]  ( .D(n3759), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][2] ), .QN(n4908) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[2]  ( .D(n3758), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][2] ), .QN(n4940) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[2]  ( .D(n3756), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][2] ), .QN(n5004) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[2]  ( .D(n3755), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][2] ), .QN(n5036) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[2]  ( .D(n3745), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[2] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[2]  ( .D(n3743), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[2] ), 
        .QN(n5545) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[2]  ( .D(n3742), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[34] ), 
        .QN(n5600) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[2]  ( .D(n3741), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[2] ), .QN(
        \UUT/Mpath/the_alu/N80 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[2]  ( .D(n3740), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [2])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[2]  ( .D(n3739), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [2]), .QN(
        n2699) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[3]  ( .D(n3733), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][3] ), .QN(n4457)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[3]  ( .D(n3732), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][3] ), .QN(n4489)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[3]  ( .D(n3727), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][3] ), .QN(n4649) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[3]  ( .D(n3726), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][3] ), .QN(n4681) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[3]  ( .D(n3723), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][3] ), .QN(n4777) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[3]  ( .D(n3722), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][3] ), .QN(n4809) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[3]  ( .D(n3719), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][3] ), .QN(n4905) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[3]  ( .D(n3718), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][3] ), .QN(n4937) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[3]  ( .D(n3716), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][3] ), .QN(n5001) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[3]  ( .D(n3715), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][3] ), .QN(n5033) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[3]  ( .D(n3706), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[3] ), .QN(
        \UUT/Mpath/the_alu/N77 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[3]  ( .D(n3705), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[3] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[3]  ( .D(n3703), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[3] ), 
        .QN(n5539) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[3]  ( .D(n3701), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[3] ), .QN(
        \UUT/Mpath/the_alu/N78 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[3]  ( .D(n3699), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [3]), .QN(
        n2696) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[4]  ( .D(n3693), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][4] ), .QN(n4456)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[4]  ( .D(n3692), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][4] ), .QN(n4488)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[4]  ( .D(n3687), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][4] ), .QN(n4648) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[4]  ( .D(n3686), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][4] ), .QN(n4680) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[4]  ( .D(n3683), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][4] ), .QN(n4776) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[4]  ( .D(n3682), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][4] ), .QN(n4808) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[4]  ( .D(n3679), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][4] ), .QN(n4904) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[4]  ( .D(n3678), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][4] ), .QN(n4936) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[4]  ( .D(n3676), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][4] ), .QN(n5000) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[4]  ( .D(n3675), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][4] ), .QN(n5032) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[4]  ( .D(n3666), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[4] ), .QN(
        \UUT/Mpath/the_alu/N75 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[4]  ( .D(n3665), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[4] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[4]  ( .D(n3663), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[4] ), 
        .QN(n5537) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[4]  ( .D(n3662), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[36] ), 
        .QN(n5596) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[4]  ( .D(n3661), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[4] ), .QN(
        \UUT/Mpath/the_alu/N76 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[4]  ( .D(n3660), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [4])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[4]  ( .D(n3659), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [4]), .QN(
        n2693) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[5]  ( .D(n3653), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][5] ), .QN(n4455)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[5]  ( .D(n3652), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][5] ), .QN(n4487)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[5]  ( .D(n3647), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][5] ), .QN(n4647) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[5]  ( .D(n3646), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][5] ), .QN(n4679) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[5]  ( .D(n3643), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][5] ), .QN(n4775) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[5]  ( .D(n3642), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][5] ), .QN(n4807) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[5]  ( .D(n3639), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][5] ), .QN(n4903) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[5]  ( .D(n3638), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][5] ), .QN(n4935) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[5]  ( .D(n3636), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][5] ), .QN(n4999) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[5]  ( .D(n3635), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][5] ), .QN(n5031) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[5]  ( .D(n3625), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[5] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[5]  ( .D(n3623), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[5] ), 
        .QN(n5535) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[5]  ( .D(n3622), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[37] ), 
        .QN(n5595) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[5]  ( .D(n3619), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [5]), .QN(
        n2690) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[6]  ( .D(n3613), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][6] ), .QN(n4454)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[6]  ( .D(n3612), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][6] ), .QN(n4486)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[6]  ( .D(n3607), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][6] ), .QN(n4646) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[6]  ( .D(n3606), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][6] ), .QN(n4678) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[6]  ( .D(n3603), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][6] ), .QN(n4774) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[6]  ( .D(n3602), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][6] ), .QN(n4806) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[6]  ( .D(n3599), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][6] ), .QN(n4902) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[6]  ( .D(n3598), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][6] ), .QN(n4934) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[6]  ( .D(n3596), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][6] ), .QN(n4998) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[6]  ( .D(n3595), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][6] ), .QN(n5030) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[6]  ( .D(n3585), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[6] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[6]  ( .D(n3583), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[6] ), 
        .QN(n5533) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[6]  ( .D(n3582), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[38] ), 
        .QN(n5594) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[6]  ( .D(n3580), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [6])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[7]  ( .D(n3573), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][7] ), .QN(n4453)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[7]  ( .D(n3572), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][7] ), .QN(n4485)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[7]  ( .D(n3567), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][7] ), .QN(n4645) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[7]  ( .D(n3566), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][7] ), .QN(n4677) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[7]  ( .D(n3563), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][7] ), .QN(n4773) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[7]  ( .D(n3562), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][7] ), .QN(n4805) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[7]  ( .D(n3559), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][7] ), .QN(n4901) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[7]  ( .D(n3558), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][7] ), .QN(n4933) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[7]  ( .D(n3556), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][7] ), .QN(n4997) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[7]  ( .D(n3555), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][7] ), .QN(n5029) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[7]  ( .D(n3545), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[7] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[7]  ( .D(n3543), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[7] ), 
        .QN(n5531) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[7]  ( .D(n3542), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[39] ), 
        .QN(n5593) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[7]  ( .D(n3541), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[7] ), .QN(
        \UUT/Mpath/the_alu/N70 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[7]  ( .D(n3539), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [7]), .QN(
        n2684) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[8]  ( .D(n3533), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][8] ), .QN(n4452)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[8]  ( .D(n3532), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][8] ), .QN(n4484)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[8]  ( .D(n3527), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][8] ), .QN(n4644) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[8]  ( .D(n3526), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][8] ), .QN(n4676) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[8]  ( .D(n3523), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][8] ), .QN(n4772) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[8]  ( .D(n3522), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][8] ), .QN(n4804) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[8]  ( .D(n3519), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][8] ), .QN(n4900) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[8]  ( .D(n3518), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][8] ), .QN(n4932) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[8]  ( .D(n3516), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][8] ), .QN(n4996) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[8]  ( .D(n3515), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][8] ), .QN(n5028) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[8]  ( .D(n3505), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[8] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[8]  ( .D(n3503), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[8] ), 
        .QN(n5529) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[8]  ( .D(n3502), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[40] ), 
        .QN(n5592) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[8]  ( .D(n3501), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[8] ), .QN(
        \UUT/Mpath/the_alu/N68 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[8]  ( .D(n3500), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [8])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[8]  ( .D(n3499), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [8]), .QN(
        n2681) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[9]  ( .D(n3493), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][9] ), .QN(n4451)
         );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[9]  ( .D(n3492), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][9] ), .QN(n4483)
         );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[9]  ( .D(n3487), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][9] ), .QN(n4643) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[9]  ( .D(n3486), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][9] ), .QN(n4675) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[9]  ( .D(n3483), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][9] ), .QN(n4771) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[9]  ( .D(n3482), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][9] ), .QN(n4803) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[9]  ( .D(n3479), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][9] ), .QN(n4899) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[9]  ( .D(n3478), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][9] ), .QN(n4931) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[9]  ( .D(n3476), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][9] ), .QN(n4995) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[9]  ( .D(n3475), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][9] ), .QN(n5027) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[9]  ( .D(n3465), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[9] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[9]  ( .D(n3463), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[9] ), 
        .QN(n5527) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[9]  ( .D(n3462), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[41] ), 
        .QN(n5591) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[9]  ( .D(n3461), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[9] ), .QN(
        \UUT/Mpath/the_alu/N66 ) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[10]  ( .D(n3454), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][10] ), .QN(n4481) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[10]  ( .D(n3453), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][10] ), .QN(n4513) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[10]  ( .D(n3448), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][10] ), .QN(
        n4673) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[10]  ( .D(n3447), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][10] ), .QN(
        n4705) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[10]  ( .D(n3444), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][10] ), .QN(
        n4801) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[10]  ( .D(n3443), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][10] ), .QN(
        n4833) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[10]  ( .D(n3440), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][10] ), .QN(
        n4929) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[10]  ( .D(n3439), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][10] ), .QN(
        n4961) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[10]  ( .D(n3437), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][10] ), .QN(
        n5025) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[10]  ( .D(n3436), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][10] ), .QN(
        n5057) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[10]  ( .D(n3426), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[10] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[10]  ( .D(n3424), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[10] ), .QN(
        n5587) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[10]  ( .D(n3423), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[42] ), .QN(
        n5621) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[10]  ( .D(n3421), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [10])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[11]  ( .D(n3415), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][11] ), .QN(n4480) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[11]  ( .D(n3414), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][11] ), .QN(n4512) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[11]  ( .D(n3409), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][11] ), .QN(
        n4672) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[11]  ( .D(n3408), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][11] ), .QN(
        n4704) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[11]  ( .D(n3405), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][11] ), .QN(
        n4800) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[11]  ( .D(n3404), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][11] ), .QN(
        n4832) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[11]  ( .D(n3401), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][11] ), .QN(
        n4928) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[11]  ( .D(n3400), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][11] ), .QN(
        n4960) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[11]  ( .D(n3398), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][11] ), .QN(
        n5024) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[11]  ( .D(n3397), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][11] ), .QN(
        n5056) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[11]  ( .D(n3387), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[11] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[11]  ( .D(n3385), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[11] ), .QN(
        n5585) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[11]  ( .D(n3384), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[43] ), .QN(
        n5620) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[11]  ( .D(n3383), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[11] ), .QN(
        \UUT/Mpath/the_alu/N62 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[11]  ( .D(n3381), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [11]), .QN(
        n2674) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[12]  ( .D(n3375), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][12] ), .QN(n4479) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[12]  ( .D(n3374), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][12] ), .QN(n4511) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[12]  ( .D(n3369), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][12] ), .QN(
        n4671) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[12]  ( .D(n3368), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][12] ), .QN(
        n4703) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[12]  ( .D(n3365), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][12] ), .QN(
        n4799) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[12]  ( .D(n3364), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][12] ), .QN(
        n4831) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[12]  ( .D(n3361), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][12] ), .QN(
        n4927) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[12]  ( .D(n3360), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][12] ), .QN(
        n4959) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[12]  ( .D(n3358), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][12] ), .QN(
        n5023) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[12]  ( .D(n3357), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][12] ), .QN(
        n5055) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[12]  ( .D(n3347), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[12] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[12]  ( .D(n3345), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[12] ), .QN(
        n5583) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[12]  ( .D(n3344), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[44] ), .QN(
        n5619) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[12]  ( .D(n3342), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [12])
         );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[12]  ( .D(n3341), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [12]), .QN(
        n2671) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[13]  ( .D(n3335), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][13] ), .QN(n4478) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[13]  ( .D(n3334), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][13] ), .QN(n4510) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[13]  ( .D(n3329), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][13] ), .QN(
        n4670) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[13]  ( .D(n3328), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][13] ), .QN(
        n4702) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[13]  ( .D(n3325), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][13] ), .QN(
        n4798) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[13]  ( .D(n3324), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][13] ), .QN(
        n4830) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[13]  ( .D(n3321), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][13] ), .QN(
        n4926) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[13]  ( .D(n3320), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][13] ), .QN(
        n4958) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[13]  ( .D(n3318), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][13] ), .QN(
        n5022) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[13]  ( .D(n3317), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][13] ), .QN(
        n5054) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[13]  ( .D(n3307), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[13] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[13]  ( .D(n3305), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[13] ), .QN(
        n5581) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[13]  ( .D(n3304), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[45] ), .QN(
        n5618) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[13]  ( .D(n3302), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [13]), .QN(
        n2669) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[14]  ( .D(n3295), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][14] ), .QN(n4477) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[14]  ( .D(n3294), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][14] ), .QN(n4509) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[14]  ( .D(n3289), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][14] ), .QN(
        n4669) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[14]  ( .D(n3288), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][14] ), .QN(
        n4701) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[14]  ( .D(n3285), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][14] ), .QN(
        n4797) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[14]  ( .D(n3284), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][14] ), .QN(
        n4829) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[14]  ( .D(n3281), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][14] ), .QN(
        n4925) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[14]  ( .D(n3280), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][14] ), .QN(
        n4957) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[14]  ( .D(n3278), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][14] ), .QN(
        n5021) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[14]  ( .D(n3277), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][14] ), .QN(
        n5053) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[14]  ( .D(n3267), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[14] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[14]  ( .D(n3265), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[14] ), .QN(
        n5579) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[14]  ( .D(n3264), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[46] ), .QN(
        n5617) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[14]  ( .D(n3262), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [14]), .QN(
        n2666) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[14]  ( .D(n3261), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [14])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[15]  ( .D(n3255), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][15] ), .QN(n4476) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[15]  ( .D(n3254), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][15] ), .QN(n4508) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[15]  ( .D(n3249), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][15] ), .QN(
        n4668) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[15]  ( .D(n3248), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][15] ), .QN(
        n4700) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[15]  ( .D(n3245), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][15] ), .QN(
        n4796) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[15]  ( .D(n3244), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][15] ), .QN(
        n4828) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[15]  ( .D(n3241), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][15] ), .QN(
        n4924) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[15]  ( .D(n3240), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][15] ), .QN(
        n4956) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[15]  ( .D(n3238), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][15] ), .QN(
        n5020) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[15]  ( .D(n3237), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][15] ), .QN(
        n5052) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[15]  ( .D(n3227), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[15] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[15]  ( .D(n3225), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[15] ), .QN(
        n5577) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[15]  ( .D(n3224), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[47] ), .QN(
        n5616) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[15]  ( .D(n3223), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[15] ), .QN(
        \UUT/Mpath/the_alu/N54 ) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[16]  ( .D(n3215), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][16] ), .QN(n4475) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[16]  ( .D(n3214), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][16] ), .QN(n4507) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[16]  ( .D(n3209), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][16] ), .QN(
        n4667) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[16]  ( .D(n3208), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][16] ), .QN(
        n4699) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[16]  ( .D(n3205), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][16] ), .QN(
        n4795) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[16]  ( .D(n3204), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][16] ), .QN(
        n4827) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[16]  ( .D(n3201), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][16] ), .QN(
        n4923) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[16]  ( .D(n3200), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][16] ), .QN(
        n4955) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[16]  ( .D(n3198), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][16] ), .QN(
        n5019) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[16]  ( .D(n3197), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][16] ), .QN(
        n5051) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[16]  ( .D(n3187), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[16] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[16]  ( .D(n3185), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[16] ), .QN(
        n5575) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[16]  ( .D(n3184), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[48] ), .QN(
        n5615) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[16]  ( .D(n3183), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[16] ), .QN(
        \UUT/Mpath/the_alu/N52 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[16]  ( .D(n3182), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [16]), .QN(
        n2660) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[16]  ( .D(n3181), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [16])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[17]  ( .D(n3175), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][17] ), .QN(n4474) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[17]  ( .D(n3174), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][17] ), .QN(n4506) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[17]  ( .D(n3169), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][17] ), .QN(
        n4666) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[17]  ( .D(n3168), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][17] ), .QN(
        n4698) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[17]  ( .D(n3165), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][17] ), .QN(
        n4794) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[17]  ( .D(n3164), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][17] ), .QN(
        n4826) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[17]  ( .D(n3161), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][17] ), .QN(
        n4922) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[17]  ( .D(n3160), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][17] ), .QN(
        n4954) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[17]  ( .D(n3158), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][17] ), .QN(
        n5018) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[17]  ( .D(n3157), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][17] ), .QN(
        n5050) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[17]  ( .D(n3147), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[17] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[17]  ( .D(n3145), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[17] ), .QN(
        n5573) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[17]  ( .D(n3144), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[49] ), .QN(
        n5614) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[17]  ( .D(n3143), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[17] ), .QN(
        \UUT/Mpath/the_alu/N50 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[17]  ( .D(n3142), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [17]), .QN(
        n2657) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[18]  ( .D(n3135), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][18] ), .QN(n4473) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[18]  ( .D(n3134), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][18] ), .QN(n4505) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[18]  ( .D(n3129), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][18] ), .QN(
        n4665) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[18]  ( .D(n3128), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][18] ), .QN(
        n4697) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[18]  ( .D(n3125), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][18] ), .QN(
        n4793) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[18]  ( .D(n3124), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][18] ), .QN(
        n4825) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[18]  ( .D(n3121), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][18] ), .QN(
        n4921) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[18]  ( .D(n3120), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][18] ), .QN(
        n4953) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[18]  ( .D(n3118), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][18] ), .QN(
        n5017) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[18]  ( .D(n3117), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][18] ), .QN(
        n5049) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[18]  ( .D(n3107), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[18] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[18]  ( .D(n3105), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[18] ), .QN(
        n5571) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[18]  ( .D(n3104), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[50] ), .QN(
        n5613) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[18]  ( .D(n3102), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [18]), .QN(
        n2654) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[18]  ( .D(n3101), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [18])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[19]  ( .D(n3095), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][19] ), .QN(n4472) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[19]  ( .D(n3094), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][19] ), .QN(n4504) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[19]  ( .D(n3089), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][19] ), .QN(
        n4664) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[19]  ( .D(n3088), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][19] ), .QN(
        n4696) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[19]  ( .D(n3085), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][19] ), .QN(
        n4792) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[19]  ( .D(n3084), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][19] ), .QN(
        n4824) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[19]  ( .D(n3081), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][19] ), .QN(
        n4920) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[19]  ( .D(n3080), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][19] ), .QN(
        n4952) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[19]  ( .D(n3078), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][19] ), .QN(
        n5016) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[19]  ( .D(n3077), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][19] ), .QN(
        n5048) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[19]  ( .D(n3067), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[19] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[19]  ( .D(n3065), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[19] ), .QN(
        n5569) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[19]  ( .D(n3064), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[51] ), .QN(
        n5612) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[19]  ( .D(n3063), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[19] ), .QN(
        \UUT/Mpath/the_alu/N46 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[19]  ( .D(n3062), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [19]), .QN(
        n2651) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[20]  ( .D(n3055), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][20] ), .QN(n4470) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[20]  ( .D(n3054), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][20] ), .QN(n4502) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[20]  ( .D(n3049), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][20] ), .QN(
        n4662) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[20]  ( .D(n3048), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][20] ), .QN(
        n4694) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[20]  ( .D(n3045), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][20] ), .QN(
        n4790) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[20]  ( .D(n3044), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][20] ), .QN(
        n4822) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[20]  ( .D(n3041), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][20] ), .QN(
        n4918) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[20]  ( .D(n3040), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][20] ), .QN(
        n4950) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[20]  ( .D(n3038), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][20] ), .QN(
        n5014) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[20]  ( .D(n3037), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][20] ), .QN(
        n5046) );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[20]  ( .D(n3025), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[20] ), .QN(
        n5565) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[20]  ( .D(n3024), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[52] ), .QN(
        n5610) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[20]  ( .D(n3023), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[20] ), .QN(
        \UUT/Mpath/the_alu/N44 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[20]  ( .D(n3022), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [20]), .QN(
        n2648) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[20]  ( .D(n3021), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [20])
         );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[21]  ( .D(n3015), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][21] ), .QN(n4469) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[21]  ( .D(n3014), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][21] ), .QN(n4501) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[21]  ( .D(n3009), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][21] ), .QN(
        n4661) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[21]  ( .D(n3008), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][21] ), .QN(
        n4693) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[21]  ( .D(n3005), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][21] ), .QN(
        n4789) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[21]  ( .D(n3004), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][21] ), .QN(
        n4821) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[21]  ( .D(n3001), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][21] ), .QN(
        n4917) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[21]  ( .D(n3000), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][21] ), .QN(
        n4949) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[21]  ( .D(n2998), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][21] ), .QN(
        n5013) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[21]  ( .D(n2997), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][21] ), .QN(
        n5045) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[21]  ( .D(n2988), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[21] ), .QN(
        \UUT/Mpath/the_alu/N41 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[21]  ( .D(n2987), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[21] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[21]  ( .D(n2985), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[21] ), .QN(
        n5563) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[21]  ( .D(n2984), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[53] ), .QN(
        n5609) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[21]  ( .D(n2983), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[21] ), .QN(
        \UUT/Mpath/the_alu/N42 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[21]  ( .D(n2982), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [21]), .QN(
        n2645) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[22]  ( .D(n2975), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][22] ), .QN(n4468) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[22]  ( .D(n2974), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][22] ), .QN(n4500) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[22]  ( .D(n2969), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][22] ), .QN(
        n4660) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[22]  ( .D(n2968), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][22] ), .QN(
        n4692) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[22]  ( .D(n2965), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][22] ), .QN(
        n4788) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[22]  ( .D(n2964), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][22] ), .QN(
        n4820) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[22]  ( .D(n2961), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][22] ), .QN(
        n4916) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[22]  ( .D(n2960), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][22] ), .QN(
        n4948) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[22]  ( .D(n2958), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][22] ), .QN(
        n5012) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[22]  ( .D(n2957), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][22] ), .QN(
        n5044) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[22]  ( .D(n2948), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[22] ), .QN(
        \UUT/Mpath/the_alu/N39 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[22]  ( .D(n2947), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[22] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[22]  ( .D(n2945), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[22] ), .QN(
        n5561) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[22]  ( .D(n2944), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[54] ), .QN(
        n5608) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[22]  ( .D(n2943), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[22] ), .QN(
        \UUT/Mpath/the_alu/N40 ) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[22]  ( .D(n2942), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [22]), .QN(
        n2642) );
  DFFR_X1 \UUT/regfile/rx_5/data_out_reg[24]  ( .D(n2935), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[5][24] ), .QN(n4466) );
  DFFR_X1 \UUT/regfile/rx_4/data_out_reg[24]  ( .D(n2934), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[4][24] ), .QN(n4498) );
  DFFR_X1 \UUT/regfile/rx_29/data_out_reg[24]  ( .D(n2929), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[29][24] ), .QN(
        n4658) );
  DFFR_X1 \UUT/regfile/rx_28/data_out_reg[24]  ( .D(n2928), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[28][24] ), .QN(
        n4690) );
  DFFR_X1 \UUT/regfile/rx_25/data_out_reg[24]  ( .D(n2925), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[25][24] ), .QN(
        n4786) );
  DFFR_X1 \UUT/regfile/rx_24/data_out_reg[24]  ( .D(n2924), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[24][24] ), .QN(
        n4818) );
  DFFR_X1 \UUT/regfile/rx_21/data_out_reg[24]  ( .D(n2921), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[21][24] ), .QN(
        n4914) );
  DFFR_X1 \UUT/regfile/rx_20/data_out_reg[24]  ( .D(n2920), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[20][24] ), .QN(
        n4946) );
  DFFR_X1 \UUT/regfile/rx_19/data_out_reg[24]  ( .D(n2918), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[19][24] ), .QN(
        n5010) );
  DFFR_X1 \UUT/regfile/rx_18/data_out_reg[24]  ( .D(n2917), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/regfile/reg_out[18][24] ), .QN(
        n5042) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[24]  ( .D(n2908), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[24] ), .QN(
        \UUT/Mpath/the_alu/N35 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[24]  ( .D(n2907), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[24] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[24]  ( .D(n2905), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[24] ), .QN(
        n5557) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[24]  ( .D(n2904), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[56] ), .QN(
        n5606) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[24]  ( .D(n2903), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[24] ), .QN(
        \UUT/Mpath/the_alu/N36 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[24]  ( .D(n2902), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [24])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[25]  ( .D(n2901), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[25] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[25]  ( .D(n2899), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[25] ), .QN(
        n5555) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[25]  ( .D(n2898), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[57] ), .QN(
        n5605) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[25]  ( .D(n2897), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[25] ), .QN(
        \UUT/Mpath/the_alu/N34 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[26]  ( .D(n2895), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[26] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[26]  ( .D(n2893), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[26] ), .QN(
        n5553) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[26]  ( .D(n2892), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[58] ), .QN(
        n5604) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[26]  ( .D(n2891), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[26] ), .QN(
        \UUT/Mpath/the_alu/N32 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[26]  ( .D(n2890), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [26])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[27]  ( .D(n2889), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[27] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[27]  ( .D(n2887), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[27] ), .QN(
        n5551) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[27]  ( .D(n2886), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[59] ), .QN(
        n5603) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[27]  ( .D(n2885), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[27] ), .QN(
        \UUT/Mpath/the_alu/N30 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[28]  ( .D(n2883), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[28] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[28]  ( .D(n2881), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[28] ), .QN(
        n5549) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[28]  ( .D(n2880), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[60] ), .QN(
        n5602) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[28]  ( .D(n2879), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[28] ), .QN(
        \UUT/Mpath/the_alu/N28 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[28]  ( .D(n2878), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [28])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[29]  ( .D(n2877), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[29] )
         );
  DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[29]  ( .D(n2875), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[29] ), .QN(
        n5547) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[29]  ( .D(n2874), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[29] ), .QN(
        \UUT/Mpath/the_alu/N26 ) );
  DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[31]  ( .D(n2872), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[63] ), .QN(
        n5598) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[0]  ( .D(n2867), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [0])
         );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[30]  ( .D(n2866), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[30] ), 
        .QN(n2624) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[29]  ( .D(n2865), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[29] ), 
        .QN(n2623) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[28]  ( .D(n2864), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[28] ), 
        .QN(n2622) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[27]  ( .D(n2863), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[27] ), 
        .QN(n2621) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[26]  ( .D(n2862), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[26] ), 
        .QN(n2620) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[25]  ( .D(n2861), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[25] ), 
        .QN(n2619) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[24]  ( .D(n2860), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[24] ), 
        .QN(n2618) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[23]  ( .D(n2859), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[23] ), 
        .QN(n2617) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[22]  ( .D(n2858), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[22] ), 
        .QN(n2616) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[21]  ( .D(n2857), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[21] ), 
        .QN(n2615) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[20]  ( .D(n2856), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[20] ), 
        .QN(n2614) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[19]  ( .D(n2855), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[19] ), 
        .QN(n2613) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[18]  ( .D(n2854), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[18] ), 
        .QN(n2612) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[17]  ( .D(n2853), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[17] ), 
        .QN(n2611) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[16]  ( .D(n2852), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_memhandle/smdr_out[16] ), 
        .QN(n2610) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[7]  ( .D(n2843), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[7]), .QN(n6293) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[6]  ( .D(n2842), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[6]), .QN(n6297) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[5]  ( .D(n2841), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[5]), .QN(n6300) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[4]  ( .D(n2840), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[4]), .QN(n6303) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[3]  ( .D(n2839), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[3]), .QN(n6306) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[2]  ( .D(n2838), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[2]), .QN(n6309) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[1]  ( .D(n2837), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[1]), .QN(n6285) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[0]  ( .D(n2836), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(D_DATA_OUTBUS[0]), .QN(n6289) );
  OAI22_X1 U3 ( .A1(n6289), .A2(n46), .B1(n47), .B2(n48), .ZN(n2836) );
  OAI22_X1 U4 ( .A1(n6285), .A2(n46), .B1(n49), .B2(n48), .ZN(n2837) );
  OAI22_X1 U5 ( .A1(n6309), .A2(n46), .B1(n50), .B2(n48), .ZN(n2838) );
  OAI22_X1 U6 ( .A1(n6306), .A2(n46), .B1(n51), .B2(n48), .ZN(n2839) );
  OAI22_X1 U7 ( .A1(n6303), .A2(n46), .B1(n52), .B2(n48), .ZN(n2840) );
  OAI22_X1 U8 ( .A1(n6300), .A2(n46), .B1(n53), .B2(n48), .ZN(n2841) );
  OAI22_X1 U9 ( .A1(n6297), .A2(n46), .B1(n54), .B2(n48), .ZN(n2842) );
  OAI22_X1 U10 ( .A1(n6293), .A2(n46), .B1(n55), .B2(n48), .ZN(n2843) );
  OAI22_X1 U11 ( .A1(n6290), .A2(n46), .B1(n56), .B2(n48), .ZN(n2844) );
  OAI22_X1 U12 ( .A1(n6288), .A2(n46), .B1(n57), .B2(n48), .ZN(n2845) );
  OAI22_X1 U13 ( .A1(n6308), .A2(n46), .B1(n58), .B2(n48), .ZN(n2846) );
  OAI22_X1 U14 ( .A1(n6305), .A2(n46), .B1(n59), .B2(n48), .ZN(n2847) );
  OAI22_X1 U15 ( .A1(n6302), .A2(n46), .B1(n60), .B2(n48), .ZN(n2848) );
  OAI22_X1 U16 ( .A1(n6299), .A2(n46), .B1(n61), .B2(n48), .ZN(n2849) );
  OAI22_X1 U38 ( .A1(n6296), .A2(n46), .B1(n62), .B2(n48), .ZN(n2850) );
  OAI22_X1 U39 ( .A1(n6292), .A2(n46), .B1(n63), .B2(n48), .ZN(n2851) );
  OAI22_X1 U40 ( .A1(n46), .A2(n2610), .B1(n64), .B2(n48), .ZN(n2852) );
  OAI22_X1 U41 ( .A1(n46), .A2(n2611), .B1(n65), .B2(n48), .ZN(n2853) );
  OAI22_X1 U42 ( .A1(n46), .A2(n2612), .B1(n66), .B2(n48), .ZN(n2854) );
  OAI22_X1 U43 ( .A1(n46), .A2(n2613), .B1(n67), .B2(n48), .ZN(n2855) );
  OAI22_X1 U44 ( .A1(n46), .A2(n2614), .B1(n68), .B2(n48), .ZN(n2856) );
  OAI22_X1 U45 ( .A1(n46), .A2(n2615), .B1(n69), .B2(n48), .ZN(n2857) );
  OAI22_X1 U46 ( .A1(n46), .A2(n2616), .B1(n70), .B2(n48), .ZN(n2858) );
  OAI22_X1 U47 ( .A1(n46), .A2(n2617), .B1(n71), .B2(n48), .ZN(n2859) );
  OAI22_X1 U48 ( .A1(n46), .A2(n2618), .B1(n72), .B2(n48), .ZN(n2860) );
  OAI22_X1 U49 ( .A1(n46), .A2(n2619), .B1(n73), .B2(n48), .ZN(n2861) );
  OAI22_X1 U50 ( .A1(n46), .A2(n2620), .B1(n74), .B2(n48), .ZN(n2862) );
  OAI22_X1 U51 ( .A1(n46), .A2(n2621), .B1(n75), .B2(n48), .ZN(n2863) );
  OAI22_X1 U52 ( .A1(n46), .A2(n2622), .B1(n76), .B2(n48), .ZN(n2864) );
  OAI22_X1 U53 ( .A1(n46), .A2(n2623), .B1(n77), .B2(n48), .ZN(n2865) );
  OAI22_X1 U54 ( .A1(n46), .A2(n2624), .B1(n78), .B2(n48), .ZN(n2866) );
  OAI221_X1 U55 ( .B1(n79), .B2(n80), .C1(n47), .C2(n81), .A(n82), .ZN(n2867)
         );
  NAND2_X1 U56 ( .A1(\UUT/Mpath/the_mult/x_operand2 [0]), .A2(n6340), .ZN(n82)
         );
  OAI221_X1 U57 ( .B1(n84), .B2(n80), .C1(n71), .C2(n81), .A(n85), .ZN(n2868)
         );
  NAND2_X1 U58 ( .A1(n7048), .A2(n6340), .ZN(n85) );
  NAND2_X1 U60 ( .A1(\UUT/Mpath/the_mult/x_operand2 [31]), .A2(n6340), .ZN(n88) );
  OAI211_X1 U61 ( .C1(n5902), .C2(n89), .A(n90), .B(n91), .ZN(n2870) );
  OAI221_X1 U63 ( .B1(n78), .B2(n94), .C1(\UUT/Mpath/the_alu/N24 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n95), .ZN(n2871) );
  AOI21_X1 U64 ( .B1(n96), .B2(\UUT/Mcontrol/d_sampled_finstr [14]), .A(n97), 
        .ZN(n95) );
  INV_X1 U65 ( .A(n6840), .ZN(n78) );
  OAI221_X1 U67 ( .B1(n103), .B2(n104), .C1(n5598), .C2(n105), .A(n106), .ZN(
        n2872) );
  OAI211_X1 U69 ( .C1(n5903), .C2(n89), .A(n90), .B(n110), .ZN(n2873) );
  AOI22_X1 U70 ( .A1(n92), .A2(n111), .B1(\UUT/Mpath/the_mult/x_operand2 [29]), 
        .B2(n6340), .ZN(n110) );
  OAI221_X1 U71 ( .B1(n77), .B2(n94), .C1(\UUT/Mpath/the_alu/N26 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n112), .ZN(n2874) );
  AOI21_X1 U72 ( .B1(n96), .B2(\UUT/Mcontrol/d_sampled_finstr [13]), .A(n97), 
        .ZN(n112) );
  INV_X1 U73 ( .A(n111), .ZN(n77) );
  OAI221_X1 U75 ( .B1(n115), .B2(n116), .C1(n5547), .C2(n117), .A(n118), .ZN(
        n2875) );
  AOI22_X1 U76 ( .A1(n119), .A2(n120), .B1(\UUT/Mpath/the_mult/Mad_out [29]), 
        .B2(n121), .ZN(n118) );
  OAI22_X1 U77 ( .A1(n7383), .A2(n123), .B1(n5548), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2876) );
  OAI221_X1 U78 ( .B1(n5318), .B2(n6350), .C1(n125), .C2(n123), .A(n126), .ZN(
        n2877) );
  AOI22_X1 U79 ( .A1(n127), .A2(n128), .B1(n129), .B2(n130), .ZN(n126) );
  INV_X1 U80 ( .A(\UUT/Mpath/the_mult/x_operand1[29] ), .ZN(n123) );
  OAI211_X1 U81 ( .C1(n5905), .C2(n89), .A(n90), .B(n131), .ZN(n2878) );
  AOI22_X1 U82 ( .A1(n92), .A2(n132), .B1(\UUT/Mpath/the_mult/x_operand2 [28]), 
        .B2(n6340), .ZN(n131) );
  OAI221_X1 U83 ( .B1(n76), .B2(n94), .C1(\UUT/Mpath/the_alu/N28 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n133), .ZN(n2879) );
  AOI21_X1 U84 ( .B1(n96), .B2(\UUT/Mcontrol/d_sampled_finstr [12]), .A(n97), 
        .ZN(n133) );
  INV_X1 U85 ( .A(n132), .ZN(n76) );
  OAI222_X1 U86 ( .A1(n134), .A2(n5332), .B1(n135), .B2(n101), .C1(n5368), 
        .C2(n102), .ZN(n132) );
  OAI221_X1 U87 ( .B1(n103), .B2(n136), .C1(n5602), .C2(n105), .A(n137), .ZN(
        n2880) );
  AOI22_X1 U88 ( .A1(n107), .A2(n138), .B1(\UUT/Mpath/the_mult/Mad_out [60]), 
        .B2(n109), .ZN(n137) );
  OAI221_X1 U89 ( .B1(n115), .B2(n139), .C1(n5549), .C2(n117), .A(n140), .ZN(
        n2881) );
  AOI22_X1 U90 ( .A1(n119), .A2(n138), .B1(\UUT/Mpath/the_mult/Mad_out [28]), 
        .B2(n121), .ZN(n140) );
  OAI22_X1 U92 ( .A1(n7387), .A2(n141), .B1(n5550), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2882) );
  OAI221_X1 U93 ( .B1(n5319), .B2(n6350), .C1(n125), .C2(n141), .A(n142), .ZN(
        n2883) );
  AOI22_X1 U94 ( .A1(n127), .A2(n143), .B1(n129), .B2(n144), .ZN(n142) );
  INV_X1 U95 ( .A(\UUT/Mpath/the_mult/x_operand1[28] ), .ZN(n141) );
  OAI211_X1 U96 ( .C1(n5906), .C2(n89), .A(n90), .B(n145), .ZN(n2884) );
  AOI22_X1 U97 ( .A1(n92), .A2(n146), .B1(n6973), .B2(n6340), .ZN(n145) );
  NAND2_X1 U98 ( .A1(n125), .A2(n147), .ZN(n90) );
  OAI221_X1 U99 ( .B1(n75), .B2(n94), .C1(\UUT/Mpath/the_alu/N30 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n148), .ZN(n2885) );
  AOI21_X1 U100 ( .B1(n96), .B2(\UUT/Mcontrol/d_sampled_finstr [11]), .A(n97), 
        .ZN(n148) );
  AND2_X1 U101 ( .A1(\UUT/Mcontrol/N22 ), .A2(n147), .ZN(n97) );
  NAND2_X1 U102 ( .A1(n149), .A2(n150), .ZN(n147) );
  INV_X1 U103 ( .A(n146), .ZN(n75) );
  OAI222_X1 U104 ( .A1(n151), .A2(n99), .B1(n152), .B2(n101), .C1(n5371), .C2(
        n102), .ZN(n146) );
  OAI221_X1 U105 ( .B1(n103), .B2(n153), .C1(n5603), .C2(n105), .A(n154), .ZN(
        n2886) );
  AOI22_X1 U106 ( .A1(n107), .A2(n155), .B1(\UUT/Mpath/the_mult/Mad_out [59]), 
        .B2(n109), .ZN(n154) );
  OAI221_X1 U107 ( .B1(n115), .B2(n156), .C1(n5551), .C2(n117), .A(n157), .ZN(
        n2887) );
  AOI22_X1 U108 ( .A1(n119), .A2(n155), .B1(\UUT/Mpath/the_mult/Mad_out [27]), 
        .B2(n121), .ZN(n157) );
  OAI22_X1 U110 ( .A1(n7388), .A2(n158), .B1(n5552), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2888) );
  OAI221_X1 U111 ( .B1(n5320), .B2(n6350), .C1(n125), .C2(n158), .A(n159), 
        .ZN(n2889) );
  AOI22_X1 U112 ( .A1(n127), .A2(n160), .B1(n129), .B2(n161), .ZN(n159) );
  INV_X1 U113 ( .A(\UUT/Mpath/the_mult/x_operand1[27] ), .ZN(n158) );
  OAI221_X1 U114 ( .B1(n162), .B2(n6340), .C1(n5762), .C2(n89), .A(n163), .ZN(
        n2890) );
  AOI22_X1 U115 ( .A1(n92), .A2(n164), .B1(\UUT/Mpath/the_mult/x_operand2 [26]), .B2(n6340), .ZN(n163) );
  INV_X1 U116 ( .A(n165), .ZN(n162) );
  OAI221_X1 U117 ( .B1(n74), .B2(n94), .C1(\UUT/Mpath/the_alu/N32 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n166), .ZN(n2891) );
  AOI22_X1 U118 ( .A1(\UUT/Mcontrol/N22 ), .A2(n165), .B1(n96), .B2(
        \UUT/Mcontrol/d_sampled_finstr [10]), .ZN(n166) );
  OAI21_X1 U119 ( .B1(n5760), .B2(n167), .A(n149), .ZN(n165) );
  INV_X1 U120 ( .A(n164), .ZN(n74) );
  OAI222_X1 U121 ( .A1(n168), .A2(n5332), .B1(n169), .B2(n101), .C1(n5374), 
        .C2(n102), .ZN(n164) );
  OAI221_X1 U122 ( .B1(n103), .B2(n170), .C1(n5604), .C2(n105), .A(n171), .ZN(
        n2892) );
  AOI22_X1 U123 ( .A1(n107), .A2(n172), .B1(\UUT/Mpath/the_mult/Mad_out [58]), 
        .B2(n109), .ZN(n171) );
  OAI221_X1 U124 ( .B1(n115), .B2(n173), .C1(n5553), .C2(n117), .A(n174), .ZN(
        n2893) );
  AOI22_X1 U125 ( .A1(n119), .A2(n172), .B1(\UUT/Mpath/the_mult/Mad_out [26]), 
        .B2(n121), .ZN(n174) );
  OAI22_X1 U127 ( .A1(n7388), .A2(n175), .B1(n5554), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2894) );
  OAI221_X1 U128 ( .B1(n5321), .B2(n6350), .C1(n125), .C2(n175), .A(n176), 
        .ZN(n2895) );
  AOI22_X1 U129 ( .A1(n127), .A2(n177), .B1(n129), .B2(n178), .ZN(n176) );
  INV_X1 U130 ( .A(\UUT/Mpath/the_mult/x_operand1[26] ), .ZN(n175) );
  OAI221_X1 U131 ( .B1(n179), .B2(n6340), .C1(n5769), .C2(n89), .A(n180), .ZN(
        n2896) );
  AOI22_X1 U132 ( .A1(n92), .A2(n181), .B1(n6963), .B2(n6340), .ZN(n180) );
  INV_X1 U133 ( .A(n182), .ZN(n179) );
  OAI221_X1 U134 ( .B1(n73), .B2(n94), .C1(\UUT/Mpath/the_alu/N34 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n183), .ZN(n2897) );
  AOI22_X1 U135 ( .A1(\UUT/Mcontrol/N22 ), .A2(n182), .B1(n96), .B2(
        \UUT/Mcontrol/d_sampled_finstr [9]), .ZN(n183) );
  OAI21_X1 U136 ( .B1(n5768), .B2(n167), .A(n149), .ZN(n182) );
  INV_X1 U137 ( .A(n181), .ZN(n73) );
  OAI222_X1 U138 ( .A1(n184), .A2(n99), .B1(n185), .B2(n101), .C1(n5377), .C2(
        n102), .ZN(n181) );
  OAI221_X1 U139 ( .B1(n103), .B2(n186), .C1(n5605), .C2(n105), .A(n187), .ZN(
        n2898) );
  AOI22_X1 U140 ( .A1(n107), .A2(n188), .B1(\UUT/Mpath/the_mult/Mad_out [57]), 
        .B2(n109), .ZN(n187) );
  OAI221_X1 U141 ( .B1(n115), .B2(n189), .C1(n5555), .C2(n117), .A(n190), .ZN(
        n2899) );
  AOI22_X1 U142 ( .A1(n119), .A2(n188), .B1(\UUT/Mpath/the_mult/Mad_out [25]), 
        .B2(n121), .ZN(n190) );
  OAI22_X1 U144 ( .A1(n7388), .A2(n191), .B1(n5556), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2900) );
  OAI221_X1 U145 ( .B1(n5322), .B2(n6350), .C1(n125), .C2(n191), .A(n192), 
        .ZN(n2901) );
  AOI22_X1 U146 ( .A1(n127), .A2(n193), .B1(n129), .B2(n194), .ZN(n192) );
  INV_X1 U147 ( .A(\UUT/Mpath/the_mult/x_operand1[25] ), .ZN(n191) );
  OAI221_X1 U148 ( .B1(n195), .B2(n6340), .C1(n5776), .C2(n89), .A(n196), .ZN(
        n2902) );
  AOI22_X1 U149 ( .A1(n197), .A2(n92), .B1(\UUT/Mpath/the_mult/x_operand2 [24]), .B2(n6340), .ZN(n196) );
  INV_X1 U150 ( .A(n81), .ZN(n92) );
  NAND3_X1 U151 ( .A1(n7096), .A2(n125), .A3(n198), .ZN(n89) );
  INV_X1 U152 ( .A(n199), .ZN(n195) );
  OAI221_X1 U153 ( .B1(n72), .B2(n94), .C1(\UUT/Mpath/the_alu/N36 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n200), .ZN(n2903) );
  AOI22_X1 U154 ( .A1(\UUT/Mcontrol/N22 ), .A2(n199), .B1(n96), .B2(
        \UUT/Mcontrol/d_sampled_finstr [8]), .ZN(n200) );
  OAI21_X1 U155 ( .B1(n5775), .B2(n167), .A(n149), .ZN(n199) );
  INV_X1 U156 ( .A(n201), .ZN(n149) );
  OAI21_X1 U157 ( .B1(n202), .B2(n203), .A(n204), .ZN(n201) );
  NAND2_X1 U158 ( .A1(n205), .A2(n206), .ZN(n167) );
  INV_X1 U159 ( .A(n5754), .ZN(n206) );
  INV_X1 U160 ( .A(n197), .ZN(n72) );
  OAI222_X1 U161 ( .A1(n207), .A2(n99), .B1(n208), .B2(n101), .C1(n5380), .C2(
        n102), .ZN(n197) );
  OAI221_X1 U162 ( .B1(n103), .B2(n209), .C1(n5606), .C2(n105), .A(n210), .ZN(
        n2904) );
  AOI22_X1 U163 ( .A1(n107), .A2(n211), .B1(\UUT/Mpath/the_mult/Mad_out [56]), 
        .B2(n109), .ZN(n210) );
  OAI221_X1 U164 ( .B1(n115), .B2(n212), .C1(n5557), .C2(n117), .A(n213), .ZN(
        n2905) );
  AOI22_X1 U165 ( .A1(n119), .A2(n211), .B1(\UUT/Mpath/the_mult/Mad_out [24]), 
        .B2(n121), .ZN(n213) );
  OAI22_X1 U167 ( .A1(n7388), .A2(n214), .B1(n5558), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2906) );
  OAI221_X1 U168 ( .B1(n5323), .B2(n6350), .C1(n125), .C2(n214), .A(n215), 
        .ZN(n2907) );
  AOI22_X1 U169 ( .A1(n127), .A2(n216), .B1(n129), .B2(n217), .ZN(n215) );
  INV_X1 U170 ( .A(\UUT/Mpath/the_mult/x_operand1[24] ), .ZN(n214) );
  OAI221_X1 U171 ( .B1(n5323), .B2(n218), .C1(\UUT/Mpath/the_alu/N35 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n219), .ZN(n2908) );
  AOI22_X1 U172 ( .A1(n220), .A2(n216), .B1(n221), .B2(n217), .ZN(n219) );
  OAI22_X1 U173 ( .A1(n5298), .A2(n6393), .B1(n208), .B2(n223), .ZN(n2909) );
  OAI22_X1 U174 ( .A1(n5266), .A2(n6396), .B1(n208), .B2(n225), .ZN(n2910) );
  OAI22_X1 U175 ( .A1(n5234), .A2(n6387), .B1(n208), .B2(n227), .ZN(n2911) );
  OAI22_X1 U176 ( .A1(n5202), .A2(n6395), .B1(n208), .B2(n229), .ZN(n2912) );
  OAI22_X1 U177 ( .A1(n5170), .A2(n6390), .B1(n208), .B2(n231), .ZN(n2913) );
  OAI22_X1 U178 ( .A1(n5138), .A2(n6385), .B1(n208), .B2(n233), .ZN(n2914) );
  OAI22_X1 U179 ( .A1(n5106), .A2(n6389), .B1(n208), .B2(n235), .ZN(n2915) );
  OAI22_X1 U180 ( .A1(n5074), .A2(n6382), .B1(n208), .B2(n237), .ZN(n2916) );
  OAI22_X1 U181 ( .A1(n5042), .A2(n6380), .B1(n208), .B2(n239), .ZN(n2917) );
  OAI22_X1 U182 ( .A1(n5010), .A2(n6379), .B1(n208), .B2(n241), .ZN(n2918) );
  OAI22_X1 U183 ( .A1(n4978), .A2(n6376), .B1(n208), .B2(n243), .ZN(n2919) );
  OAI22_X1 U184 ( .A1(n4946), .A2(n6375), .B1(n208), .B2(n245), .ZN(n2920) );
  OAI22_X1 U185 ( .A1(n4914), .A2(n6372), .B1(n208), .B2(n247), .ZN(n2921) );
  OAI22_X1 U186 ( .A1(n4882), .A2(n6371), .B1(n208), .B2(n249), .ZN(n2922) );
  OAI22_X1 U187 ( .A1(n4850), .A2(n6368), .B1(n208), .B2(n251), .ZN(n2923) );
  OAI22_X1 U188 ( .A1(n4818), .A2(n6367), .B1(n208), .B2(n253), .ZN(n2924) );
  OAI22_X1 U189 ( .A1(n4786), .A2(n6364), .B1(n208), .B2(n255), .ZN(n2925) );
  OAI22_X1 U190 ( .A1(n4754), .A2(n6362), .B1(n208), .B2(n257), .ZN(n2926) );
  OAI22_X1 U191 ( .A1(n4722), .A2(n6361), .B1(n208), .B2(n259), .ZN(n2927) );
  OAI22_X1 U192 ( .A1(n4690), .A2(n6365), .B1(n208), .B2(n261), .ZN(n2928) );
  OAI22_X1 U193 ( .A1(n4658), .A2(n6366), .B1(n208), .B2(n263), .ZN(n2929) );
  OAI22_X1 U194 ( .A1(n4626), .A2(n6369), .B1(n208), .B2(n265), .ZN(n2930) );
  OAI22_X1 U195 ( .A1(n4594), .A2(n6370), .B1(n208), .B2(n267), .ZN(n2931) );
  OAI22_X1 U196 ( .A1(n4562), .A2(n6373), .B1(n208), .B2(n269), .ZN(n2932) );
  OAI22_X1 U197 ( .A1(n4530), .A2(n6374), .B1(n208), .B2(n271), .ZN(n2933) );
  OAI22_X1 U198 ( .A1(n4498), .A2(n6377), .B1(n208), .B2(n273), .ZN(n2934) );
  OAI22_X1 U199 ( .A1(n4466), .A2(n6378), .B1(n208), .B2(n275), .ZN(n2935) );
  OAI22_X1 U200 ( .A1(n4434), .A2(n6381), .B1(n208), .B2(n277), .ZN(n2936) );
  OAI22_X1 U201 ( .A1(n4402), .A2(n6384), .B1(n208), .B2(n279), .ZN(n2937) );
  OAI22_X1 U202 ( .A1(n4370), .A2(n6383), .B1(n208), .B2(n281), .ZN(n2938) );
  OAI22_X1 U203 ( .A1(n4338), .A2(n6391), .B1(n208), .B2(n283), .ZN(n2939) );
  OAI221_X1 U205 ( .B1(n5870), .B2(n284), .C1(n5623), .C2(n5381), .A(n285), 
        .ZN(n216) );
  OAI22_X1 U206 ( .A1(n5381), .A2(\UUT/Mcontrol/N22 ), .B1(n207), .B2(n7397), 
        .ZN(n2940) );
  INV_X1 U210 ( .A(n5606), .ZN(n292) );
  INV_X1 U211 ( .A(n5557), .ZN(n290) );
  OAI221_X1 U212 ( .B1(n294), .B2(n80), .C1(n70), .C2(n81), .A(n295), .ZN(
        n2941) );
  NAND2_X1 U213 ( .A1(\UUT/Mpath/the_mult/x_operand2 [22]), .A2(n6340), .ZN(
        n295) );
  OAI222_X1 U216 ( .A1(n70), .A2(n94), .B1(n294), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N40 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n2943) );
  INV_X1 U217 ( .A(n303), .ZN(n70) );
  OAI222_X1 U218 ( .A1(n304), .A2(n99), .B1(n305), .B2(n101), .C1(n5386), .C2(
        n102), .ZN(n303) );
  OAI221_X1 U219 ( .B1(n103), .B2(n306), .C1(n5608), .C2(n105), .A(n307), .ZN(
        n2944) );
  AOI22_X1 U220 ( .A1(n107), .A2(n308), .B1(\UUT/Mpath/the_mult/Mad_out [54]), 
        .B2(n109), .ZN(n307) );
  OAI221_X1 U221 ( .B1(n115), .B2(n309), .C1(n5561), .C2(n117), .A(n310), .ZN(
        n2945) );
  AOI22_X1 U222 ( .A1(n119), .A2(n308), .B1(\UUT/Mpath/the_mult/Mad_out [22]), 
        .B2(n121), .ZN(n310) );
  OAI22_X1 U224 ( .A1(n7387), .A2(n311), .B1(n5562), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2946) );
  OAI221_X1 U225 ( .B1(n312), .B2(n6350), .C1(n125), .C2(n311), .A(n313), .ZN(
        n2947) );
  AOI22_X1 U226 ( .A1(n127), .A2(n314), .B1(n129), .B2(n315), .ZN(n313) );
  INV_X1 U227 ( .A(\UUT/Mpath/the_mult/x_operand1[22] ), .ZN(n311) );
  OAI221_X1 U228 ( .B1(n312), .B2(n218), .C1(\UUT/Mpath/the_alu/N39 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n316), .ZN(n2948) );
  AOI22_X1 U229 ( .A1(n220), .A2(n314), .B1(n221), .B2(n315), .ZN(n316) );
  OAI22_X1 U230 ( .A1(n5300), .A2(n6393), .B1(n305), .B2(n223), .ZN(n2949) );
  OAI22_X1 U231 ( .A1(n5268), .A2(n6396), .B1(n305), .B2(n225), .ZN(n2950) );
  OAI22_X1 U232 ( .A1(n5236), .A2(n6387), .B1(n305), .B2(n227), .ZN(n2951) );
  OAI22_X1 U233 ( .A1(n5204), .A2(n6395), .B1(n305), .B2(n229), .ZN(n2952) );
  OAI22_X1 U234 ( .A1(n5172), .A2(n6390), .B1(n305), .B2(n231), .ZN(n2953) );
  OAI22_X1 U235 ( .A1(n5140), .A2(n6385), .B1(n305), .B2(n233), .ZN(n2954) );
  OAI22_X1 U236 ( .A1(n5108), .A2(n6389), .B1(n305), .B2(n235), .ZN(n2955) );
  OAI22_X1 U237 ( .A1(n5076), .A2(n6382), .B1(n305), .B2(n237), .ZN(n2956) );
  OAI22_X1 U238 ( .A1(n5044), .A2(n6380), .B1(n305), .B2(n239), .ZN(n2957) );
  OAI22_X1 U239 ( .A1(n5012), .A2(n6379), .B1(n305), .B2(n241), .ZN(n2958) );
  OAI22_X1 U240 ( .A1(n4980), .A2(n6376), .B1(n305), .B2(n243), .ZN(n2959) );
  OAI22_X1 U241 ( .A1(n4948), .A2(n6375), .B1(n305), .B2(n245), .ZN(n2960) );
  OAI22_X1 U242 ( .A1(n4916), .A2(n6372), .B1(n305), .B2(n247), .ZN(n2961) );
  OAI22_X1 U243 ( .A1(n4884), .A2(n6371), .B1(n305), .B2(n249), .ZN(n2962) );
  OAI22_X1 U244 ( .A1(n4852), .A2(n6368), .B1(n305), .B2(n251), .ZN(n2963) );
  OAI22_X1 U245 ( .A1(n4820), .A2(n6367), .B1(n305), .B2(n253), .ZN(n2964) );
  OAI22_X1 U246 ( .A1(n4788), .A2(n6364), .B1(n305), .B2(n255), .ZN(n2965) );
  OAI22_X1 U247 ( .A1(n4756), .A2(n6362), .B1(n305), .B2(n257), .ZN(n2966) );
  OAI22_X1 U248 ( .A1(n4724), .A2(n6361), .B1(n305), .B2(n259), .ZN(n2967) );
  OAI22_X1 U249 ( .A1(n4692), .A2(n6365), .B1(n305), .B2(n261), .ZN(n2968) );
  OAI22_X1 U250 ( .A1(n4660), .A2(n6366), .B1(n305), .B2(n263), .ZN(n2969) );
  OAI22_X1 U251 ( .A1(n4628), .A2(n6369), .B1(n305), .B2(n265), .ZN(n2970) );
  OAI22_X1 U252 ( .A1(n4596), .A2(n6370), .B1(n305), .B2(n267), .ZN(n2971) );
  OAI22_X1 U253 ( .A1(n4564), .A2(n6373), .B1(n305), .B2(n269), .ZN(n2972) );
  OAI22_X1 U254 ( .A1(n4532), .A2(n6374), .B1(n305), .B2(n271), .ZN(n2973) );
  OAI22_X1 U255 ( .A1(n4500), .A2(n6377), .B1(n305), .B2(n273), .ZN(n2974) );
  OAI22_X1 U256 ( .A1(n4468), .A2(n6378), .B1(n305), .B2(n275), .ZN(n2975) );
  OAI22_X1 U257 ( .A1(n4436), .A2(n6381), .B1(n305), .B2(n277), .ZN(n2976) );
  OAI22_X1 U258 ( .A1(n4404), .A2(n6384), .B1(n305), .B2(n279), .ZN(n2977) );
  OAI22_X1 U259 ( .A1(n4372), .A2(n6383), .B1(n305), .B2(n281), .ZN(n2978) );
  OAI22_X1 U260 ( .A1(n4340), .A2(n6391), .B1(n305), .B2(n283), .ZN(n2979) );
  OAI221_X1 U262 ( .B1(n317), .B2(n284), .C1(n5623), .C2(n5387), .A(n285), 
        .ZN(n314) );
  INV_X1 U263 ( .A(D_DATA_INBUS[22]), .ZN(n317) );
  OAI22_X1 U264 ( .A1(n5387), .A2(\UUT/Mcontrol/N22 ), .B1(n304), .B2(n7397), 
        .ZN(n2980) );
  INV_X1 U265 ( .A(n315), .ZN(n304) );
  OAI211_X1 U266 ( .C1(n5980), .C2(n287), .A(n318), .B(n319), .ZN(n315) );
  AOI222_X1 U267 ( .A1(\UUT/Mpath/the_mult/x_mult_out[22] ), .A2(n6357), .B1(
        n320), .B2(n321), .C1(n291), .C2(n322), .ZN(n319) );
  INV_X1 U268 ( .A(n5608), .ZN(n322) );
  AOI22_X1 U270 ( .A1(n6397), .A2(n323), .B1(n324), .B2(n6115), .ZN(n318) );
  INV_X1 U271 ( .A(n5561), .ZN(n323) );
  OAI221_X1 U272 ( .B1(n325), .B2(n80), .C1(n69), .C2(n81), .A(n326), .ZN(
        n2981) );
  NAND2_X1 U273 ( .A1(n7053), .A2(n6340), .ZN(n326) );
  OAI222_X1 U276 ( .A1(n69), .A2(n94), .B1(n325), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N42 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n2983) );
  INV_X1 U277 ( .A(n328), .ZN(n69) );
  OAI222_X1 U278 ( .A1(n329), .A2(n99), .B1(n330), .B2(n101), .C1(n5389), .C2(
        n102), .ZN(n328) );
  OAI221_X1 U279 ( .B1(n103), .B2(n331), .C1(n5609), .C2(n105), .A(n332), .ZN(
        n2984) );
  AOI22_X1 U280 ( .A1(n107), .A2(n333), .B1(\UUT/Mpath/the_mult/Mad_out [53]), 
        .B2(n109), .ZN(n332) );
  OAI221_X1 U281 ( .B1(n115), .B2(n334), .C1(n5563), .C2(n117), .A(n335), .ZN(
        n2985) );
  AOI22_X1 U282 ( .A1(n119), .A2(n333), .B1(\UUT/Mpath/the_mult/Mad_out [21]), 
        .B2(n121), .ZN(n335) );
  OAI22_X1 U284 ( .A1(n7387), .A2(n336), .B1(n5564), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n2986) );
  OAI221_X1 U285 ( .B1(n337), .B2(n124), .C1(n125), .C2(n336), .A(n338), .ZN(
        n2987) );
  AOI22_X1 U286 ( .A1(n127), .A2(n339), .B1(n129), .B2(n340), .ZN(n338) );
  INV_X1 U287 ( .A(\UUT/Mpath/the_mult/x_operand1[21] ), .ZN(n336) );
  OAI221_X1 U288 ( .B1(n337), .B2(n218), .C1(\UUT/Mpath/the_alu/N41 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n341), .ZN(n2988) );
  AOI22_X1 U289 ( .A1(n220), .A2(n339), .B1(n221), .B2(n340), .ZN(n341) );
  OAI22_X1 U290 ( .A1(n5301), .A2(n6393), .B1(n330), .B2(n223), .ZN(n2989) );
  OAI22_X1 U291 ( .A1(n5269), .A2(n224), .B1(n330), .B2(n225), .ZN(n2990) );
  OAI22_X1 U292 ( .A1(n5237), .A2(n6387), .B1(n330), .B2(n227), .ZN(n2991) );
  OAI22_X1 U293 ( .A1(n5205), .A2(n6395), .B1(n330), .B2(n229), .ZN(n2992) );
  OAI22_X1 U294 ( .A1(n5173), .A2(n230), .B1(n330), .B2(n231), .ZN(n2993) );
  OAI22_X1 U295 ( .A1(n5141), .A2(n232), .B1(n330), .B2(n233), .ZN(n2994) );
  OAI22_X1 U296 ( .A1(n5109), .A2(n6389), .B1(n330), .B2(n235), .ZN(n2995) );
  OAI22_X1 U297 ( .A1(n5077), .A2(n236), .B1(n330), .B2(n237), .ZN(n2996) );
  OAI22_X1 U298 ( .A1(n5045), .A2(n238), .B1(n330), .B2(n239), .ZN(n2997) );
  OAI22_X1 U299 ( .A1(n5013), .A2(n240), .B1(n330), .B2(n241), .ZN(n2998) );
  OAI22_X1 U300 ( .A1(n4981), .A2(n242), .B1(n330), .B2(n243), .ZN(n2999) );
  OAI22_X1 U301 ( .A1(n4949), .A2(n244), .B1(n330), .B2(n245), .ZN(n3000) );
  OAI22_X1 U302 ( .A1(n4917), .A2(n246), .B1(n330), .B2(n247), .ZN(n3001) );
  OAI22_X1 U303 ( .A1(n4885), .A2(n248), .B1(n330), .B2(n249), .ZN(n3002) );
  OAI22_X1 U304 ( .A1(n4853), .A2(n250), .B1(n330), .B2(n251), .ZN(n3003) );
  OAI22_X1 U305 ( .A1(n4821), .A2(n252), .B1(n330), .B2(n253), .ZN(n3004) );
  OAI22_X1 U306 ( .A1(n4789), .A2(n6364), .B1(n330), .B2(n255), .ZN(n3005) );
  OAI22_X1 U307 ( .A1(n4757), .A2(n256), .B1(n330), .B2(n257), .ZN(n3006) );
  OAI22_X1 U308 ( .A1(n4725), .A2(n6361), .B1(n330), .B2(n259), .ZN(n3007) );
  OAI22_X1 U309 ( .A1(n4693), .A2(n260), .B1(n330), .B2(n261), .ZN(n3008) );
  OAI22_X1 U310 ( .A1(n4661), .A2(n262), .B1(n330), .B2(n263), .ZN(n3009) );
  OAI22_X1 U311 ( .A1(n4629), .A2(n264), .B1(n330), .B2(n265), .ZN(n3010) );
  OAI22_X1 U312 ( .A1(n4597), .A2(n266), .B1(n330), .B2(n267), .ZN(n3011) );
  OAI22_X1 U313 ( .A1(n4565), .A2(n268), .B1(n330), .B2(n269), .ZN(n3012) );
  OAI22_X1 U314 ( .A1(n4533), .A2(n270), .B1(n330), .B2(n271), .ZN(n3013) );
  OAI22_X1 U315 ( .A1(n4501), .A2(n272), .B1(n330), .B2(n273), .ZN(n3014) );
  OAI22_X1 U316 ( .A1(n4469), .A2(n274), .B1(n330), .B2(n275), .ZN(n3015) );
  OAI22_X1 U317 ( .A1(n4437), .A2(n276), .B1(n330), .B2(n277), .ZN(n3016) );
  OAI22_X1 U318 ( .A1(n4405), .A2(n278), .B1(n330), .B2(n279), .ZN(n3017) );
  OAI22_X1 U319 ( .A1(n4373), .A2(n280), .B1(n330), .B2(n281), .ZN(n3018) );
  OAI22_X1 U320 ( .A1(n4341), .A2(n282), .B1(n330), .B2(n283), .ZN(n3019) );
  OAI221_X1 U322 ( .B1(n342), .B2(n284), .C1(n5623), .C2(n5390), .A(n285), 
        .ZN(n339) );
  INV_X1 U323 ( .A(D_DATA_INBUS[21]), .ZN(n342) );
  OAI22_X1 U324 ( .A1(n5390), .A2(\UUT/Mcontrol/N22 ), .B1(n329), .B2(n7396), 
        .ZN(n3020) );
  INV_X1 U325 ( .A(n340), .ZN(n329) );
  OAI211_X1 U326 ( .C1(n5990), .C2(n287), .A(n343), .B(n344), .ZN(n340) );
  AOI222_X1 U327 ( .A1(\UUT/Mpath/the_mult/x_mult_out[21] ), .A2(n6357), .B1(
        n320), .B2(n345), .C1(n291), .C2(n346), .ZN(n344) );
  INV_X1 U328 ( .A(n5609), .ZN(n346) );
  AOI22_X1 U330 ( .A1(n6397), .A2(n347), .B1(n324), .B2(n6116), .ZN(n343) );
  INV_X1 U331 ( .A(n5563), .ZN(n347) );
  OAI221_X1 U332 ( .B1(n348), .B2(n80), .C1(n68), .C2(n81), .A(n349), .ZN(
        n3021) );
  NAND2_X1 U333 ( .A1(\UUT/Mpath/the_mult/x_operand2 [20]), .A2(n6340), .ZN(
        n349) );
  OAI222_X1 U336 ( .A1(n68), .A2(n94), .B1(n348), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N44 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3023) );
  INV_X1 U337 ( .A(n351), .ZN(n68) );
  OAI222_X1 U338 ( .A1(n352), .A2(n99), .B1(n353), .B2(n101), .C1(n5392), .C2(
        n102), .ZN(n351) );
  OAI221_X1 U339 ( .B1(n103), .B2(n354), .C1(n5610), .C2(n105), .A(n355), .ZN(
        n3024) );
  AOI22_X1 U340 ( .A1(n107), .A2(n356), .B1(\UUT/Mpath/the_mult/Mad_out [52]), 
        .B2(n109), .ZN(n355) );
  OAI221_X1 U341 ( .B1(n115), .B2(n357), .C1(n5565), .C2(n117), .A(n358), .ZN(
        n3025) );
  AOI22_X1 U342 ( .A1(n119), .A2(n356), .B1(\UUT/Mpath/the_mult/Mad_out [20]), 
        .B2(n121), .ZN(n358) );
  OAI22_X1 U344 ( .A1(n7387), .A2(n359), .B1(n5566), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3026) );
  OAI221_X1 U345 ( .B1(n360), .B2(n124), .C1(n125), .C2(n359), .A(n361), .ZN(
        n3027) );
  AOI22_X1 U346 ( .A1(n127), .A2(n362), .B1(n129), .B2(n363), .ZN(n361) );
  OAI221_X1 U348 ( .B1(n360), .B2(n218), .C1(\UUT/Mpath/the_alu/N43 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n364), .ZN(n3028) );
  AOI22_X1 U349 ( .A1(n220), .A2(n362), .B1(n221), .B2(n363), .ZN(n364) );
  OAI22_X1 U350 ( .A1(n5302), .A2(n6393), .B1(n353), .B2(n223), .ZN(n3029) );
  OAI22_X1 U351 ( .A1(n5270), .A2(n6396), .B1(n353), .B2(n225), .ZN(n3030) );
  OAI22_X1 U352 ( .A1(n5238), .A2(n6387), .B1(n353), .B2(n227), .ZN(n3031) );
  OAI22_X1 U353 ( .A1(n5206), .A2(n6395), .B1(n353), .B2(n229), .ZN(n3032) );
  OAI22_X1 U354 ( .A1(n5174), .A2(n6390), .B1(n353), .B2(n231), .ZN(n3033) );
  OAI22_X1 U355 ( .A1(n5142), .A2(n6385), .B1(n353), .B2(n233), .ZN(n3034) );
  OAI22_X1 U356 ( .A1(n5110), .A2(n6389), .B1(n353), .B2(n235), .ZN(n3035) );
  OAI22_X1 U357 ( .A1(n5078), .A2(n6382), .B1(n353), .B2(n237), .ZN(n3036) );
  OAI22_X1 U358 ( .A1(n5046), .A2(n6380), .B1(n353), .B2(n239), .ZN(n3037) );
  OAI22_X1 U359 ( .A1(n5014), .A2(n6379), .B1(n353), .B2(n241), .ZN(n3038) );
  OAI22_X1 U360 ( .A1(n4982), .A2(n6376), .B1(n353), .B2(n243), .ZN(n3039) );
  OAI22_X1 U361 ( .A1(n4950), .A2(n6375), .B1(n353), .B2(n245), .ZN(n3040) );
  OAI22_X1 U362 ( .A1(n4918), .A2(n6372), .B1(n353), .B2(n247), .ZN(n3041) );
  OAI22_X1 U363 ( .A1(n4886), .A2(n6371), .B1(n353), .B2(n249), .ZN(n3042) );
  OAI22_X1 U364 ( .A1(n4854), .A2(n6368), .B1(n353), .B2(n251), .ZN(n3043) );
  OAI22_X1 U365 ( .A1(n4822), .A2(n6367), .B1(n353), .B2(n253), .ZN(n3044) );
  OAI22_X1 U366 ( .A1(n4790), .A2(n6364), .B1(n353), .B2(n255), .ZN(n3045) );
  OAI22_X1 U367 ( .A1(n4758), .A2(n6362), .B1(n353), .B2(n257), .ZN(n3046) );
  OAI22_X1 U368 ( .A1(n4726), .A2(n6361), .B1(n353), .B2(n259), .ZN(n3047) );
  OAI22_X1 U369 ( .A1(n4694), .A2(n6365), .B1(n353), .B2(n261), .ZN(n3048) );
  OAI22_X1 U370 ( .A1(n4662), .A2(n6366), .B1(n353), .B2(n263), .ZN(n3049) );
  OAI22_X1 U371 ( .A1(n4630), .A2(n6369), .B1(n353), .B2(n265), .ZN(n3050) );
  OAI22_X1 U372 ( .A1(n4598), .A2(n6370), .B1(n353), .B2(n267), .ZN(n3051) );
  OAI22_X1 U373 ( .A1(n4566), .A2(n6373), .B1(n353), .B2(n269), .ZN(n3052) );
  OAI22_X1 U374 ( .A1(n4534), .A2(n6374), .B1(n353), .B2(n271), .ZN(n3053) );
  OAI22_X1 U375 ( .A1(n4502), .A2(n6377), .B1(n353), .B2(n273), .ZN(n3054) );
  OAI22_X1 U376 ( .A1(n4470), .A2(n6378), .B1(n353), .B2(n275), .ZN(n3055) );
  OAI22_X1 U377 ( .A1(n4438), .A2(n6381), .B1(n353), .B2(n277), .ZN(n3056) );
  OAI22_X1 U378 ( .A1(n4406), .A2(n6384), .B1(n353), .B2(n279), .ZN(n3057) );
  OAI22_X1 U379 ( .A1(n4374), .A2(n6383), .B1(n353), .B2(n281), .ZN(n3058) );
  OAI22_X1 U380 ( .A1(n4342), .A2(n6391), .B1(n353), .B2(n283), .ZN(n3059) );
  OAI221_X1 U382 ( .B1(n365), .B2(n284), .C1(n5623), .C2(n5393), .A(n285), 
        .ZN(n362) );
  INV_X1 U383 ( .A(D_DATA_INBUS[20]), .ZN(n365) );
  OAI22_X1 U384 ( .A1(n5393), .A2(\UUT/Mcontrol/N22 ), .B1(n352), .B2(n7397), 
        .ZN(n3060) );
  INV_X1 U385 ( .A(n363), .ZN(n352) );
  OAI211_X1 U386 ( .C1(n6000), .C2(n287), .A(n366), .B(n367), .ZN(n363) );
  AOI222_X1 U387 ( .A1(\UUT/Mpath/the_mult/x_mult_out[20] ), .A2(n6357), .B1(
        n320), .B2(n368), .C1(n291), .C2(n369), .ZN(n367) );
  INV_X1 U388 ( .A(n5610), .ZN(n369) );
  AOI22_X1 U390 ( .A1(n6397), .A2(n370), .B1(n324), .B2(n6117), .ZN(n366) );
  INV_X1 U391 ( .A(n5565), .ZN(n370) );
  OAI221_X1 U392 ( .B1(n371), .B2(n80), .C1(n67), .C2(n81), .A(n372), .ZN(
        n3061) );
  NAND2_X1 U393 ( .A1(n6938), .A2(n6340), .ZN(n372) );
  INV_X1 U394 ( .A(n373), .ZN(n67) );
  AOI222_X1 U396 ( .A1(\UUT/jar_in [19]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [19]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [19]), 
        .C2(n301), .ZN(n374) );
  INV_X1 U397 ( .A(\UUT/break_code[19] ), .ZN(n371) );
  OAI211_X1 U398 ( .C1(\UUT/Mpath/the_alu/N46 ), .C2(\UUT/Mcontrol/N22 ), .A(
        n375), .B(n376), .ZN(n3063) );
  AOI222_X1 U399 ( .A1(n377), .A2(n373), .B1(n378), .B2(n6015), .C1(n96), .C2(
        \UUT/Mcontrol/d_sampled_finstr [3]), .ZN(n376) );
  OAI222_X1 U400 ( .A1(n379), .A2(n5332), .B1(n380), .B2(n101), .C1(n5398), 
        .C2(n102), .ZN(n373) );
  OAI221_X1 U401 ( .B1(n103), .B2(n381), .C1(n5612), .C2(n105), .A(n382), .ZN(
        n3064) );
  AOI22_X1 U402 ( .A1(n107), .A2(n383), .B1(\UUT/Mpath/the_mult/Mad_out [51]), 
        .B2(n109), .ZN(n382) );
  OAI221_X1 U403 ( .B1(n115), .B2(n384), .C1(n5569), .C2(n117), .A(n385), .ZN(
        n3065) );
  AOI22_X1 U404 ( .A1(n119), .A2(n383), .B1(\UUT/Mpath/the_mult/Mad_out [19]), 
        .B2(n121), .ZN(n385) );
  OAI22_X1 U406 ( .A1(n7387), .A2(n386), .B1(n5570), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3066) );
  OAI221_X1 U407 ( .B1(n387), .B2(n124), .C1(n125), .C2(n386), .A(n388), .ZN(
        n3067) );
  AOI22_X1 U408 ( .A1(n127), .A2(n389), .B1(n129), .B2(n390), .ZN(n388) );
  INV_X1 U409 ( .A(\UUT/Mpath/the_mult/x_operand1[19] ), .ZN(n386) );
  OAI221_X1 U410 ( .B1(n387), .B2(n218), .C1(\UUT/Mpath/the_alu/N45 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n391), .ZN(n3068) );
  AOI22_X1 U411 ( .A1(n220), .A2(n389), .B1(n221), .B2(n390), .ZN(n391) );
  OAI22_X1 U412 ( .A1(n5304), .A2(n6393), .B1(n380), .B2(n223), .ZN(n3069) );
  OAI22_X1 U413 ( .A1(n5272), .A2(n224), .B1(n380), .B2(n225), .ZN(n3070) );
  OAI22_X1 U414 ( .A1(n5240), .A2(n6387), .B1(n380), .B2(n227), .ZN(n3071) );
  OAI22_X1 U415 ( .A1(n5208), .A2(n6395), .B1(n380), .B2(n229), .ZN(n3072) );
  OAI22_X1 U416 ( .A1(n5176), .A2(n230), .B1(n380), .B2(n231), .ZN(n3073) );
  OAI22_X1 U417 ( .A1(n5144), .A2(n232), .B1(n380), .B2(n233), .ZN(n3074) );
  OAI22_X1 U418 ( .A1(n5112), .A2(n6389), .B1(n380), .B2(n235), .ZN(n3075) );
  OAI22_X1 U419 ( .A1(n5080), .A2(n236), .B1(n380), .B2(n237), .ZN(n3076) );
  OAI22_X1 U420 ( .A1(n5048), .A2(n238), .B1(n380), .B2(n239), .ZN(n3077) );
  OAI22_X1 U421 ( .A1(n5016), .A2(n240), .B1(n380), .B2(n241), .ZN(n3078) );
  OAI22_X1 U422 ( .A1(n4984), .A2(n242), .B1(n380), .B2(n243), .ZN(n3079) );
  OAI22_X1 U423 ( .A1(n4952), .A2(n244), .B1(n380), .B2(n245), .ZN(n3080) );
  OAI22_X1 U424 ( .A1(n4920), .A2(n246), .B1(n380), .B2(n247), .ZN(n3081) );
  OAI22_X1 U425 ( .A1(n4888), .A2(n248), .B1(n380), .B2(n249), .ZN(n3082) );
  OAI22_X1 U426 ( .A1(n4856), .A2(n250), .B1(n380), .B2(n251), .ZN(n3083) );
  OAI22_X1 U427 ( .A1(n4824), .A2(n252), .B1(n380), .B2(n253), .ZN(n3084) );
  OAI22_X1 U428 ( .A1(n4792), .A2(n6364), .B1(n380), .B2(n255), .ZN(n3085) );
  OAI22_X1 U429 ( .A1(n4760), .A2(n256), .B1(n380), .B2(n257), .ZN(n3086) );
  OAI22_X1 U430 ( .A1(n4728), .A2(n6361), .B1(n380), .B2(n259), .ZN(n3087) );
  OAI22_X1 U431 ( .A1(n4696), .A2(n260), .B1(n380), .B2(n261), .ZN(n3088) );
  OAI22_X1 U432 ( .A1(n4664), .A2(n262), .B1(n380), .B2(n263), .ZN(n3089) );
  OAI22_X1 U433 ( .A1(n4632), .A2(n264), .B1(n380), .B2(n265), .ZN(n3090) );
  OAI22_X1 U434 ( .A1(n4600), .A2(n266), .B1(n380), .B2(n267), .ZN(n3091) );
  OAI22_X1 U435 ( .A1(n4568), .A2(n268), .B1(n380), .B2(n269), .ZN(n3092) );
  OAI22_X1 U436 ( .A1(n4536), .A2(n270), .B1(n380), .B2(n271), .ZN(n3093) );
  OAI22_X1 U437 ( .A1(n4504), .A2(n272), .B1(n380), .B2(n273), .ZN(n3094) );
  OAI22_X1 U438 ( .A1(n4472), .A2(n274), .B1(n380), .B2(n275), .ZN(n3095) );
  OAI22_X1 U439 ( .A1(n4440), .A2(n276), .B1(n380), .B2(n277), .ZN(n3096) );
  OAI22_X1 U440 ( .A1(n4408), .A2(n278), .B1(n380), .B2(n279), .ZN(n3097) );
  OAI22_X1 U441 ( .A1(n4376), .A2(n280), .B1(n380), .B2(n281), .ZN(n3098) );
  OAI22_X1 U442 ( .A1(n4344), .A2(n282), .B1(n380), .B2(n283), .ZN(n3099) );
  OAI221_X1 U444 ( .B1(n392), .B2(n284), .C1(n5623), .C2(n5399), .A(n285), 
        .ZN(n389) );
  INV_X1 U445 ( .A(D_DATA_INBUS[19]), .ZN(n392) );
  OAI22_X1 U446 ( .A1(n5399), .A2(\UUT/Mcontrol/N22 ), .B1(n379), .B2(n7397), 
        .ZN(n3100) );
  INV_X1 U447 ( .A(n390), .ZN(n379) );
  OAI211_X1 U448 ( .C1(n6013), .C2(n287), .A(n393), .B(n394), .ZN(n390) );
  AOI222_X1 U449 ( .A1(\UUT/Mpath/the_mult/x_mult_out[19] ), .A2(n6357), .B1(
        n320), .B2(n395), .C1(n291), .C2(n396), .ZN(n394) );
  INV_X1 U450 ( .A(n5612), .ZN(n396) );
  AOI22_X1 U452 ( .A1(n6397), .A2(n397), .B1(n324), .B2(n6118), .ZN(n393) );
  INV_X1 U453 ( .A(n5569), .ZN(n397) );
  OAI221_X1 U454 ( .B1(n398), .B2(n80), .C1(n66), .C2(n81), .A(n399), .ZN(
        n3101) );
  NAND2_X1 U455 ( .A1(\UUT/Mpath/the_mult/x_operand2 [18]), .A2(n6340), .ZN(
        n399) );
  INV_X1 U456 ( .A(n400), .ZN(n66) );
  AOI222_X1 U458 ( .A1(\UUT/jar_in [18]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [18]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [18]), 
        .C2(n301), .ZN(n401) );
  INV_X1 U459 ( .A(\UUT/break_code[18] ), .ZN(n398) );
  OAI211_X1 U460 ( .C1(\UUT/Mpath/the_alu/N48 ), .C2(\UUT/Mcontrol/N22 ), .A(
        n375), .B(n402), .ZN(n3103) );
  AOI222_X1 U461 ( .A1(n377), .A2(n400), .B1(n6027), .B2(n378), .C1(n96), .C2(
        \UUT/Mcontrol/d_sampled_finstr [2]), .ZN(n402) );
  OAI222_X1 U462 ( .A1(n403), .A2(n99), .B1(n404), .B2(n101), .C1(n5401), .C2(
        n102), .ZN(n400) );
  OAI221_X1 U463 ( .B1(n103), .B2(n405), .C1(n5613), .C2(n105), .A(n406), .ZN(
        n3104) );
  AOI22_X1 U464 ( .A1(n107), .A2(n407), .B1(\UUT/Mpath/the_mult/Mad_out [50]), 
        .B2(n109), .ZN(n406) );
  OAI221_X1 U465 ( .B1(n115), .B2(n408), .C1(n5571), .C2(n117), .A(n409), .ZN(
        n3105) );
  AOI22_X1 U466 ( .A1(n119), .A2(n407), .B1(\UUT/Mpath/the_mult/Mad_out [18]), 
        .B2(n121), .ZN(n409) );
  OAI22_X1 U468 ( .A1(n7387), .A2(n410), .B1(n5572), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3106) );
  OAI221_X1 U469 ( .B1(n411), .B2(n124), .C1(n125), .C2(n410), .A(n412), .ZN(
        n3107) );
  AOI22_X1 U470 ( .A1(n127), .A2(n413), .B1(n129), .B2(n414), .ZN(n412) );
  INV_X1 U471 ( .A(\UUT/Mpath/the_mult/x_operand1[18] ), .ZN(n410) );
  OAI221_X1 U472 ( .B1(n411), .B2(n218), .C1(\UUT/Mpath/the_alu/N47 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n415), .ZN(n3108) );
  AOI22_X1 U473 ( .A1(n220), .A2(n413), .B1(n221), .B2(n414), .ZN(n415) );
  OAI22_X1 U474 ( .A1(n5305), .A2(n6393), .B1(n404), .B2(n223), .ZN(n3109) );
  OAI22_X1 U475 ( .A1(n5273), .A2(n6396), .B1(n404), .B2(n225), .ZN(n3110) );
  OAI22_X1 U476 ( .A1(n5241), .A2(n6387), .B1(n404), .B2(n227), .ZN(n3111) );
  OAI22_X1 U477 ( .A1(n5209), .A2(n6395), .B1(n404), .B2(n229), .ZN(n3112) );
  OAI22_X1 U478 ( .A1(n5177), .A2(n6390), .B1(n404), .B2(n231), .ZN(n3113) );
  OAI22_X1 U479 ( .A1(n5145), .A2(n6385), .B1(n404), .B2(n233), .ZN(n3114) );
  OAI22_X1 U480 ( .A1(n5113), .A2(n6389), .B1(n404), .B2(n235), .ZN(n3115) );
  OAI22_X1 U481 ( .A1(n5081), .A2(n6382), .B1(n404), .B2(n237), .ZN(n3116) );
  OAI22_X1 U482 ( .A1(n5049), .A2(n6380), .B1(n404), .B2(n239), .ZN(n3117) );
  OAI22_X1 U483 ( .A1(n5017), .A2(n6379), .B1(n404), .B2(n241), .ZN(n3118) );
  OAI22_X1 U484 ( .A1(n4985), .A2(n6376), .B1(n404), .B2(n243), .ZN(n3119) );
  OAI22_X1 U485 ( .A1(n4953), .A2(n6375), .B1(n404), .B2(n245), .ZN(n3120) );
  OAI22_X1 U486 ( .A1(n4921), .A2(n6372), .B1(n404), .B2(n247), .ZN(n3121) );
  OAI22_X1 U487 ( .A1(n4889), .A2(n6371), .B1(n404), .B2(n249), .ZN(n3122) );
  OAI22_X1 U488 ( .A1(n4857), .A2(n6368), .B1(n404), .B2(n251), .ZN(n3123) );
  OAI22_X1 U489 ( .A1(n4825), .A2(n6367), .B1(n404), .B2(n253), .ZN(n3124) );
  OAI22_X1 U490 ( .A1(n4793), .A2(n6364), .B1(n404), .B2(n255), .ZN(n3125) );
  OAI22_X1 U491 ( .A1(n4761), .A2(n6362), .B1(n404), .B2(n257), .ZN(n3126) );
  OAI22_X1 U492 ( .A1(n4729), .A2(n6361), .B1(n404), .B2(n259), .ZN(n3127) );
  OAI22_X1 U493 ( .A1(n4697), .A2(n6365), .B1(n404), .B2(n261), .ZN(n3128) );
  OAI22_X1 U494 ( .A1(n4665), .A2(n6366), .B1(n404), .B2(n263), .ZN(n3129) );
  OAI22_X1 U495 ( .A1(n4633), .A2(n6369), .B1(n404), .B2(n265), .ZN(n3130) );
  OAI22_X1 U496 ( .A1(n4601), .A2(n6370), .B1(n404), .B2(n267), .ZN(n3131) );
  OAI22_X1 U497 ( .A1(n4569), .A2(n6373), .B1(n404), .B2(n269), .ZN(n3132) );
  OAI22_X1 U498 ( .A1(n4537), .A2(n6374), .B1(n404), .B2(n271), .ZN(n3133) );
  OAI22_X1 U499 ( .A1(n4505), .A2(n6377), .B1(n404), .B2(n273), .ZN(n3134) );
  OAI22_X1 U500 ( .A1(n4473), .A2(n6378), .B1(n404), .B2(n275), .ZN(n3135) );
  OAI22_X1 U501 ( .A1(n4441), .A2(n6381), .B1(n404), .B2(n277), .ZN(n3136) );
  OAI22_X1 U502 ( .A1(n4409), .A2(n6384), .B1(n404), .B2(n279), .ZN(n3137) );
  OAI22_X1 U503 ( .A1(n4377), .A2(n6383), .B1(n404), .B2(n281), .ZN(n3138) );
  OAI22_X1 U504 ( .A1(n4345), .A2(n6391), .B1(n404), .B2(n283), .ZN(n3139) );
  OAI221_X1 U506 ( .B1(n416), .B2(n284), .C1(n5623), .C2(n5402), .A(n285), 
        .ZN(n413) );
  INV_X1 U507 ( .A(D_DATA_INBUS[18]), .ZN(n416) );
  OAI22_X1 U508 ( .A1(n5402), .A2(\UUT/Mcontrol/N22 ), .B1(n403), .B2(n7396), 
        .ZN(n3140) );
  INV_X1 U509 ( .A(n414), .ZN(n403) );
  OAI211_X1 U510 ( .C1(n6026), .C2(n287), .A(n417), .B(n418), .ZN(n414) );
  AOI222_X1 U511 ( .A1(\UUT/Mpath/the_mult/x_mult_out[18] ), .A2(n6357), .B1(
        n320), .B2(n419), .C1(n291), .C2(n420), .ZN(n418) );
  INV_X1 U512 ( .A(n5613), .ZN(n420) );
  AOI22_X1 U514 ( .A1(n6397), .A2(n421), .B1(n324), .B2(n6119), .ZN(n417) );
  INV_X1 U515 ( .A(n5571), .ZN(n421) );
  OAI221_X1 U516 ( .B1(n422), .B2(n80), .C1(n65), .C2(n81), .A(n423), .ZN(
        n3141) );
  NAND2_X1 U517 ( .A1(n6915), .A2(n6340), .ZN(n423) );
  INV_X1 U518 ( .A(n424), .ZN(n65) );
  AOI222_X1 U520 ( .A1(\UUT/jar_in [17]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [17]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [17]), 
        .C2(n301), .ZN(n425) );
  INV_X1 U521 ( .A(\UUT/break_code[17] ), .ZN(n422) );
  OAI211_X1 U522 ( .C1(\UUT/Mpath/the_alu/N50 ), .C2(\UUT/Mcontrol/N22 ), .A(
        n375), .B(n426), .ZN(n3143) );
  AOI222_X1 U523 ( .A1(n377), .A2(n424), .B1(n6048), .B2(n378), .C1(n96), .C2(
        \UUT/Mcontrol/d_sampled_finstr [1]), .ZN(n426) );
  OAI222_X1 U524 ( .A1(n427), .A2(n99), .B1(n428), .B2(n101), .C1(n5404), .C2(
        n102), .ZN(n424) );
  OAI221_X1 U525 ( .B1(n103), .B2(n429), .C1(n5614), .C2(n105), .A(n430), .ZN(
        n3144) );
  AOI22_X1 U526 ( .A1(n107), .A2(n431), .B1(\UUT/Mpath/the_mult/Mad_out [49]), 
        .B2(n109), .ZN(n430) );
  OAI221_X1 U527 ( .B1(n115), .B2(n432), .C1(n5573), .C2(n117), .A(n433), .ZN(
        n3145) );
  AOI22_X1 U528 ( .A1(n119), .A2(n431), .B1(\UUT/Mpath/the_mult/Mad_out [17]), 
        .B2(n121), .ZN(n433) );
  OAI22_X1 U530 ( .A1(n7386), .A2(n434), .B1(n5574), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3146) );
  OAI221_X1 U531 ( .B1(n435), .B2(n124), .C1(n125), .C2(n434), .A(n436), .ZN(
        n3147) );
  AOI22_X1 U532 ( .A1(n127), .A2(n437), .B1(n129), .B2(n438), .ZN(n436) );
  INV_X1 U533 ( .A(\UUT/Mpath/the_mult/x_operand1[17] ), .ZN(n434) );
  OAI221_X1 U534 ( .B1(n435), .B2(n218), .C1(\UUT/Mpath/the_alu/N49 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n439), .ZN(n3148) );
  AOI22_X1 U535 ( .A1(n220), .A2(n437), .B1(n221), .B2(n438), .ZN(n439) );
  OAI22_X1 U536 ( .A1(n5306), .A2(n6393), .B1(n428), .B2(n223), .ZN(n3149) );
  OAI22_X1 U537 ( .A1(n5274), .A2(n6396), .B1(n428), .B2(n225), .ZN(n3150) );
  OAI22_X1 U538 ( .A1(n5242), .A2(n6387), .B1(n428), .B2(n227), .ZN(n3151) );
  OAI22_X1 U539 ( .A1(n5210), .A2(n6395), .B1(n428), .B2(n229), .ZN(n3152) );
  OAI22_X1 U540 ( .A1(n5178), .A2(n6390), .B1(n428), .B2(n231), .ZN(n3153) );
  OAI22_X1 U541 ( .A1(n5146), .A2(n6385), .B1(n428), .B2(n233), .ZN(n3154) );
  OAI22_X1 U542 ( .A1(n5114), .A2(n6389), .B1(n428), .B2(n235), .ZN(n3155) );
  OAI22_X1 U543 ( .A1(n5082), .A2(n6382), .B1(n428), .B2(n237), .ZN(n3156) );
  OAI22_X1 U544 ( .A1(n5050), .A2(n6380), .B1(n428), .B2(n239), .ZN(n3157) );
  OAI22_X1 U545 ( .A1(n5018), .A2(n6379), .B1(n428), .B2(n241), .ZN(n3158) );
  OAI22_X1 U546 ( .A1(n4986), .A2(n6376), .B1(n428), .B2(n243), .ZN(n3159) );
  OAI22_X1 U547 ( .A1(n4954), .A2(n6375), .B1(n428), .B2(n245), .ZN(n3160) );
  OAI22_X1 U548 ( .A1(n4922), .A2(n6372), .B1(n428), .B2(n247), .ZN(n3161) );
  OAI22_X1 U549 ( .A1(n4890), .A2(n6371), .B1(n428), .B2(n249), .ZN(n3162) );
  OAI22_X1 U550 ( .A1(n4858), .A2(n6368), .B1(n428), .B2(n251), .ZN(n3163) );
  OAI22_X1 U551 ( .A1(n4826), .A2(n6367), .B1(n428), .B2(n253), .ZN(n3164) );
  OAI22_X1 U552 ( .A1(n4794), .A2(n6364), .B1(n428), .B2(n255), .ZN(n3165) );
  OAI22_X1 U553 ( .A1(n4762), .A2(n6362), .B1(n428), .B2(n257), .ZN(n3166) );
  OAI22_X1 U554 ( .A1(n4730), .A2(n6361), .B1(n428), .B2(n259), .ZN(n3167) );
  OAI22_X1 U555 ( .A1(n4698), .A2(n6365), .B1(n428), .B2(n261), .ZN(n3168) );
  OAI22_X1 U556 ( .A1(n4666), .A2(n6366), .B1(n428), .B2(n263), .ZN(n3169) );
  OAI22_X1 U557 ( .A1(n4634), .A2(n6369), .B1(n428), .B2(n265), .ZN(n3170) );
  OAI22_X1 U558 ( .A1(n4602), .A2(n6370), .B1(n428), .B2(n267), .ZN(n3171) );
  OAI22_X1 U559 ( .A1(n4570), .A2(n6373), .B1(n428), .B2(n269), .ZN(n3172) );
  OAI22_X1 U560 ( .A1(n4538), .A2(n6374), .B1(n428), .B2(n271), .ZN(n3173) );
  OAI22_X1 U561 ( .A1(n4506), .A2(n6377), .B1(n428), .B2(n273), .ZN(n3174) );
  OAI22_X1 U562 ( .A1(n4474), .A2(n6378), .B1(n428), .B2(n275), .ZN(n3175) );
  OAI22_X1 U563 ( .A1(n4442), .A2(n6381), .B1(n428), .B2(n277), .ZN(n3176) );
  OAI22_X1 U564 ( .A1(n4410), .A2(n6384), .B1(n428), .B2(n279), .ZN(n3177) );
  OAI22_X1 U565 ( .A1(n4378), .A2(n6383), .B1(n428), .B2(n281), .ZN(n3178) );
  OAI22_X1 U566 ( .A1(n4346), .A2(n6391), .B1(n428), .B2(n283), .ZN(n3179) );
  OAI221_X1 U568 ( .B1(n440), .B2(n284), .C1(n5623), .C2(n5405), .A(n285), 
        .ZN(n437) );
  INV_X1 U569 ( .A(D_DATA_INBUS[17]), .ZN(n440) );
  OAI22_X1 U570 ( .A1(n5405), .A2(\UUT/Mcontrol/N22 ), .B1(n427), .B2(n7396), 
        .ZN(n3180) );
  INV_X1 U571 ( .A(n438), .ZN(n427) );
  OAI211_X1 U572 ( .C1(n6047), .C2(n287), .A(n441), .B(n442), .ZN(n438) );
  AOI222_X1 U573 ( .A1(\UUT/Mpath/the_mult/x_mult_out[17] ), .A2(n6357), .B1(
        n320), .B2(n443), .C1(n291), .C2(n444), .ZN(n442) );
  INV_X1 U574 ( .A(n5614), .ZN(n444) );
  AOI22_X1 U576 ( .A1(n6397), .A2(n445), .B1(n324), .B2(n6120), .ZN(n441) );
  INV_X1 U577 ( .A(n5573), .ZN(n445) );
  OAI221_X1 U578 ( .B1(n446), .B2(n80), .C1(n64), .C2(n81), .A(n447), .ZN(
        n3181) );
  NAND2_X1 U579 ( .A1(\UUT/Mpath/the_mult/x_operand2 [16]), .A2(n6340), .ZN(
        n447) );
  INV_X1 U580 ( .A(n448), .ZN(n64) );
  INV_X1 U583 ( .A(\UUT/break_code[16] ), .ZN(n446) );
  OAI211_X1 U584 ( .C1(\UUT/Mpath/the_alu/N52 ), .C2(\UUT/Mcontrol/N22 ), .A(
        n375), .B(n450), .ZN(n3183) );
  AOI222_X1 U585 ( .A1(n377), .A2(n448), .B1(n6060), .B2(n378), .C1(n96), .C2(
        \UUT/Mcontrol/d_sampled_finstr [0]), .ZN(n450) );
  AND2_X1 U587 ( .A1(n452), .A2(n6996), .ZN(n378) );
  OAI222_X1 U588 ( .A1(n454), .A2(n99), .B1(n455), .B2(n101), .C1(n5407), .C2(
        n102), .ZN(n448) );
  INV_X1 U589 ( .A(n94), .ZN(n377) );
  AOI22_X1 U590 ( .A1(n456), .A2(n457), .B1(n6016), .B2(n452), .ZN(n375) );
  NOR3_X1 U591 ( .A1(n7382), .A2(n7095), .A3(n203), .ZN(n452) );
  OAI221_X1 U592 ( .B1(n103), .B2(n458), .C1(n5615), .C2(n105), .A(n459), .ZN(
        n3184) );
  AOI22_X1 U593 ( .A1(n107), .A2(n460), .B1(\UUT/Mpath/the_mult/Mad_out [48]), 
        .B2(n109), .ZN(n459) );
  OAI221_X1 U594 ( .B1(n115), .B2(n461), .C1(n5575), .C2(n117), .A(n462), .ZN(
        n3185) );
  AOI22_X1 U595 ( .A1(n119), .A2(n460), .B1(\UUT/Mpath/the_mult/Mad_out [16]), 
        .B2(n121), .ZN(n462) );
  OAI22_X1 U597 ( .A1(n7386), .A2(n463), .B1(n5576), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3186) );
  OAI221_X1 U598 ( .B1(n464), .B2(n124), .C1(n125), .C2(n463), .A(n465), .ZN(
        n3187) );
  AOI22_X1 U599 ( .A1(n127), .A2(n466), .B1(n129), .B2(n467), .ZN(n465) );
  INV_X1 U600 ( .A(\UUT/Mpath/the_mult/x_operand1[16] ), .ZN(n463) );
  OAI221_X1 U601 ( .B1(n464), .B2(n218), .C1(\UUT/Mpath/the_alu/N51 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n468), .ZN(n3188) );
  AOI22_X1 U602 ( .A1(n220), .A2(n466), .B1(n221), .B2(n467), .ZN(n468) );
  OAI22_X1 U603 ( .A1(n5307), .A2(n6393), .B1(n455), .B2(n223), .ZN(n3189) );
  OAI22_X1 U604 ( .A1(n5275), .A2(n6396), .B1(n455), .B2(n225), .ZN(n3190) );
  OAI22_X1 U605 ( .A1(n5243), .A2(n6387), .B1(n455), .B2(n227), .ZN(n3191) );
  OAI22_X1 U606 ( .A1(n5211), .A2(n6395), .B1(n455), .B2(n229), .ZN(n3192) );
  OAI22_X1 U607 ( .A1(n5179), .A2(n6390), .B1(n455), .B2(n231), .ZN(n3193) );
  OAI22_X1 U608 ( .A1(n5147), .A2(n6385), .B1(n455), .B2(n233), .ZN(n3194) );
  OAI22_X1 U609 ( .A1(n5115), .A2(n6389), .B1(n455), .B2(n235), .ZN(n3195) );
  OAI22_X1 U610 ( .A1(n5083), .A2(n6382), .B1(n455), .B2(n237), .ZN(n3196) );
  OAI22_X1 U611 ( .A1(n5051), .A2(n6380), .B1(n455), .B2(n239), .ZN(n3197) );
  OAI22_X1 U612 ( .A1(n5019), .A2(n6379), .B1(n455), .B2(n241), .ZN(n3198) );
  OAI22_X1 U613 ( .A1(n4987), .A2(n6376), .B1(n455), .B2(n243), .ZN(n3199) );
  OAI22_X1 U614 ( .A1(n4955), .A2(n6375), .B1(n455), .B2(n245), .ZN(n3200) );
  OAI22_X1 U615 ( .A1(n4923), .A2(n6372), .B1(n455), .B2(n247), .ZN(n3201) );
  OAI22_X1 U616 ( .A1(n4891), .A2(n6371), .B1(n455), .B2(n249), .ZN(n3202) );
  OAI22_X1 U617 ( .A1(n4859), .A2(n6368), .B1(n455), .B2(n251), .ZN(n3203) );
  OAI22_X1 U618 ( .A1(n4827), .A2(n6367), .B1(n455), .B2(n253), .ZN(n3204) );
  OAI22_X1 U619 ( .A1(n4795), .A2(n6364), .B1(n455), .B2(n255), .ZN(n3205) );
  OAI22_X1 U620 ( .A1(n4763), .A2(n6362), .B1(n455), .B2(n257), .ZN(n3206) );
  OAI22_X1 U621 ( .A1(n4731), .A2(n6361), .B1(n455), .B2(n259), .ZN(n3207) );
  OAI22_X1 U622 ( .A1(n4699), .A2(n6365), .B1(n455), .B2(n261), .ZN(n3208) );
  OAI22_X1 U623 ( .A1(n4667), .A2(n6366), .B1(n455), .B2(n263), .ZN(n3209) );
  OAI22_X1 U624 ( .A1(n4635), .A2(n6369), .B1(n455), .B2(n265), .ZN(n3210) );
  OAI22_X1 U625 ( .A1(n4603), .A2(n6370), .B1(n455), .B2(n267), .ZN(n3211) );
  OAI22_X1 U626 ( .A1(n4571), .A2(n6373), .B1(n455), .B2(n269), .ZN(n3212) );
  OAI22_X1 U627 ( .A1(n4539), .A2(n6374), .B1(n455), .B2(n271), .ZN(n3213) );
  OAI22_X1 U628 ( .A1(n4507), .A2(n6377), .B1(n455), .B2(n273), .ZN(n3214) );
  OAI22_X1 U629 ( .A1(n4475), .A2(n6378), .B1(n455), .B2(n275), .ZN(n3215) );
  OAI22_X1 U630 ( .A1(n4443), .A2(n6381), .B1(n455), .B2(n277), .ZN(n3216) );
  OAI22_X1 U631 ( .A1(n4411), .A2(n6384), .B1(n455), .B2(n279), .ZN(n3217) );
  OAI22_X1 U632 ( .A1(n4379), .A2(n6383), .B1(n455), .B2(n281), .ZN(n3218) );
  OAI22_X1 U633 ( .A1(n4347), .A2(n6391), .B1(n455), .B2(n283), .ZN(n3219) );
  OAI221_X1 U635 ( .B1(n469), .B2(n284), .C1(n5623), .C2(n5408), .A(n285), 
        .ZN(n466) );
  INV_X1 U636 ( .A(D_DATA_INBUS[16]), .ZN(n469) );
  OAI22_X1 U637 ( .A1(n5408), .A2(\UUT/Mcontrol/N22 ), .B1(n454), .B2(n7396), 
        .ZN(n3220) );
  INV_X1 U638 ( .A(n467), .ZN(n454) );
  OAI211_X1 U639 ( .C1(n6059), .C2(n287), .A(n470), .B(n471), .ZN(n467) );
  AOI222_X1 U640 ( .A1(\UUT/Mpath/the_mult/x_mult_out[16] ), .A2(n6357), .B1(
        n320), .B2(n472), .C1(n291), .C2(n473), .ZN(n471) );
  INV_X1 U641 ( .A(n5615), .ZN(n473) );
  AOI22_X1 U643 ( .A1(n6397), .A2(n474), .B1(n324), .B2(n6121), .ZN(n470) );
  INV_X1 U644 ( .A(n5575), .ZN(n474) );
  OAI221_X1 U645 ( .B1(n475), .B2(n80), .C1(n63), .C2(n81), .A(n476), .ZN(
        n3221) );
  NAND2_X1 U646 ( .A1(n7091), .A2(n6340), .ZN(n476) );
  AOI222_X1 U648 ( .A1(\UUT/jar_in [15]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [15]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [15]), 
        .C2(n301), .ZN(n478) );
  OAI222_X1 U649 ( .A1(n63), .A2(n94), .B1(n477), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N54 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3223) );
  INV_X1 U651 ( .A(n483), .ZN(n63) );
  OAI222_X1 U652 ( .A1(n484), .A2(n5332), .B1(n485), .B2(n101), .C1(n5410), 
        .C2(n102), .ZN(n483) );
  OAI221_X1 U653 ( .B1(n103), .B2(n486), .C1(n5616), .C2(n105), .A(n487), .ZN(
        n3224) );
  AOI22_X1 U654 ( .A1(n107), .A2(n488), .B1(\UUT/Mpath/the_mult/Mad_out [47]), 
        .B2(n109), .ZN(n487) );
  OAI221_X1 U655 ( .B1(n115), .B2(n489), .C1(n5577), .C2(n117), .A(n490), .ZN(
        n3225) );
  AOI22_X1 U656 ( .A1(n119), .A2(n488), .B1(\UUT/Mpath/the_mult/Mad_out [15]), 
        .B2(n121), .ZN(n490) );
  OAI22_X1 U658 ( .A1(n7385), .A2(n491), .B1(n5578), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3226) );
  OAI221_X1 U659 ( .B1(n492), .B2(n124), .C1(n125), .C2(n491), .A(n493), .ZN(
        n3227) );
  AOI22_X1 U660 ( .A1(n127), .A2(n494), .B1(n129), .B2(n495), .ZN(n493) );
  INV_X1 U661 ( .A(\UUT/Mpath/the_mult/x_operand1[15] ), .ZN(n491) );
  OAI221_X1 U662 ( .B1(n492), .B2(n218), .C1(\UUT/Mpath/the_alu/N53 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n496), .ZN(n3228) );
  AOI22_X1 U663 ( .A1(n220), .A2(n494), .B1(n221), .B2(n495), .ZN(n496) );
  INV_X1 U664 ( .A(n485), .ZN(n494) );
  OAI22_X1 U665 ( .A1(n5308), .A2(n6393), .B1(n485), .B2(n223), .ZN(n3229) );
  OAI22_X1 U666 ( .A1(n5276), .A2(n6396), .B1(n485), .B2(n225), .ZN(n3230) );
  OAI22_X1 U667 ( .A1(n5244), .A2(n6387), .B1(n485), .B2(n227), .ZN(n3231) );
  OAI22_X1 U668 ( .A1(n5212), .A2(n6395), .B1(n485), .B2(n229), .ZN(n3232) );
  OAI22_X1 U669 ( .A1(n5180), .A2(n6390), .B1(n485), .B2(n231), .ZN(n3233) );
  OAI22_X1 U670 ( .A1(n5148), .A2(n6385), .B1(n485), .B2(n233), .ZN(n3234) );
  OAI22_X1 U671 ( .A1(n5116), .A2(n6389), .B1(n485), .B2(n235), .ZN(n3235) );
  OAI22_X1 U672 ( .A1(n5084), .A2(n6382), .B1(n485), .B2(n237), .ZN(n3236) );
  OAI22_X1 U673 ( .A1(n5052), .A2(n6380), .B1(n485), .B2(n239), .ZN(n3237) );
  OAI22_X1 U674 ( .A1(n5020), .A2(n6379), .B1(n485), .B2(n241), .ZN(n3238) );
  OAI22_X1 U675 ( .A1(n4988), .A2(n6376), .B1(n485), .B2(n243), .ZN(n3239) );
  OAI22_X1 U676 ( .A1(n4956), .A2(n6375), .B1(n485), .B2(n245), .ZN(n3240) );
  OAI22_X1 U677 ( .A1(n4924), .A2(n6372), .B1(n485), .B2(n247), .ZN(n3241) );
  OAI22_X1 U678 ( .A1(n4892), .A2(n6371), .B1(n485), .B2(n249), .ZN(n3242) );
  OAI22_X1 U679 ( .A1(n4860), .A2(n6368), .B1(n485), .B2(n251), .ZN(n3243) );
  OAI22_X1 U680 ( .A1(n4828), .A2(n6367), .B1(n485), .B2(n253), .ZN(n3244) );
  OAI22_X1 U681 ( .A1(n4796), .A2(n6364), .B1(n485), .B2(n255), .ZN(n3245) );
  OAI22_X1 U682 ( .A1(n4764), .A2(n6362), .B1(n485), .B2(n257), .ZN(n3246) );
  OAI22_X1 U683 ( .A1(n4732), .A2(n6361), .B1(n485), .B2(n259), .ZN(n3247) );
  OAI22_X1 U684 ( .A1(n4700), .A2(n6365), .B1(n485), .B2(n261), .ZN(n3248) );
  OAI22_X1 U685 ( .A1(n4668), .A2(n6366), .B1(n485), .B2(n263), .ZN(n3249) );
  OAI22_X1 U686 ( .A1(n4636), .A2(n6369), .B1(n485), .B2(n265), .ZN(n3250) );
  OAI22_X1 U687 ( .A1(n4604), .A2(n6370), .B1(n485), .B2(n267), .ZN(n3251) );
  OAI22_X1 U688 ( .A1(n4572), .A2(n6373), .B1(n485), .B2(n269), .ZN(n3252) );
  OAI22_X1 U689 ( .A1(n4540), .A2(n6374), .B1(n485), .B2(n271), .ZN(n3253) );
  OAI22_X1 U690 ( .A1(n4508), .A2(n6377), .B1(n485), .B2(n273), .ZN(n3254) );
  OAI22_X1 U691 ( .A1(n4476), .A2(n6378), .B1(n485), .B2(n275), .ZN(n3255) );
  OAI22_X1 U692 ( .A1(n4444), .A2(n6381), .B1(n485), .B2(n277), .ZN(n3256) );
  OAI22_X1 U693 ( .A1(n4412), .A2(n6384), .B1(n485), .B2(n279), .ZN(n3257) );
  OAI22_X1 U694 ( .A1(n4380), .A2(n6383), .B1(n485), .B2(n281), .ZN(n3258) );
  OAI22_X1 U695 ( .A1(n4348), .A2(n6391), .B1(n485), .B2(n283), .ZN(n3259) );
  OAI22_X1 U697 ( .A1(n501), .A2(n5668), .B1(n5411), .B2(n5623), .ZN(n500) );
  INV_X1 U698 ( .A(n5666), .ZN(n497) );
  OAI22_X1 U699 ( .A1(n5411), .A2(\UUT/Mcontrol/N22 ), .B1(n484), .B2(n7396), 
        .ZN(n3260) );
  INV_X1 U700 ( .A(n495), .ZN(n484) );
  OAI211_X1 U701 ( .C1(n6070), .C2(n287), .A(n502), .B(n503), .ZN(n495) );
  AOI222_X1 U702 ( .A1(\UUT/Mpath/the_mult/x_mult_out[15] ), .A2(n6357), .B1(
        n320), .B2(n504), .C1(n291), .C2(n505), .ZN(n503) );
  INV_X1 U703 ( .A(n5616), .ZN(n505) );
  AOI22_X1 U705 ( .A1(n6397), .A2(n506), .B1(n324), .B2(n6122), .ZN(n502) );
  INV_X1 U706 ( .A(n5577), .ZN(n506) );
  OAI221_X1 U707 ( .B1(n507), .B2(n80), .C1(n62), .C2(n81), .A(n508), .ZN(
        n3261) );
  NAND2_X1 U708 ( .A1(\UUT/Mpath/the_mult/x_operand2 [14]), .A2(n6340), .ZN(
        n508) );
  AOI222_X1 U710 ( .A1(\UUT/jar_in [14]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [14]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [14]), 
        .C2(n301), .ZN(n509) );
  OAI222_X1 U711 ( .A1(n62), .A2(n94), .B1(n507), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N56 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3263) );
  INV_X1 U712 ( .A(\UUT/break_code[14] ), .ZN(n507) );
  INV_X1 U713 ( .A(n510), .ZN(n62) );
  OAI222_X1 U714 ( .A1(n511), .A2(n99), .B1(n512), .B2(n101), .C1(n5413), .C2(
        n102), .ZN(n510) );
  OAI221_X1 U715 ( .B1(n103), .B2(n513), .C1(n5617), .C2(n105), .A(n514), .ZN(
        n3264) );
  AOI22_X1 U716 ( .A1(n107), .A2(n515), .B1(\UUT/Mpath/the_mult/Mad_out [46]), 
        .B2(n109), .ZN(n514) );
  OAI221_X1 U717 ( .B1(n115), .B2(n516), .C1(n5579), .C2(n117), .A(n517), .ZN(
        n3265) );
  AOI22_X1 U718 ( .A1(n119), .A2(n515), .B1(\UUT/Mpath/the_mult/Mad_out [14]), 
        .B2(n121), .ZN(n517) );
  OAI22_X1 U720 ( .A1(n7386), .A2(n518), .B1(n5580), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3266) );
  OAI221_X1 U721 ( .B1(n519), .B2(n124), .C1(n125), .C2(n518), .A(n520), .ZN(
        n3267) );
  AOI22_X1 U722 ( .A1(n127), .A2(n521), .B1(n129), .B2(n522), .ZN(n520) );
  INV_X1 U723 ( .A(\UUT/Mpath/the_mult/x_operand1[14] ), .ZN(n518) );
  OAI221_X1 U724 ( .B1(n519), .B2(n218), .C1(\UUT/Mpath/the_alu/N55 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n523), .ZN(n3268) );
  AOI22_X1 U725 ( .A1(n220), .A2(n521), .B1(n221), .B2(n522), .ZN(n523) );
  INV_X1 U726 ( .A(n512), .ZN(n521) );
  OAI22_X1 U727 ( .A1(n5309), .A2(n6393), .B1(n512), .B2(n223), .ZN(n3269) );
  OAI22_X1 U728 ( .A1(n5277), .A2(n6396), .B1(n512), .B2(n225), .ZN(n3270) );
  OAI22_X1 U729 ( .A1(n5245), .A2(n6387), .B1(n512), .B2(n227), .ZN(n3271) );
  OAI22_X1 U730 ( .A1(n5213), .A2(n6395), .B1(n512), .B2(n229), .ZN(n3272) );
  OAI22_X1 U731 ( .A1(n5181), .A2(n6390), .B1(n512), .B2(n231), .ZN(n3273) );
  OAI22_X1 U732 ( .A1(n5149), .A2(n6385), .B1(n512), .B2(n233), .ZN(n3274) );
  OAI22_X1 U733 ( .A1(n5117), .A2(n6389), .B1(n512), .B2(n235), .ZN(n3275) );
  OAI22_X1 U734 ( .A1(n5085), .A2(n6382), .B1(n512), .B2(n237), .ZN(n3276) );
  OAI22_X1 U735 ( .A1(n5053), .A2(n6380), .B1(n512), .B2(n239), .ZN(n3277) );
  OAI22_X1 U736 ( .A1(n5021), .A2(n6379), .B1(n512), .B2(n241), .ZN(n3278) );
  OAI22_X1 U737 ( .A1(n4989), .A2(n6376), .B1(n512), .B2(n243), .ZN(n3279) );
  OAI22_X1 U738 ( .A1(n4957), .A2(n6375), .B1(n512), .B2(n245), .ZN(n3280) );
  OAI22_X1 U739 ( .A1(n4925), .A2(n6372), .B1(n512), .B2(n247), .ZN(n3281) );
  OAI22_X1 U740 ( .A1(n4893), .A2(n6371), .B1(n512), .B2(n249), .ZN(n3282) );
  OAI22_X1 U741 ( .A1(n4861), .A2(n6368), .B1(n512), .B2(n251), .ZN(n3283) );
  OAI22_X1 U742 ( .A1(n4829), .A2(n6367), .B1(n512), .B2(n253), .ZN(n3284) );
  OAI22_X1 U743 ( .A1(n4797), .A2(n6364), .B1(n512), .B2(n255), .ZN(n3285) );
  OAI22_X1 U744 ( .A1(n4765), .A2(n6362), .B1(n512), .B2(n257), .ZN(n3286) );
  OAI22_X1 U745 ( .A1(n4733), .A2(n6361), .B1(n512), .B2(n259), .ZN(n3287) );
  OAI22_X1 U746 ( .A1(n4701), .A2(n6365), .B1(n512), .B2(n261), .ZN(n3288) );
  OAI22_X1 U747 ( .A1(n4669), .A2(n6366), .B1(n512), .B2(n263), .ZN(n3289) );
  OAI22_X1 U748 ( .A1(n4637), .A2(n6369), .B1(n512), .B2(n265), .ZN(n3290) );
  OAI22_X1 U749 ( .A1(n4605), .A2(n6370), .B1(n512), .B2(n267), .ZN(n3291) );
  OAI22_X1 U750 ( .A1(n4573), .A2(n6373), .B1(n512), .B2(n269), .ZN(n3292) );
  OAI22_X1 U751 ( .A1(n4541), .A2(n6374), .B1(n512), .B2(n271), .ZN(n3293) );
  OAI22_X1 U752 ( .A1(n4509), .A2(n6377), .B1(n512), .B2(n273), .ZN(n3294) );
  OAI22_X1 U753 ( .A1(n4477), .A2(n6378), .B1(n512), .B2(n275), .ZN(n3295) );
  OAI22_X1 U754 ( .A1(n4445), .A2(n6381), .B1(n512), .B2(n277), .ZN(n3296) );
  OAI22_X1 U755 ( .A1(n4413), .A2(n6384), .B1(n512), .B2(n279), .ZN(n3297) );
  OAI22_X1 U756 ( .A1(n4381), .A2(n6383), .B1(n512), .B2(n281), .ZN(n3298) );
  OAI22_X1 U757 ( .A1(n4349), .A2(n6391), .B1(n512), .B2(n283), .ZN(n3299) );
  OAI22_X1 U759 ( .A1(n501), .A2(n5677), .B1(n5414), .B2(n5623), .ZN(n525) );
  INV_X1 U760 ( .A(n5676), .ZN(n524) );
  OAI22_X1 U761 ( .A1(n5414), .A2(\UUT/Mcontrol/N22 ), .B1(n511), .B2(n7396), 
        .ZN(n3300) );
  INV_X1 U762 ( .A(n522), .ZN(n511) );
  OAI211_X1 U763 ( .C1(n6084), .C2(n287), .A(n526), .B(n527), .ZN(n522) );
  AOI222_X1 U764 ( .A1(\UUT/Mpath/the_mult/x_mult_out[14] ), .A2(n6357), .B1(
        n320), .B2(n528), .C1(n291), .C2(n529), .ZN(n527) );
  INV_X1 U765 ( .A(n5617), .ZN(n529) );
  AOI22_X1 U767 ( .A1(n6397), .A2(n530), .B1(n324), .B2(n6123), .ZN(n526) );
  INV_X1 U768 ( .A(n5579), .ZN(n530) );
  OAI221_X1 U769 ( .B1(n531), .B2(n80), .C1(n61), .C2(n81), .A(n532), .ZN(
        n3301) );
  NAND2_X1 U770 ( .A1(n7006), .A2(n6340), .ZN(n532) );
  AOI222_X1 U772 ( .A1(\UUT/jar_in [13]), .A2(n299), .B1(n300), .B2(
        \UUT/branch_rega [13]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [13]), 
        .C2(n301), .ZN(n533) );
  OAI222_X1 U773 ( .A1(n61), .A2(n94), .B1(n531), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N58 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3303) );
  INV_X1 U774 ( .A(\UUT/break_code[13] ), .ZN(n531) );
  INV_X1 U775 ( .A(n534), .ZN(n61) );
  OAI222_X1 U776 ( .A1(n535), .A2(n99), .B1(n536), .B2(n101), .C1(n5416), .C2(
        n102), .ZN(n534) );
  OAI221_X1 U777 ( .B1(n103), .B2(n537), .C1(n5618), .C2(n105), .A(n538), .ZN(
        n3304) );
  AOI22_X1 U778 ( .A1(n107), .A2(n539), .B1(\UUT/Mpath/the_mult/Mad_out [45]), 
        .B2(n109), .ZN(n538) );
  OAI221_X1 U779 ( .B1(n115), .B2(n540), .C1(n5581), .C2(n117), .A(n541), .ZN(
        n3305) );
  AOI22_X1 U780 ( .A1(n119), .A2(n539), .B1(\UUT/Mpath/the_mult/Mad_out [13]), 
        .B2(n121), .ZN(n541) );
  OAI22_X1 U782 ( .A1(n7385), .A2(n542), .B1(n5582), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3306) );
  OAI221_X1 U783 ( .B1(n543), .B2(n124), .C1(n125), .C2(n542), .A(n544), .ZN(
        n3307) );
  AOI22_X1 U784 ( .A1(n127), .A2(n545), .B1(n129), .B2(n546), .ZN(n544) );
  INV_X1 U785 ( .A(\UUT/Mpath/the_mult/x_operand1[13] ), .ZN(n542) );
  OAI221_X1 U786 ( .B1(n543), .B2(n218), .C1(\UUT/Mpath/the_alu/N57 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n547), .ZN(n3308) );
  AOI22_X1 U787 ( .A1(n220), .A2(n545), .B1(n221), .B2(n546), .ZN(n547) );
  INV_X1 U788 ( .A(n536), .ZN(n545) );
  OAI22_X1 U789 ( .A1(n5310), .A2(n6393), .B1(n536), .B2(n223), .ZN(n3309) );
  OAI22_X1 U790 ( .A1(n5278), .A2(n6396), .B1(n536), .B2(n225), .ZN(n3310) );
  OAI22_X1 U791 ( .A1(n5246), .A2(n6387), .B1(n536), .B2(n227), .ZN(n3311) );
  OAI22_X1 U792 ( .A1(n5214), .A2(n6395), .B1(n536), .B2(n229), .ZN(n3312) );
  OAI22_X1 U793 ( .A1(n5182), .A2(n6390), .B1(n536), .B2(n231), .ZN(n3313) );
  OAI22_X1 U794 ( .A1(n5150), .A2(n6385), .B1(n536), .B2(n233), .ZN(n3314) );
  OAI22_X1 U795 ( .A1(n5118), .A2(n6389), .B1(n536), .B2(n235), .ZN(n3315) );
  OAI22_X1 U796 ( .A1(n5086), .A2(n6382), .B1(n536), .B2(n237), .ZN(n3316) );
  OAI22_X1 U797 ( .A1(n5054), .A2(n6380), .B1(n536), .B2(n239), .ZN(n3317) );
  OAI22_X1 U798 ( .A1(n5022), .A2(n6379), .B1(n536), .B2(n241), .ZN(n3318) );
  OAI22_X1 U799 ( .A1(n4990), .A2(n6376), .B1(n536), .B2(n243), .ZN(n3319) );
  OAI22_X1 U800 ( .A1(n4958), .A2(n6375), .B1(n536), .B2(n245), .ZN(n3320) );
  OAI22_X1 U801 ( .A1(n4926), .A2(n6372), .B1(n536), .B2(n247), .ZN(n3321) );
  OAI22_X1 U802 ( .A1(n4894), .A2(n6371), .B1(n536), .B2(n249), .ZN(n3322) );
  OAI22_X1 U803 ( .A1(n4862), .A2(n6368), .B1(n536), .B2(n251), .ZN(n3323) );
  OAI22_X1 U804 ( .A1(n4830), .A2(n6367), .B1(n536), .B2(n253), .ZN(n3324) );
  OAI22_X1 U805 ( .A1(n4798), .A2(n6364), .B1(n536), .B2(n255), .ZN(n3325) );
  OAI22_X1 U806 ( .A1(n4766), .A2(n6362), .B1(n536), .B2(n257), .ZN(n3326) );
  OAI22_X1 U807 ( .A1(n4734), .A2(n6361), .B1(n536), .B2(n259), .ZN(n3327) );
  OAI22_X1 U808 ( .A1(n4702), .A2(n6365), .B1(n536), .B2(n261), .ZN(n3328) );
  OAI22_X1 U809 ( .A1(n4670), .A2(n6366), .B1(n536), .B2(n263), .ZN(n3329) );
  OAI22_X1 U810 ( .A1(n4638), .A2(n6369), .B1(n536), .B2(n265), .ZN(n3330) );
  OAI22_X1 U811 ( .A1(n4606), .A2(n6370), .B1(n536), .B2(n267), .ZN(n3331) );
  OAI22_X1 U812 ( .A1(n4574), .A2(n6373), .B1(n536), .B2(n269), .ZN(n3332) );
  OAI22_X1 U813 ( .A1(n4542), .A2(n6374), .B1(n536), .B2(n271), .ZN(n3333) );
  OAI22_X1 U814 ( .A1(n4510), .A2(n6377), .B1(n536), .B2(n273), .ZN(n3334) );
  OAI22_X1 U815 ( .A1(n4478), .A2(n6378), .B1(n536), .B2(n275), .ZN(n3335) );
  OAI22_X1 U816 ( .A1(n4446), .A2(n6381), .B1(n536), .B2(n277), .ZN(n3336) );
  OAI22_X1 U817 ( .A1(n4414), .A2(n6384), .B1(n536), .B2(n279), .ZN(n3337) );
  OAI22_X1 U818 ( .A1(n4382), .A2(n6383), .B1(n536), .B2(n281), .ZN(n3338) );
  OAI22_X1 U819 ( .A1(n4350), .A2(n6391), .B1(n536), .B2(n283), .ZN(n3339) );
  OAI22_X1 U821 ( .A1(n501), .A2(n5687), .B1(n5417), .B2(n5623), .ZN(n549) );
  INV_X1 U822 ( .A(n5686), .ZN(n548) );
  OAI22_X1 U823 ( .A1(n5417), .A2(\UUT/Mcontrol/N22 ), .B1(n535), .B2(n7395), 
        .ZN(n3340) );
  INV_X1 U824 ( .A(n546), .ZN(n535) );
  OAI211_X1 U825 ( .C1(n6094), .C2(n287), .A(n550), .B(n551), .ZN(n546) );
  AOI222_X1 U826 ( .A1(\UUT/Mpath/the_mult/x_mult_out[13] ), .A2(n6357), .B1(
        n320), .B2(n552), .C1(n291), .C2(n553), .ZN(n551) );
  INV_X1 U827 ( .A(n5618), .ZN(n553) );
  AOI22_X1 U829 ( .A1(n6397), .A2(n554), .B1(n324), .B2(n6124), .ZN(n550) );
  INV_X1 U830 ( .A(n5581), .ZN(n554) );
  OAI22_X1 U831 ( .A1(n555), .A2(n556), .B1(n297), .B2(n2671), .ZN(n3341) );
  INV_X1 U832 ( .A(\UUT/Mcontrol/Program_counter/N28 ), .ZN(n555) );
  OAI221_X1 U833 ( .B1(n557), .B2(n80), .C1(n60), .C2(n81), .A(n558), .ZN(
        n3342) );
  NAND2_X1 U834 ( .A1(\UUT/Mpath/the_mult/x_operand2 [12]), .A2(n6340), .ZN(
        n558) );
  OAI222_X1 U835 ( .A1(n60), .A2(n94), .B1(n557), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N60 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3343) );
  INV_X1 U836 ( .A(\UUT/break_code[12] ), .ZN(n557) );
  INV_X1 U837 ( .A(n559), .ZN(n60) );
  OAI222_X1 U838 ( .A1(n560), .A2(n99), .B1(n561), .B2(n101), .C1(n5419), .C2(
        n102), .ZN(n559) );
  OAI221_X1 U839 ( .B1(n103), .B2(n562), .C1(n5619), .C2(n105), .A(n563), .ZN(
        n3344) );
  AOI22_X1 U840 ( .A1(n107), .A2(n564), .B1(\UUT/Mpath/the_mult/Mad_out [44]), 
        .B2(n109), .ZN(n563) );
  OAI221_X1 U841 ( .B1(n115), .B2(n565), .C1(n5583), .C2(n117), .A(n566), .ZN(
        n3345) );
  AOI22_X1 U842 ( .A1(n119), .A2(n564), .B1(\UUT/Mpath/the_mult/Mad_out [12]), 
        .B2(n121), .ZN(n566) );
  OAI22_X1 U844 ( .A1(n7385), .A2(n567), .B1(n5584), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3346) );
  OAI221_X1 U845 ( .B1(n568), .B2(n124), .C1(n125), .C2(n567), .A(n569), .ZN(
        n3347) );
  AOI22_X1 U846 ( .A1(n127), .A2(n570), .B1(n129), .B2(n571), .ZN(n569) );
  INV_X1 U847 ( .A(\UUT/Mpath/the_mult/x_operand1[12] ), .ZN(n567) );
  OAI221_X1 U848 ( .B1(n568), .B2(n218), .C1(\UUT/Mpath/the_alu/N59 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n572), .ZN(n3348) );
  AOI22_X1 U849 ( .A1(n220), .A2(n570), .B1(n221), .B2(n571), .ZN(n572) );
  INV_X1 U850 ( .A(n561), .ZN(n570) );
  OAI22_X1 U851 ( .A1(n5311), .A2(n6393), .B1(n561), .B2(n223), .ZN(n3349) );
  OAI22_X1 U852 ( .A1(n5279), .A2(n6396), .B1(n561), .B2(n225), .ZN(n3350) );
  OAI22_X1 U853 ( .A1(n5247), .A2(n6387), .B1(n561), .B2(n227), .ZN(n3351) );
  OAI22_X1 U854 ( .A1(n5215), .A2(n6395), .B1(n561), .B2(n229), .ZN(n3352) );
  OAI22_X1 U855 ( .A1(n5183), .A2(n6390), .B1(n561), .B2(n231), .ZN(n3353) );
  OAI22_X1 U856 ( .A1(n5151), .A2(n6385), .B1(n561), .B2(n233), .ZN(n3354) );
  OAI22_X1 U857 ( .A1(n5119), .A2(n6389), .B1(n561), .B2(n235), .ZN(n3355) );
  OAI22_X1 U858 ( .A1(n5087), .A2(n6382), .B1(n561), .B2(n237), .ZN(n3356) );
  OAI22_X1 U859 ( .A1(n5055), .A2(n6380), .B1(n561), .B2(n239), .ZN(n3357) );
  OAI22_X1 U860 ( .A1(n5023), .A2(n6379), .B1(n561), .B2(n241), .ZN(n3358) );
  OAI22_X1 U861 ( .A1(n4991), .A2(n6376), .B1(n561), .B2(n243), .ZN(n3359) );
  OAI22_X1 U862 ( .A1(n4959), .A2(n6375), .B1(n561), .B2(n245), .ZN(n3360) );
  OAI22_X1 U863 ( .A1(n4927), .A2(n6372), .B1(n561), .B2(n247), .ZN(n3361) );
  OAI22_X1 U864 ( .A1(n4895), .A2(n6371), .B1(n561), .B2(n249), .ZN(n3362) );
  OAI22_X1 U865 ( .A1(n4863), .A2(n6368), .B1(n561), .B2(n251), .ZN(n3363) );
  OAI22_X1 U866 ( .A1(n4831), .A2(n6367), .B1(n561), .B2(n253), .ZN(n3364) );
  OAI22_X1 U867 ( .A1(n4799), .A2(n6364), .B1(n561), .B2(n255), .ZN(n3365) );
  OAI22_X1 U868 ( .A1(n4767), .A2(n6362), .B1(n561), .B2(n257), .ZN(n3366) );
  OAI22_X1 U869 ( .A1(n4735), .A2(n6361), .B1(n561), .B2(n259), .ZN(n3367) );
  OAI22_X1 U870 ( .A1(n4703), .A2(n6365), .B1(n561), .B2(n261), .ZN(n3368) );
  OAI22_X1 U871 ( .A1(n4671), .A2(n6366), .B1(n561), .B2(n263), .ZN(n3369) );
  OAI22_X1 U872 ( .A1(n4639), .A2(n6369), .B1(n561), .B2(n265), .ZN(n3370) );
  OAI22_X1 U873 ( .A1(n4607), .A2(n6370), .B1(n561), .B2(n267), .ZN(n3371) );
  OAI22_X1 U874 ( .A1(n4575), .A2(n6373), .B1(n561), .B2(n269), .ZN(n3372) );
  OAI22_X1 U875 ( .A1(n4543), .A2(n6374), .B1(n561), .B2(n271), .ZN(n3373) );
  OAI22_X1 U876 ( .A1(n4511), .A2(n6377), .B1(n561), .B2(n273), .ZN(n3374) );
  OAI22_X1 U877 ( .A1(n4479), .A2(n6378), .B1(n561), .B2(n275), .ZN(n3375) );
  OAI22_X1 U878 ( .A1(n4447), .A2(n6381), .B1(n561), .B2(n277), .ZN(n3376) );
  OAI22_X1 U879 ( .A1(n4415), .A2(n6384), .B1(n561), .B2(n279), .ZN(n3377) );
  OAI22_X1 U880 ( .A1(n4383), .A2(n6383), .B1(n561), .B2(n281), .ZN(n3378) );
  OAI22_X1 U881 ( .A1(n4351), .A2(n6391), .B1(n561), .B2(n283), .ZN(n3379) );
  OAI22_X1 U883 ( .A1(n501), .A2(n5697), .B1(n5420), .B2(n5623), .ZN(n574) );
  INV_X1 U884 ( .A(n5696), .ZN(n573) );
  OAI22_X1 U885 ( .A1(n5420), .A2(\UUT/Mcontrol/N22 ), .B1(n560), .B2(n7395), 
        .ZN(n3380) );
  INV_X1 U886 ( .A(n571), .ZN(n560) );
  OAI211_X1 U887 ( .C1(n6125), .C2(n287), .A(n575), .B(n576), .ZN(n571) );
  AOI222_X1 U888 ( .A1(\UUT/Mpath/the_mult/x_mult_out[12] ), .A2(n6357), .B1(
        n320), .B2(n577), .C1(n291), .C2(n578), .ZN(n576) );
  INV_X1 U889 ( .A(n5619), .ZN(n578) );
  AOI22_X1 U891 ( .A1(n6397), .A2(n579), .B1(n324), .B2(n6126), .ZN(n575) );
  INV_X1 U892 ( .A(n5583), .ZN(n579) );
  OAI22_X1 U893 ( .A1(n580), .A2(n556), .B1(n297), .B2(n2674), .ZN(n3381) );
  INV_X1 U894 ( .A(\UUT/Mcontrol/Program_counter/N26 ), .ZN(n580) );
  OAI221_X1 U895 ( .B1(n581), .B2(n80), .C1(n59), .C2(n81), .A(n582), .ZN(
        n3382) );
  NAND2_X1 U896 ( .A1(n7058), .A2(n6340), .ZN(n582) );
  OAI222_X1 U897 ( .A1(n59), .A2(n94), .B1(n581), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N62 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3383) );
  INV_X1 U898 ( .A(\UUT/break_code[11] ), .ZN(n581) );
  INV_X1 U899 ( .A(n583), .ZN(n59) );
  OAI222_X1 U900 ( .A1(n584), .A2(n99), .B1(n585), .B2(n101), .C1(n5422), .C2(
        n102), .ZN(n583) );
  OAI221_X1 U901 ( .B1(n103), .B2(n586), .C1(n5620), .C2(n105), .A(n587), .ZN(
        n3384) );
  AOI22_X1 U902 ( .A1(n107), .A2(n588), .B1(\UUT/Mpath/the_mult/Mad_out [43]), 
        .B2(n109), .ZN(n587) );
  OAI221_X1 U903 ( .B1(n115), .B2(n589), .C1(n5585), .C2(n117), .A(n590), .ZN(
        n3385) );
  AOI22_X1 U904 ( .A1(n119), .A2(n588), .B1(\UUT/Mpath/the_mult/Mad_out [11]), 
        .B2(n121), .ZN(n590) );
  OAI22_X1 U906 ( .A1(n7385), .A2(n591), .B1(n5586), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3386) );
  OAI221_X1 U907 ( .B1(n592), .B2(n124), .C1(n125), .C2(n591), .A(n593), .ZN(
        n3387) );
  AOI22_X1 U908 ( .A1(n127), .A2(n594), .B1(n129), .B2(n595), .ZN(n593) );
  INV_X1 U909 ( .A(\UUT/Mpath/the_mult/x_operand1[11] ), .ZN(n591) );
  OAI221_X1 U910 ( .B1(n592), .B2(n218), .C1(\UUT/Mpath/the_alu/N61 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n596), .ZN(n3388) );
  AOI22_X1 U911 ( .A1(n220), .A2(n594), .B1(n221), .B2(n595), .ZN(n596) );
  INV_X1 U912 ( .A(n585), .ZN(n594) );
  OAI22_X1 U913 ( .A1(n5312), .A2(n6393), .B1(n585), .B2(n223), .ZN(n3389) );
  OAI22_X1 U914 ( .A1(n5280), .A2(n6396), .B1(n585), .B2(n225), .ZN(n3390) );
  OAI22_X1 U915 ( .A1(n5248), .A2(n6387), .B1(n585), .B2(n227), .ZN(n3391) );
  OAI22_X1 U916 ( .A1(n5216), .A2(n6395), .B1(n585), .B2(n229), .ZN(n3392) );
  OAI22_X1 U917 ( .A1(n5184), .A2(n6390), .B1(n585), .B2(n231), .ZN(n3393) );
  OAI22_X1 U918 ( .A1(n5152), .A2(n6385), .B1(n585), .B2(n233), .ZN(n3394) );
  OAI22_X1 U919 ( .A1(n5120), .A2(n6389), .B1(n585), .B2(n235), .ZN(n3395) );
  OAI22_X1 U920 ( .A1(n5088), .A2(n6382), .B1(n585), .B2(n237), .ZN(n3396) );
  OAI22_X1 U921 ( .A1(n5056), .A2(n6380), .B1(n585), .B2(n239), .ZN(n3397) );
  OAI22_X1 U922 ( .A1(n5024), .A2(n6379), .B1(n585), .B2(n241), .ZN(n3398) );
  OAI22_X1 U923 ( .A1(n4992), .A2(n6376), .B1(n585), .B2(n243), .ZN(n3399) );
  OAI22_X1 U924 ( .A1(n4960), .A2(n6375), .B1(n585), .B2(n245), .ZN(n3400) );
  OAI22_X1 U925 ( .A1(n4928), .A2(n6372), .B1(n585), .B2(n247), .ZN(n3401) );
  OAI22_X1 U926 ( .A1(n4896), .A2(n6371), .B1(n585), .B2(n249), .ZN(n3402) );
  OAI22_X1 U927 ( .A1(n4864), .A2(n6368), .B1(n585), .B2(n251), .ZN(n3403) );
  OAI22_X1 U928 ( .A1(n4832), .A2(n6367), .B1(n585), .B2(n253), .ZN(n3404) );
  OAI22_X1 U929 ( .A1(n4800), .A2(n6364), .B1(n585), .B2(n255), .ZN(n3405) );
  OAI22_X1 U930 ( .A1(n4768), .A2(n6362), .B1(n585), .B2(n257), .ZN(n3406) );
  OAI22_X1 U931 ( .A1(n4736), .A2(n6361), .B1(n585), .B2(n259), .ZN(n3407) );
  OAI22_X1 U932 ( .A1(n4704), .A2(n6365), .B1(n585), .B2(n261), .ZN(n3408) );
  OAI22_X1 U933 ( .A1(n4672), .A2(n6366), .B1(n585), .B2(n263), .ZN(n3409) );
  OAI22_X1 U934 ( .A1(n4640), .A2(n6369), .B1(n585), .B2(n265), .ZN(n3410) );
  OAI22_X1 U935 ( .A1(n4608), .A2(n6370), .B1(n585), .B2(n267), .ZN(n3411) );
  OAI22_X1 U936 ( .A1(n4576), .A2(n6373), .B1(n585), .B2(n269), .ZN(n3412) );
  OAI22_X1 U937 ( .A1(n4544), .A2(n6374), .B1(n585), .B2(n271), .ZN(n3413) );
  OAI22_X1 U938 ( .A1(n4512), .A2(n6377), .B1(n585), .B2(n273), .ZN(n3414) );
  OAI22_X1 U939 ( .A1(n4480), .A2(n6378), .B1(n585), .B2(n275), .ZN(n3415) );
  OAI22_X1 U940 ( .A1(n4448), .A2(n6381), .B1(n585), .B2(n277), .ZN(n3416) );
  OAI22_X1 U941 ( .A1(n4416), .A2(n6384), .B1(n585), .B2(n279), .ZN(n3417) );
  OAI22_X1 U942 ( .A1(n4384), .A2(n6383), .B1(n585), .B2(n281), .ZN(n3418) );
  OAI22_X1 U943 ( .A1(n4352), .A2(n6391), .B1(n585), .B2(n283), .ZN(n3419) );
  OAI22_X1 U945 ( .A1(n501), .A2(n5707), .B1(n5423), .B2(n5623), .ZN(n598) );
  INV_X1 U946 ( .A(n5706), .ZN(n597) );
  OAI22_X1 U947 ( .A1(n5423), .A2(\UUT/Mcontrol/N22 ), .B1(n584), .B2(n7395), 
        .ZN(n3420) );
  INV_X1 U948 ( .A(n595), .ZN(n584) );
  OAI211_X1 U949 ( .C1(n6127), .C2(n287), .A(n599), .B(n600), .ZN(n595) );
  AOI222_X1 U950 ( .A1(\UUT/Mpath/the_mult/x_mult_out[11] ), .A2(n6357), .B1(
        n320), .B2(n601), .C1(n291), .C2(n602), .ZN(n600) );
  INV_X1 U951 ( .A(n5620), .ZN(n602) );
  AOI22_X1 U953 ( .A1(n6397), .A2(n603), .B1(n324), .B2(n6128), .ZN(n599) );
  INV_X1 U954 ( .A(n5585), .ZN(n603) );
  OAI221_X1 U955 ( .B1(n604), .B2(n80), .C1(n58), .C2(n81), .A(n605), .ZN(
        n3421) );
  NAND2_X1 U956 ( .A1(\UUT/Mpath/the_mult/x_operand2 [10]), .A2(n6340), .ZN(
        n605) );
  OAI222_X1 U957 ( .A1(n58), .A2(n94), .B1(n604), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N64 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3422) );
  INV_X1 U958 ( .A(\UUT/break_code[10] ), .ZN(n604) );
  INV_X1 U959 ( .A(n606), .ZN(n58) );
  OAI222_X1 U960 ( .A1(n607), .A2(n5332), .B1(n608), .B2(n101), .C1(n5425), 
        .C2(n102), .ZN(n606) );
  OAI221_X1 U961 ( .B1(n103), .B2(n609), .C1(n5621), .C2(n105), .A(n610), .ZN(
        n3423) );
  AOI22_X1 U962 ( .A1(n107), .A2(n611), .B1(\UUT/Mpath/the_mult/Mad_out [42]), 
        .B2(n109), .ZN(n610) );
  OAI221_X1 U963 ( .B1(n115), .B2(n612), .C1(n5587), .C2(n117), .A(n613), .ZN(
        n3424) );
  AOI22_X1 U964 ( .A1(n119), .A2(n611), .B1(\UUT/Mpath/the_mult/Mad_out [10]), 
        .B2(n121), .ZN(n613) );
  OAI22_X1 U966 ( .A1(n7386), .A2(n614), .B1(n5588), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3425) );
  OAI221_X1 U967 ( .B1(n615), .B2(n124), .C1(n125), .C2(n614), .A(n616), .ZN(
        n3426) );
  AOI22_X1 U968 ( .A1(n127), .A2(n617), .B1(n129), .B2(n618), .ZN(n616) );
  INV_X1 U969 ( .A(\UUT/Mpath/the_mult/x_operand1[10] ), .ZN(n614) );
  OAI221_X1 U970 ( .B1(n615), .B2(n218), .C1(\UUT/Mpath/the_alu/N63 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n619), .ZN(n3427) );
  AOI22_X1 U971 ( .A1(n220), .A2(n617), .B1(n221), .B2(n618), .ZN(n619) );
  INV_X1 U972 ( .A(n608), .ZN(n617) );
  OAI22_X1 U973 ( .A1(n5313), .A2(n6393), .B1(n608), .B2(n223), .ZN(n3428) );
  OAI22_X1 U974 ( .A1(n5281), .A2(n6396), .B1(n608), .B2(n225), .ZN(n3429) );
  OAI22_X1 U975 ( .A1(n5249), .A2(n6387), .B1(n608), .B2(n227), .ZN(n3430) );
  OAI22_X1 U976 ( .A1(n5217), .A2(n6395), .B1(n608), .B2(n229), .ZN(n3431) );
  OAI22_X1 U977 ( .A1(n5185), .A2(n6390), .B1(n608), .B2(n231), .ZN(n3432) );
  OAI22_X1 U978 ( .A1(n5153), .A2(n6385), .B1(n608), .B2(n233), .ZN(n3433) );
  OAI22_X1 U979 ( .A1(n5121), .A2(n6389), .B1(n608), .B2(n235), .ZN(n3434) );
  OAI22_X1 U980 ( .A1(n5089), .A2(n6382), .B1(n608), .B2(n237), .ZN(n3435) );
  OAI22_X1 U981 ( .A1(n5057), .A2(n6380), .B1(n608), .B2(n239), .ZN(n3436) );
  OAI22_X1 U982 ( .A1(n5025), .A2(n6379), .B1(n608), .B2(n241), .ZN(n3437) );
  OAI22_X1 U983 ( .A1(n4993), .A2(n6376), .B1(n608), .B2(n243), .ZN(n3438) );
  OAI22_X1 U984 ( .A1(n4961), .A2(n6375), .B1(n608), .B2(n245), .ZN(n3439) );
  OAI22_X1 U985 ( .A1(n4929), .A2(n6372), .B1(n608), .B2(n247), .ZN(n3440) );
  OAI22_X1 U986 ( .A1(n4897), .A2(n6371), .B1(n608), .B2(n249), .ZN(n3441) );
  OAI22_X1 U987 ( .A1(n4865), .A2(n6368), .B1(n608), .B2(n251), .ZN(n3442) );
  OAI22_X1 U988 ( .A1(n4833), .A2(n6367), .B1(n608), .B2(n253), .ZN(n3443) );
  OAI22_X1 U989 ( .A1(n4801), .A2(n6364), .B1(n608), .B2(n255), .ZN(n3444) );
  OAI22_X1 U990 ( .A1(n4769), .A2(n6362), .B1(n608), .B2(n257), .ZN(n3445) );
  OAI22_X1 U991 ( .A1(n4737), .A2(n6361), .B1(n608), .B2(n259), .ZN(n3446) );
  OAI22_X1 U992 ( .A1(n4705), .A2(n6365), .B1(n608), .B2(n261), .ZN(n3447) );
  OAI22_X1 U993 ( .A1(n4673), .A2(n6366), .B1(n608), .B2(n263), .ZN(n3448) );
  OAI22_X1 U994 ( .A1(n4641), .A2(n6369), .B1(n608), .B2(n265), .ZN(n3449) );
  OAI22_X1 U995 ( .A1(n4609), .A2(n6370), .B1(n608), .B2(n267), .ZN(n3450) );
  OAI22_X1 U996 ( .A1(n4577), .A2(n6373), .B1(n608), .B2(n269), .ZN(n3451) );
  OAI22_X1 U997 ( .A1(n4545), .A2(n6374), .B1(n608), .B2(n271), .ZN(n3452) );
  OAI22_X1 U998 ( .A1(n4513), .A2(n6377), .B1(n608), .B2(n273), .ZN(n3453) );
  OAI22_X1 U999 ( .A1(n4481), .A2(n6378), .B1(n608), .B2(n275), .ZN(n3454) );
  OAI22_X1 U1000 ( .A1(n4449), .A2(n6381), .B1(n608), .B2(n277), .ZN(n3455) );
  OAI22_X1 U1001 ( .A1(n4417), .A2(n6384), .B1(n608), .B2(n279), .ZN(n3456) );
  OAI22_X1 U1002 ( .A1(n4385), .A2(n6383), .B1(n608), .B2(n281), .ZN(n3457) );
  OAI22_X1 U1003 ( .A1(n4353), .A2(n6391), .B1(n608), .B2(n283), .ZN(n3458) );
  OAI22_X1 U1005 ( .A1(n501), .A2(n5728), .B1(n5426), .B2(n5623), .ZN(n621) );
  INV_X1 U1006 ( .A(n5727), .ZN(n620) );
  OAI22_X1 U1007 ( .A1(n5426), .A2(\UUT/Mcontrol/N22 ), .B1(n607), .B2(n7395), 
        .ZN(n3459) );
  INV_X1 U1008 ( .A(n618), .ZN(n607) );
  OAI211_X1 U1009 ( .C1(n6129), .C2(n287), .A(n622), .B(n623), .ZN(n618) );
  AOI222_X1 U1010 ( .A1(\UUT/Mpath/the_mult/x_mult_out[10] ), .A2(n6357), .B1(
        n320), .B2(n624), .C1(n291), .C2(n625), .ZN(n623) );
  INV_X1 U1011 ( .A(n5621), .ZN(n625) );
  AOI22_X1 U1013 ( .A1(n6397), .A2(n626), .B1(n324), .B2(n6130), .ZN(n622) );
  INV_X1 U1014 ( .A(n5587), .ZN(n626) );
  OAI221_X1 U1015 ( .B1(n627), .B2(n80), .C1(n57), .C2(n81), .A(n628), .ZN(
        n3460) );
  NAND2_X1 U1016 ( .A1(n7032), .A2(n6340), .ZN(n628) );
  OAI222_X1 U1017 ( .A1(n57), .A2(n94), .B1(n627), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N66 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3461) );
  INV_X1 U1018 ( .A(\UUT/break_code[9] ), .ZN(n627) );
  INV_X1 U1019 ( .A(n629), .ZN(n57) );
  OAI222_X1 U1020 ( .A1(n630), .A2(n99), .B1(n631), .B2(n101), .C1(n5333), 
        .C2(n102), .ZN(n629) );
  OAI221_X1 U1021 ( .B1(n103), .B2(n632), .C1(n5591), .C2(n105), .A(n633), 
        .ZN(n3462) );
  AOI22_X1 U1022 ( .A1(n107), .A2(n634), .B1(\UUT/Mpath/the_mult/Mad_out [41]), 
        .B2(n109), .ZN(n633) );
  OAI221_X1 U1023 ( .B1(n115), .B2(n635), .C1(n5527), .C2(n117), .A(n636), 
        .ZN(n3463) );
  AOI22_X1 U1024 ( .A1(n119), .A2(n634), .B1(\UUT/Mpath/the_mult/Mad_out [9]), 
        .B2(n121), .ZN(n636) );
  OAI22_X1 U1026 ( .A1(n7383), .A2(n637), .B1(n5528), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3464) );
  OAI221_X1 U1027 ( .B1(n638), .B2(n124), .C1(n125), .C2(n637), .A(n639), .ZN(
        n3465) );
  AOI22_X1 U1028 ( .A1(n127), .A2(n640), .B1(n129), .B2(n641), .ZN(n639) );
  INV_X1 U1029 ( .A(\UUT/Mpath/the_mult/x_operand1[9] ), .ZN(n637) );
  OAI221_X1 U1030 ( .B1(n638), .B2(n218), .C1(\UUT/Mpath/the_alu/N65 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n642), .ZN(n3466) );
  AOI22_X1 U1031 ( .A1(n220), .A2(n640), .B1(n221), .B2(n641), .ZN(n642) );
  INV_X1 U1032 ( .A(n631), .ZN(n640) );
  OAI22_X1 U1033 ( .A1(n5283), .A2(n6393), .B1(n631), .B2(n223), .ZN(n3467) );
  OAI22_X1 U1034 ( .A1(n5251), .A2(n6396), .B1(n631), .B2(n225), .ZN(n3468) );
  OAI22_X1 U1035 ( .A1(n5219), .A2(n6387), .B1(n631), .B2(n227), .ZN(n3469) );
  OAI22_X1 U1036 ( .A1(n5187), .A2(n6395), .B1(n631), .B2(n229), .ZN(n3470) );
  OAI22_X1 U1037 ( .A1(n5155), .A2(n6390), .B1(n631), .B2(n231), .ZN(n3471) );
  OAI22_X1 U1038 ( .A1(n5123), .A2(n6385), .B1(n631), .B2(n233), .ZN(n3472) );
  OAI22_X1 U1039 ( .A1(n5091), .A2(n6389), .B1(n631), .B2(n235), .ZN(n3473) );
  OAI22_X1 U1040 ( .A1(n5059), .A2(n6382), .B1(n631), .B2(n237), .ZN(n3474) );
  OAI22_X1 U1041 ( .A1(n5027), .A2(n6380), .B1(n631), .B2(n239), .ZN(n3475) );
  OAI22_X1 U1042 ( .A1(n4995), .A2(n6379), .B1(n631), .B2(n241), .ZN(n3476) );
  OAI22_X1 U1043 ( .A1(n4963), .A2(n6376), .B1(n631), .B2(n243), .ZN(n3477) );
  OAI22_X1 U1044 ( .A1(n4931), .A2(n6375), .B1(n631), .B2(n245), .ZN(n3478) );
  OAI22_X1 U1045 ( .A1(n4899), .A2(n6372), .B1(n631), .B2(n247), .ZN(n3479) );
  OAI22_X1 U1046 ( .A1(n4867), .A2(n6371), .B1(n631), .B2(n249), .ZN(n3480) );
  OAI22_X1 U1047 ( .A1(n4835), .A2(n6368), .B1(n631), .B2(n251), .ZN(n3481) );
  OAI22_X1 U1048 ( .A1(n4803), .A2(n6367), .B1(n631), .B2(n253), .ZN(n3482) );
  OAI22_X1 U1049 ( .A1(n4771), .A2(n6364), .B1(n631), .B2(n255), .ZN(n3483) );
  OAI22_X1 U1050 ( .A1(n4739), .A2(n6362), .B1(n631), .B2(n257), .ZN(n3484) );
  OAI22_X1 U1051 ( .A1(n4707), .A2(n6361), .B1(n631), .B2(n259), .ZN(n3485) );
  OAI22_X1 U1052 ( .A1(n4675), .A2(n6365), .B1(n631), .B2(n261), .ZN(n3486) );
  OAI22_X1 U1053 ( .A1(n4643), .A2(n6366), .B1(n631), .B2(n263), .ZN(n3487) );
  OAI22_X1 U1054 ( .A1(n4611), .A2(n6369), .B1(n631), .B2(n265), .ZN(n3488) );
  OAI22_X1 U1055 ( .A1(n4579), .A2(n6370), .B1(n631), .B2(n267), .ZN(n3489) );
  OAI22_X1 U1056 ( .A1(n4547), .A2(n6373), .B1(n631), .B2(n269), .ZN(n3490) );
  OAI22_X1 U1057 ( .A1(n4515), .A2(n6374), .B1(n631), .B2(n271), .ZN(n3491) );
  OAI22_X1 U1058 ( .A1(n4483), .A2(n6377), .B1(n631), .B2(n273), .ZN(n3492) );
  OAI22_X1 U1059 ( .A1(n4451), .A2(n6378), .B1(n631), .B2(n275), .ZN(n3493) );
  OAI22_X1 U1060 ( .A1(n4419), .A2(n6381), .B1(n631), .B2(n277), .ZN(n3494) );
  OAI22_X1 U1061 ( .A1(n4387), .A2(n6384), .B1(n631), .B2(n279), .ZN(n3495) );
  OAI22_X1 U1062 ( .A1(n4355), .A2(n6383), .B1(n631), .B2(n281), .ZN(n3496) );
  OAI22_X1 U1063 ( .A1(n4323), .A2(n6391), .B1(n631), .B2(n283), .ZN(n3497) );
  OAI22_X1 U1065 ( .A1(n501), .A2(n5799), .B1(n5335), .B2(n5623), .ZN(n644) );
  OAI22_X1 U1066 ( .A1(n5335), .A2(\UUT/Mcontrol/N22 ), .B1(n630), .B2(n7395), 
        .ZN(n3498) );
  INV_X1 U1067 ( .A(n641), .ZN(n630) );
  OAI211_X1 U1068 ( .C1(n6096), .C2(n287), .A(n645), .B(n646), .ZN(n641) );
  AOI222_X1 U1069 ( .A1(\UUT/Mpath/the_mult/x_mult_out[9] ), .A2(n6357), .B1(
        n320), .B2(n647), .C1(n291), .C2(n648), .ZN(n646) );
  INV_X1 U1070 ( .A(n5591), .ZN(n648) );
  AOI22_X1 U1072 ( .A1(n6397), .A2(n649), .B1(n324), .B2(n6097), .ZN(n645) );
  INV_X1 U1073 ( .A(n5527), .ZN(n649) );
  OAI22_X1 U1074 ( .A1(n650), .A2(n556), .B1(n297), .B2(n2681), .ZN(n3499) );
  INV_X1 U1075 ( .A(\UUT/Mcontrol/Program_counter/N20 ), .ZN(n650) );
  OAI221_X1 U1076 ( .B1(n651), .B2(n80), .C1(n56), .C2(n81), .A(n652), .ZN(
        n3500) );
  NAND2_X1 U1077 ( .A1(\UUT/Mpath/the_mult/x_operand2 [8]), .A2(n6340), .ZN(
        n652) );
  OAI222_X1 U1078 ( .A1(n56), .A2(n94), .B1(n651), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N68 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3501) );
  INV_X1 U1079 ( .A(\UUT/break_code[8] ), .ZN(n651) );
  INV_X1 U1080 ( .A(n653), .ZN(n56) );
  OAI222_X1 U1081 ( .A1(n654), .A2(n5332), .B1(n655), .B2(n101), .C1(n5338), 
        .C2(n102), .ZN(n653) );
  OAI221_X1 U1082 ( .B1(n103), .B2(n656), .C1(n5592), .C2(n105), .A(n657), 
        .ZN(n3502) );
  AOI22_X1 U1083 ( .A1(n107), .A2(n658), .B1(\UUT/Mpath/the_mult/Mad_out [40]), 
        .B2(n109), .ZN(n657) );
  OAI221_X1 U1084 ( .B1(n115), .B2(n659), .C1(n5529), .C2(n117), .A(n660), 
        .ZN(n3503) );
  AOI22_X1 U1085 ( .A1(n119), .A2(n658), .B1(\UUT/Mpath/the_mult/Mad_out [8]), 
        .B2(n121), .ZN(n660) );
  OAI22_X1 U1087 ( .A1(n7383), .A2(n661), .B1(n5530), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3504) );
  OAI221_X1 U1088 ( .B1(n662), .B2(n124), .C1(n125), .C2(n661), .A(n663), .ZN(
        n3505) );
  AOI22_X1 U1089 ( .A1(n127), .A2(n664), .B1(n129), .B2(n665), .ZN(n663) );
  INV_X1 U1090 ( .A(\UUT/Mpath/the_mult/x_operand1[8] ), .ZN(n661) );
  OAI221_X1 U1091 ( .B1(n662), .B2(n218), .C1(\UUT/Mpath/the_alu/N67 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n666), .ZN(n3506) );
  AOI22_X1 U1092 ( .A1(n220), .A2(n664), .B1(n221), .B2(n665), .ZN(n666) );
  INV_X1 U1093 ( .A(n655), .ZN(n664) );
  OAI22_X1 U1094 ( .A1(n5284), .A2(n6393), .B1(n655), .B2(n223), .ZN(n3507) );
  OAI22_X1 U1095 ( .A1(n5252), .A2(n6396), .B1(n655), .B2(n225), .ZN(n3508) );
  OAI22_X1 U1096 ( .A1(n5220), .A2(n6387), .B1(n655), .B2(n227), .ZN(n3509) );
  OAI22_X1 U1097 ( .A1(n5188), .A2(n6395), .B1(n655), .B2(n229), .ZN(n3510) );
  OAI22_X1 U1098 ( .A1(n5156), .A2(n6390), .B1(n655), .B2(n231), .ZN(n3511) );
  OAI22_X1 U1099 ( .A1(n5124), .A2(n6385), .B1(n655), .B2(n233), .ZN(n3512) );
  OAI22_X1 U1100 ( .A1(n5092), .A2(n6389), .B1(n655), .B2(n235), .ZN(n3513) );
  OAI22_X1 U1101 ( .A1(n5060), .A2(n6382), .B1(n655), .B2(n237), .ZN(n3514) );
  OAI22_X1 U1102 ( .A1(n5028), .A2(n6380), .B1(n655), .B2(n239), .ZN(n3515) );
  OAI22_X1 U1103 ( .A1(n4996), .A2(n6379), .B1(n655), .B2(n241), .ZN(n3516) );
  OAI22_X1 U1104 ( .A1(n4964), .A2(n6376), .B1(n655), .B2(n243), .ZN(n3517) );
  OAI22_X1 U1105 ( .A1(n4932), .A2(n6375), .B1(n655), .B2(n245), .ZN(n3518) );
  OAI22_X1 U1106 ( .A1(n4900), .A2(n6372), .B1(n655), .B2(n247), .ZN(n3519) );
  OAI22_X1 U1107 ( .A1(n4868), .A2(n6371), .B1(n655), .B2(n249), .ZN(n3520) );
  OAI22_X1 U1108 ( .A1(n4836), .A2(n6368), .B1(n655), .B2(n251), .ZN(n3521) );
  OAI22_X1 U1109 ( .A1(n4804), .A2(n6367), .B1(n655), .B2(n253), .ZN(n3522) );
  OAI22_X1 U1110 ( .A1(n4772), .A2(n6364), .B1(n655), .B2(n255), .ZN(n3523) );
  OAI22_X1 U1111 ( .A1(n4740), .A2(n6362), .B1(n655), .B2(n257), .ZN(n3524) );
  OAI22_X1 U1112 ( .A1(n4708), .A2(n6361), .B1(n655), .B2(n259), .ZN(n3525) );
  OAI22_X1 U1113 ( .A1(n4676), .A2(n6365), .B1(n655), .B2(n261), .ZN(n3526) );
  OAI22_X1 U1114 ( .A1(n4644), .A2(n6366), .B1(n655), .B2(n263), .ZN(n3527) );
  OAI22_X1 U1115 ( .A1(n4612), .A2(n6369), .B1(n655), .B2(n265), .ZN(n3528) );
  OAI22_X1 U1116 ( .A1(n4580), .A2(n6370), .B1(n655), .B2(n267), .ZN(n3529) );
  OAI22_X1 U1117 ( .A1(n4548), .A2(n6373), .B1(n655), .B2(n269), .ZN(n3530) );
  OAI22_X1 U1118 ( .A1(n4516), .A2(n6374), .B1(n655), .B2(n271), .ZN(n3531) );
  OAI22_X1 U1119 ( .A1(n4484), .A2(n6377), .B1(n655), .B2(n273), .ZN(n3532) );
  OAI22_X1 U1120 ( .A1(n4452), .A2(n6378), .B1(n655), .B2(n275), .ZN(n3533) );
  OAI22_X1 U1121 ( .A1(n4420), .A2(n6381), .B1(n655), .B2(n277), .ZN(n3534) );
  OAI22_X1 U1122 ( .A1(n4388), .A2(n6384), .B1(n655), .B2(n279), .ZN(n3535) );
  OAI22_X1 U1123 ( .A1(n4356), .A2(n6383), .B1(n655), .B2(n281), .ZN(n3536) );
  OAI22_X1 U1124 ( .A1(n4324), .A2(n6391), .B1(n655), .B2(n283), .ZN(n3537) );
  OAI22_X1 U1126 ( .A1(n501), .A2(n5870), .B1(n5339), .B2(n5623), .ZN(n668) );
  NAND2_X1 U1127 ( .A1(n5624), .A2(n5623), .ZN(n501) );
  AND2_X1 U1128 ( .A1(n5625), .A2(n5623), .ZN(n498) );
  OAI22_X1 U1129 ( .A1(n5339), .A2(\UUT/Mcontrol/N22 ), .B1(n654), .B2(n7395), 
        .ZN(n3538) );
  INV_X1 U1130 ( .A(n665), .ZN(n654) );
  OAI211_X1 U1131 ( .C1(n6098), .C2(n287), .A(n669), .B(n670), .ZN(n665) );
  AOI222_X1 U1132 ( .A1(\UUT/Mpath/the_mult/x_mult_out[8] ), .A2(n6357), .B1(
        n320), .B2(n671), .C1(n291), .C2(n672), .ZN(n670) );
  INV_X1 U1133 ( .A(n5592), .ZN(n672) );
  AOI22_X1 U1135 ( .A1(n6397), .A2(n673), .B1(n324), .B2(n6099), .ZN(n669) );
  INV_X1 U1136 ( .A(n5529), .ZN(n673) );
  OAI22_X1 U1137 ( .A1(n674), .A2(n556), .B1(n297), .B2(n2684), .ZN(n3539) );
  INV_X1 U1138 ( .A(\UUT/Mcontrol/Program_counter/N18 ), .ZN(n674) );
  OAI221_X1 U1139 ( .B1(n675), .B2(n80), .C1(n55), .C2(n81), .A(n676), .ZN(
        n3540) );
  NAND2_X1 U1140 ( .A1(n6965), .A2(n6340), .ZN(n676) );
  OAI222_X1 U1141 ( .A1(n55), .A2(n94), .B1(n675), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N70 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3541) );
  INV_X1 U1142 ( .A(\UUT/break_code[7] ), .ZN(n675) );
  INV_X1 U1143 ( .A(n677), .ZN(n55) );
  OAI222_X1 U1144 ( .A1(n678), .A2(n99), .B1(n679), .B2(n101), .C1(n5341), 
        .C2(n102), .ZN(n677) );
  OAI221_X1 U1145 ( .B1(n103), .B2(n680), .C1(n5593), .C2(n105), .A(n681), 
        .ZN(n3542) );
  AOI22_X1 U1146 ( .A1(n107), .A2(n682), .B1(\UUT/Mpath/the_mult/Mad_out [39]), 
        .B2(n109), .ZN(n681) );
  OAI221_X1 U1147 ( .B1(n115), .B2(n683), .C1(n5531), .C2(n117), .A(n684), 
        .ZN(n3543) );
  AOI22_X1 U1148 ( .A1(n119), .A2(n682), .B1(\UUT/Mpath/the_mult/Mad_out [7]), 
        .B2(n121), .ZN(n684) );
  OAI22_X1 U1150 ( .A1(n7383), .A2(n685), .B1(n5532), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3544) );
  OAI221_X1 U1151 ( .B1(n686), .B2(n124), .C1(n125), .C2(n685), .A(n687), .ZN(
        n3545) );
  AOI22_X1 U1152 ( .A1(n127), .A2(n688), .B1(n129), .B2(n689), .ZN(n687) );
  INV_X1 U1153 ( .A(\UUT/Mpath/the_mult/x_operand1[7] ), .ZN(n685) );
  OAI221_X1 U1154 ( .B1(n686), .B2(n218), .C1(\UUT/Mpath/the_alu/N69 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n690), .ZN(n3546) );
  AOI22_X1 U1155 ( .A1(n220), .A2(n688), .B1(n221), .B2(n689), .ZN(n690) );
  OAI22_X1 U1156 ( .A1(n5285), .A2(n6393), .B1(n679), .B2(n223), .ZN(n3547) );
  OAI22_X1 U1157 ( .A1(n5253), .A2(n6396), .B1(n679), .B2(n225), .ZN(n3548) );
  OAI22_X1 U1158 ( .A1(n5221), .A2(n6387), .B1(n679), .B2(n227), .ZN(n3549) );
  OAI22_X1 U1159 ( .A1(n5189), .A2(n6395), .B1(n679), .B2(n229), .ZN(n3550) );
  OAI22_X1 U1160 ( .A1(n5157), .A2(n6390), .B1(n679), .B2(n231), .ZN(n3551) );
  OAI22_X1 U1161 ( .A1(n5125), .A2(n6385), .B1(n679), .B2(n233), .ZN(n3552) );
  OAI22_X1 U1162 ( .A1(n5093), .A2(n6389), .B1(n679), .B2(n235), .ZN(n3553) );
  OAI22_X1 U1163 ( .A1(n5061), .A2(n6382), .B1(n679), .B2(n237), .ZN(n3554) );
  OAI22_X1 U1164 ( .A1(n5029), .A2(n6380), .B1(n679), .B2(n239), .ZN(n3555) );
  OAI22_X1 U1165 ( .A1(n4997), .A2(n6379), .B1(n679), .B2(n241), .ZN(n3556) );
  OAI22_X1 U1166 ( .A1(n4965), .A2(n6376), .B1(n679), .B2(n243), .ZN(n3557) );
  OAI22_X1 U1167 ( .A1(n4933), .A2(n6375), .B1(n679), .B2(n245), .ZN(n3558) );
  OAI22_X1 U1168 ( .A1(n4901), .A2(n6372), .B1(n679), .B2(n247), .ZN(n3559) );
  OAI22_X1 U1169 ( .A1(n4869), .A2(n6371), .B1(n679), .B2(n249), .ZN(n3560) );
  OAI22_X1 U1170 ( .A1(n4837), .A2(n6368), .B1(n679), .B2(n251), .ZN(n3561) );
  OAI22_X1 U1171 ( .A1(n4805), .A2(n6367), .B1(n679), .B2(n253), .ZN(n3562) );
  OAI22_X1 U1172 ( .A1(n4773), .A2(n6364), .B1(n679), .B2(n255), .ZN(n3563) );
  OAI22_X1 U1173 ( .A1(n4741), .A2(n6362), .B1(n679), .B2(n257), .ZN(n3564) );
  OAI22_X1 U1174 ( .A1(n4709), .A2(n6361), .B1(n679), .B2(n259), .ZN(n3565) );
  OAI22_X1 U1175 ( .A1(n4677), .A2(n6365), .B1(n679), .B2(n261), .ZN(n3566) );
  OAI22_X1 U1176 ( .A1(n4645), .A2(n6366), .B1(n679), .B2(n263), .ZN(n3567) );
  OAI22_X1 U1177 ( .A1(n4613), .A2(n6369), .B1(n679), .B2(n265), .ZN(n3568) );
  OAI22_X1 U1178 ( .A1(n4581), .A2(n6370), .B1(n679), .B2(n267), .ZN(n3569) );
  OAI22_X1 U1179 ( .A1(n4549), .A2(n6373), .B1(n679), .B2(n269), .ZN(n3570) );
  OAI22_X1 U1180 ( .A1(n4517), .A2(n6374), .B1(n679), .B2(n271), .ZN(n3571) );
  OAI22_X1 U1181 ( .A1(n4485), .A2(n6377), .B1(n679), .B2(n273), .ZN(n3572) );
  OAI22_X1 U1182 ( .A1(n4453), .A2(n6378), .B1(n679), .B2(n275), .ZN(n3573) );
  OAI22_X1 U1183 ( .A1(n4421), .A2(n6381), .B1(n679), .B2(n277), .ZN(n3574) );
  OAI22_X1 U1184 ( .A1(n4389), .A2(n6384), .B1(n679), .B2(n279), .ZN(n3575) );
  OAI22_X1 U1185 ( .A1(n4357), .A2(n6383), .B1(n679), .B2(n281), .ZN(n3576) );
  OAI22_X1 U1186 ( .A1(n4325), .A2(n6391), .B1(n679), .B2(n283), .ZN(n3577) );
  OAI221_X1 U1188 ( .B1(n691), .B2(n692), .C1(n5623), .C2(n5342), .A(n693), 
        .ZN(n688) );
  AOI221_X1 U1189 ( .B1(D_DATA_INBUS[7]), .B2(n5663), .C1(D_DATA_INBUS[23]), 
        .C2(n5664), .A(n5665), .ZN(n691) );
  OAI22_X1 U1190 ( .A1(n5342), .A2(\UUT/Mcontrol/N22 ), .B1(n678), .B2(n7394), 
        .ZN(n3578) );
  INV_X1 U1191 ( .A(n689), .ZN(n678) );
  OAI211_X1 U1192 ( .C1(n6100), .C2(n287), .A(n694), .B(n695), .ZN(n689) );
  AOI222_X1 U1193 ( .A1(\UUT/Mpath/the_mult/x_mult_out[7] ), .A2(n6357), .B1(
        n320), .B2(n696), .C1(n291), .C2(n697), .ZN(n695) );
  INV_X1 U1194 ( .A(n5593), .ZN(n697) );
  AOI22_X1 U1196 ( .A1(n6397), .A2(n698), .B1(n324), .B2(n6101), .ZN(n694) );
  INV_X1 U1197 ( .A(n5531), .ZN(n698) );
  OAI22_X1 U1198 ( .A1(n699), .A2(n556), .B1(n297), .B2(n2687), .ZN(n3579) );
  INV_X1 U1199 ( .A(\UUT/Mcontrol/Program_counter/N16 ), .ZN(n699) );
  OAI221_X1 U1200 ( .B1(n700), .B2(n80), .C1(n54), .C2(n81), .A(n701), .ZN(
        n3580) );
  NAND2_X1 U1201 ( .A1(\UUT/Mpath/the_mult/x_operand2 [6]), .A2(n6340), .ZN(
        n701) );
  OAI222_X1 U1202 ( .A1(n54), .A2(n94), .B1(n700), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N72 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3581) );
  INV_X1 U1203 ( .A(\UUT/break_code[6] ), .ZN(n700) );
  INV_X1 U1204 ( .A(n702), .ZN(n54) );
  OAI222_X1 U1205 ( .A1(n703), .A2(n99), .B1(n704), .B2(n101), .C1(n5344), 
        .C2(n102), .ZN(n702) );
  OAI221_X1 U1206 ( .B1(n103), .B2(n705), .C1(n5594), .C2(n105), .A(n706), 
        .ZN(n3582) );
  AOI22_X1 U1207 ( .A1(n107), .A2(n707), .B1(\UUT/Mpath/the_mult/Mad_out [38]), 
        .B2(n109), .ZN(n706) );
  OAI221_X1 U1208 ( .B1(n115), .B2(n708), .C1(n5533), .C2(n117), .A(n709), 
        .ZN(n3583) );
  AOI22_X1 U1209 ( .A1(n119), .A2(n707), .B1(\UUT/Mpath/the_mult/Mad_out [6]), 
        .B2(n121), .ZN(n709) );
  OAI22_X1 U1211 ( .A1(n7383), .A2(n710), .B1(n5534), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3584) );
  OAI221_X1 U1212 ( .B1(n711), .B2(n124), .C1(n125), .C2(n710), .A(n712), .ZN(
        n3585) );
  AOI22_X1 U1213 ( .A1(n127), .A2(n713), .B1(n129), .B2(n714), .ZN(n712) );
  INV_X1 U1214 ( .A(\UUT/Mpath/the_mult/x_operand1[6] ), .ZN(n710) );
  OAI221_X1 U1215 ( .B1(n711), .B2(n218), .C1(\UUT/Mpath/the_alu/N71 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n715), .ZN(n3586) );
  AOI22_X1 U1216 ( .A1(n220), .A2(n713), .B1(n221), .B2(n714), .ZN(n715) );
  OAI22_X1 U1217 ( .A1(n5286), .A2(n6393), .B1(n704), .B2(n223), .ZN(n3587) );
  OAI22_X1 U1218 ( .A1(n5254), .A2(n6396), .B1(n704), .B2(n225), .ZN(n3588) );
  OAI22_X1 U1219 ( .A1(n5222), .A2(n6387), .B1(n704), .B2(n227), .ZN(n3589) );
  OAI22_X1 U1220 ( .A1(n5190), .A2(n6395), .B1(n704), .B2(n229), .ZN(n3590) );
  OAI22_X1 U1221 ( .A1(n5158), .A2(n6390), .B1(n704), .B2(n231), .ZN(n3591) );
  OAI22_X1 U1222 ( .A1(n5126), .A2(n6385), .B1(n704), .B2(n233), .ZN(n3592) );
  OAI22_X1 U1223 ( .A1(n5094), .A2(n6389), .B1(n704), .B2(n235), .ZN(n3593) );
  OAI22_X1 U1224 ( .A1(n5062), .A2(n6382), .B1(n704), .B2(n237), .ZN(n3594) );
  OAI22_X1 U1225 ( .A1(n5030), .A2(n6380), .B1(n704), .B2(n239), .ZN(n3595) );
  OAI22_X1 U1226 ( .A1(n4998), .A2(n6379), .B1(n704), .B2(n241), .ZN(n3596) );
  OAI22_X1 U1227 ( .A1(n4966), .A2(n6376), .B1(n704), .B2(n243), .ZN(n3597) );
  OAI22_X1 U1228 ( .A1(n4934), .A2(n6375), .B1(n704), .B2(n245), .ZN(n3598) );
  OAI22_X1 U1229 ( .A1(n4902), .A2(n6372), .B1(n704), .B2(n247), .ZN(n3599) );
  OAI22_X1 U1230 ( .A1(n4870), .A2(n6371), .B1(n704), .B2(n249), .ZN(n3600) );
  OAI22_X1 U1231 ( .A1(n4838), .A2(n6368), .B1(n704), .B2(n251), .ZN(n3601) );
  OAI22_X1 U1232 ( .A1(n4806), .A2(n6367), .B1(n704), .B2(n253), .ZN(n3602) );
  OAI22_X1 U1233 ( .A1(n4774), .A2(n6364), .B1(n704), .B2(n255), .ZN(n3603) );
  OAI22_X1 U1234 ( .A1(n4742), .A2(n6362), .B1(n704), .B2(n257), .ZN(n3604) );
  OAI22_X1 U1235 ( .A1(n4710), .A2(n6361), .B1(n704), .B2(n259), .ZN(n3605) );
  OAI22_X1 U1236 ( .A1(n4678), .A2(n6365), .B1(n704), .B2(n261), .ZN(n3606) );
  OAI22_X1 U1237 ( .A1(n4646), .A2(n6366), .B1(n704), .B2(n263), .ZN(n3607) );
  OAI22_X1 U1238 ( .A1(n4614), .A2(n6369), .B1(n704), .B2(n265), .ZN(n3608) );
  OAI22_X1 U1239 ( .A1(n4582), .A2(n6370), .B1(n704), .B2(n267), .ZN(n3609) );
  OAI22_X1 U1240 ( .A1(n4550), .A2(n6373), .B1(n704), .B2(n269), .ZN(n3610) );
  OAI22_X1 U1241 ( .A1(n4518), .A2(n6374), .B1(n704), .B2(n271), .ZN(n3611) );
  OAI22_X1 U1242 ( .A1(n4486), .A2(n6377), .B1(n704), .B2(n273), .ZN(n3612) );
  OAI22_X1 U1243 ( .A1(n4454), .A2(n6378), .B1(n704), .B2(n275), .ZN(n3613) );
  OAI22_X1 U1244 ( .A1(n4422), .A2(n6381), .B1(n704), .B2(n277), .ZN(n3614) );
  OAI22_X1 U1245 ( .A1(n4390), .A2(n6384), .B1(n704), .B2(n279), .ZN(n3615) );
  OAI22_X1 U1246 ( .A1(n4358), .A2(n6383), .B1(n704), .B2(n281), .ZN(n3616) );
  OAI22_X1 U1247 ( .A1(n4326), .A2(n6391), .B1(n704), .B2(n283), .ZN(n3617) );
  OAI211_X1 U1249 ( .C1(n5623), .C2(n5345), .A(n716), .B(n717), .ZN(n713) );
  AOI222_X1 U1250 ( .A1(n718), .A2(n719), .B1(D_DATA_INBUS[22]), .B2(n720), 
        .C1(D_DATA_INBUS[6]), .C2(n721), .ZN(n717) );
  INV_X1 U1251 ( .A(n5677), .ZN(n719) );
  AOI22_X1 U1252 ( .A1(n722), .A2(n5678), .B1(n5675), .B2(n723), .ZN(n716) );
  OAI22_X1 U1253 ( .A1(n5345), .A2(\UUT/Mcontrol/N22 ), .B1(n703), .B2(n7394), 
        .ZN(n3618) );
  INV_X1 U1254 ( .A(n714), .ZN(n703) );
  OAI211_X1 U1255 ( .C1(n6102), .C2(n287), .A(n724), .B(n725), .ZN(n714) );
  AOI222_X1 U1256 ( .A1(\UUT/Mpath/the_mult/x_mult_out[6] ), .A2(n6357), .B1(
        n320), .B2(n726), .C1(n291), .C2(n727), .ZN(n725) );
  INV_X1 U1257 ( .A(n5594), .ZN(n727) );
  AOI22_X1 U1259 ( .A1(n6397), .A2(n728), .B1(n324), .B2(n6103), .ZN(n724) );
  INV_X1 U1260 ( .A(n5533), .ZN(n728) );
  OAI22_X1 U1261 ( .A1(n729), .A2(n556), .B1(n297), .B2(n2690), .ZN(n3619) );
  INV_X1 U1262 ( .A(\UUT/Mcontrol/Program_counter/N14 ), .ZN(n729) );
  OAI221_X1 U1263 ( .B1(n730), .B2(n80), .C1(n53), .C2(n81), .A(n731), .ZN(
        n3620) );
  NAND2_X1 U1264 ( .A1(n7080), .A2(n6340), .ZN(n731) );
  OAI222_X1 U1265 ( .A1(n53), .A2(n94), .B1(n730), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N74 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3621) );
  INV_X1 U1266 ( .A(\UUT/break_code[5] ), .ZN(n730) );
  INV_X1 U1267 ( .A(n732), .ZN(n53) );
  OAI222_X1 U1268 ( .A1(n733), .A2(n5332), .B1(n734), .B2(n101), .C1(n5347), 
        .C2(n102), .ZN(n732) );
  OAI221_X1 U1269 ( .B1(n103), .B2(n735), .C1(n5595), .C2(n105), .A(n736), 
        .ZN(n3622) );
  AOI22_X1 U1270 ( .A1(n107), .A2(n737), .B1(\UUT/Mpath/the_mult/Mad_out [37]), 
        .B2(n109), .ZN(n736) );
  OAI221_X1 U1271 ( .B1(n115), .B2(n738), .C1(n5535), .C2(n117), .A(n739), 
        .ZN(n3623) );
  AOI22_X1 U1272 ( .A1(n119), .A2(n737), .B1(\UUT/Mpath/the_mult/Mad_out [5]), 
        .B2(n121), .ZN(n739) );
  OAI22_X1 U1274 ( .A1(n7382), .A2(n740), .B1(n5536), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3624) );
  OAI221_X1 U1275 ( .B1(n741), .B2(n124), .C1(n125), .C2(n740), .A(n742), .ZN(
        n3625) );
  AOI22_X1 U1276 ( .A1(n127), .A2(n743), .B1(n129), .B2(n744), .ZN(n742) );
  INV_X1 U1277 ( .A(\UUT/Mpath/the_mult/x_operand1[5] ), .ZN(n740) );
  OAI221_X1 U1278 ( .B1(n741), .B2(n218), .C1(\UUT/Mpath/the_alu/N73 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n745), .ZN(n3626) );
  AOI22_X1 U1279 ( .A1(n220), .A2(n743), .B1(n221), .B2(n744), .ZN(n745) );
  OAI22_X1 U1280 ( .A1(n5287), .A2(n6393), .B1(n734), .B2(n223), .ZN(n3627) );
  OAI22_X1 U1281 ( .A1(n5255), .A2(n6396), .B1(n734), .B2(n225), .ZN(n3628) );
  OAI22_X1 U1282 ( .A1(n5223), .A2(n6387), .B1(n734), .B2(n227), .ZN(n3629) );
  OAI22_X1 U1283 ( .A1(n5191), .A2(n6395), .B1(n734), .B2(n229), .ZN(n3630) );
  OAI22_X1 U1284 ( .A1(n5159), .A2(n6390), .B1(n734), .B2(n231), .ZN(n3631) );
  OAI22_X1 U1285 ( .A1(n5127), .A2(n6385), .B1(n734), .B2(n233), .ZN(n3632) );
  OAI22_X1 U1286 ( .A1(n5095), .A2(n6389), .B1(n734), .B2(n235), .ZN(n3633) );
  OAI22_X1 U1287 ( .A1(n5063), .A2(n6382), .B1(n734), .B2(n237), .ZN(n3634) );
  OAI22_X1 U1288 ( .A1(n5031), .A2(n6380), .B1(n734), .B2(n239), .ZN(n3635) );
  OAI22_X1 U1289 ( .A1(n4999), .A2(n6379), .B1(n734), .B2(n241), .ZN(n3636) );
  OAI22_X1 U1290 ( .A1(n4967), .A2(n6376), .B1(n734), .B2(n243), .ZN(n3637) );
  OAI22_X1 U1291 ( .A1(n4935), .A2(n6375), .B1(n734), .B2(n245), .ZN(n3638) );
  OAI22_X1 U1292 ( .A1(n4903), .A2(n6372), .B1(n734), .B2(n247), .ZN(n3639) );
  OAI22_X1 U1293 ( .A1(n4871), .A2(n6371), .B1(n734), .B2(n249), .ZN(n3640) );
  OAI22_X1 U1294 ( .A1(n4839), .A2(n6368), .B1(n734), .B2(n251), .ZN(n3641) );
  OAI22_X1 U1295 ( .A1(n4807), .A2(n6367), .B1(n734), .B2(n253), .ZN(n3642) );
  OAI22_X1 U1296 ( .A1(n4775), .A2(n6364), .B1(n734), .B2(n255), .ZN(n3643) );
  OAI22_X1 U1297 ( .A1(n4743), .A2(n6362), .B1(n734), .B2(n257), .ZN(n3644) );
  OAI22_X1 U1298 ( .A1(n4711), .A2(n6361), .B1(n734), .B2(n259), .ZN(n3645) );
  OAI22_X1 U1299 ( .A1(n4679), .A2(n6365), .B1(n734), .B2(n261), .ZN(n3646) );
  OAI22_X1 U1300 ( .A1(n4647), .A2(n6366), .B1(n734), .B2(n263), .ZN(n3647) );
  OAI22_X1 U1301 ( .A1(n4615), .A2(n6369), .B1(n734), .B2(n265), .ZN(n3648) );
  OAI22_X1 U1302 ( .A1(n4583), .A2(n6370), .B1(n734), .B2(n267), .ZN(n3649) );
  OAI22_X1 U1303 ( .A1(n4551), .A2(n6373), .B1(n734), .B2(n269), .ZN(n3650) );
  OAI22_X1 U1304 ( .A1(n4519), .A2(n6374), .B1(n734), .B2(n271), .ZN(n3651) );
  OAI22_X1 U1305 ( .A1(n4487), .A2(n6377), .B1(n734), .B2(n273), .ZN(n3652) );
  OAI22_X1 U1306 ( .A1(n4455), .A2(n6378), .B1(n734), .B2(n275), .ZN(n3653) );
  OAI22_X1 U1307 ( .A1(n4423), .A2(n6381), .B1(n734), .B2(n277), .ZN(n3654) );
  OAI22_X1 U1308 ( .A1(n4391), .A2(n6384), .B1(n734), .B2(n279), .ZN(n3655) );
  OAI22_X1 U1309 ( .A1(n4359), .A2(n6383), .B1(n734), .B2(n281), .ZN(n3656) );
  OAI22_X1 U1310 ( .A1(n4327), .A2(n6391), .B1(n734), .B2(n283), .ZN(n3657) );
  OAI211_X1 U1312 ( .C1(n5623), .C2(n5348), .A(n746), .B(n747), .ZN(n743) );
  AOI222_X1 U1313 ( .A1(n718), .A2(n748), .B1(D_DATA_INBUS[21]), .B2(n720), 
        .C1(D_DATA_INBUS[5]), .C2(n721), .ZN(n747) );
  INV_X1 U1314 ( .A(n5687), .ZN(n748) );
  AOI22_X1 U1315 ( .A1(n722), .A2(n5688), .B1(n5685), .B2(n723), .ZN(n746) );
  OAI22_X1 U1316 ( .A1(n5348), .A2(\UUT/Mcontrol/N22 ), .B1(n733), .B2(n7394), 
        .ZN(n3658) );
  INV_X1 U1317 ( .A(n744), .ZN(n733) );
  OAI211_X1 U1318 ( .C1(n6104), .C2(n287), .A(n749), .B(n750), .ZN(n744) );
  AOI222_X1 U1319 ( .A1(\UUT/Mpath/the_mult/x_mult_out[5] ), .A2(n6357), .B1(
        n320), .B2(n751), .C1(n291), .C2(n752), .ZN(n750) );
  INV_X1 U1320 ( .A(n5595), .ZN(n752) );
  AOI22_X1 U1322 ( .A1(n6397), .A2(n753), .B1(n324), .B2(n6105), .ZN(n749) );
  INV_X1 U1323 ( .A(n5535), .ZN(n753) );
  OAI22_X1 U1324 ( .A1(n754), .A2(n556), .B1(n297), .B2(n2693), .ZN(n3659) );
  INV_X1 U1325 ( .A(\UUT/Mcontrol/Program_counter/N12 ), .ZN(n754) );
  OAI221_X1 U1326 ( .B1(n755), .B2(n80), .C1(n52), .C2(n81), .A(n756), .ZN(
        n3660) );
  NAND2_X1 U1327 ( .A1(\UUT/Mpath/the_mult/x_operand2 [4]), .A2(n6340), .ZN(
        n756) );
  OAI222_X1 U1328 ( .A1(n52), .A2(n94), .B1(n755), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N76 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3661) );
  INV_X1 U1329 ( .A(n757), .ZN(n52) );
  OAI222_X1 U1330 ( .A1(n758), .A2(n99), .B1(n759), .B2(n101), .C1(n5350), 
        .C2(n102), .ZN(n757) );
  OAI221_X1 U1331 ( .B1(n103), .B2(n760), .C1(n5596), .C2(n105), .A(n761), 
        .ZN(n3662) );
  AOI22_X1 U1332 ( .A1(n107), .A2(n762), .B1(\UUT/Mpath/the_mult/Mad_out [36]), 
        .B2(n109), .ZN(n761) );
  OAI221_X1 U1333 ( .B1(n115), .B2(n763), .C1(n5537), .C2(n117), .A(n764), 
        .ZN(n3663) );
  AOI22_X1 U1334 ( .A1(n119), .A2(n762), .B1(\UUT/Mpath/the_mult/Mad_out [4]), 
        .B2(n121), .ZN(n764) );
  OAI22_X1 U1336 ( .A1(n7383), .A2(n765), .B1(n5538), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3664) );
  OAI221_X1 U1337 ( .B1(n766), .B2(n124), .C1(n125), .C2(n765), .A(n767), .ZN(
        n3665) );
  AOI22_X1 U1338 ( .A1(n127), .A2(n768), .B1(n129), .B2(n769), .ZN(n767) );
  INV_X1 U1339 ( .A(\UUT/Mpath/the_mult/x_operand1[4] ), .ZN(n765) );
  OAI221_X1 U1340 ( .B1(n766), .B2(n218), .C1(\UUT/Mpath/the_alu/N75 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n770), .ZN(n3666) );
  AOI22_X1 U1341 ( .A1(n220), .A2(n768), .B1(n221), .B2(n769), .ZN(n770) );
  OAI22_X1 U1342 ( .A1(n5288), .A2(n6393), .B1(n759), .B2(n223), .ZN(n3667) );
  OAI22_X1 U1343 ( .A1(n5256), .A2(n6396), .B1(n759), .B2(n225), .ZN(n3668) );
  OAI22_X1 U1344 ( .A1(n5224), .A2(n6387), .B1(n759), .B2(n227), .ZN(n3669) );
  OAI22_X1 U1345 ( .A1(n5192), .A2(n6395), .B1(n759), .B2(n229), .ZN(n3670) );
  OAI22_X1 U1346 ( .A1(n5160), .A2(n6390), .B1(n759), .B2(n231), .ZN(n3671) );
  OAI22_X1 U1347 ( .A1(n5128), .A2(n6385), .B1(n759), .B2(n233), .ZN(n3672) );
  OAI22_X1 U1348 ( .A1(n5096), .A2(n6389), .B1(n759), .B2(n235), .ZN(n3673) );
  OAI22_X1 U1349 ( .A1(n5064), .A2(n6382), .B1(n759), .B2(n237), .ZN(n3674) );
  OAI22_X1 U1350 ( .A1(n5032), .A2(n6380), .B1(n759), .B2(n239), .ZN(n3675) );
  OAI22_X1 U1351 ( .A1(n5000), .A2(n6379), .B1(n759), .B2(n241), .ZN(n3676) );
  OAI22_X1 U1352 ( .A1(n4968), .A2(n6376), .B1(n759), .B2(n243), .ZN(n3677) );
  OAI22_X1 U1353 ( .A1(n4936), .A2(n6375), .B1(n759), .B2(n245), .ZN(n3678) );
  OAI22_X1 U1354 ( .A1(n4904), .A2(n6372), .B1(n759), .B2(n247), .ZN(n3679) );
  OAI22_X1 U1355 ( .A1(n4872), .A2(n6371), .B1(n759), .B2(n249), .ZN(n3680) );
  OAI22_X1 U1356 ( .A1(n4840), .A2(n6368), .B1(n759), .B2(n251), .ZN(n3681) );
  OAI22_X1 U1357 ( .A1(n4808), .A2(n6367), .B1(n759), .B2(n253), .ZN(n3682) );
  OAI22_X1 U1358 ( .A1(n4776), .A2(n6364), .B1(n759), .B2(n255), .ZN(n3683) );
  OAI22_X1 U1359 ( .A1(n4744), .A2(n6362), .B1(n759), .B2(n257), .ZN(n3684) );
  OAI22_X1 U1360 ( .A1(n4712), .A2(n6361), .B1(n759), .B2(n259), .ZN(n3685) );
  OAI22_X1 U1361 ( .A1(n4680), .A2(n6365), .B1(n759), .B2(n261), .ZN(n3686) );
  OAI22_X1 U1362 ( .A1(n4648), .A2(n6366), .B1(n759), .B2(n263), .ZN(n3687) );
  OAI22_X1 U1363 ( .A1(n4616), .A2(n6369), .B1(n759), .B2(n265), .ZN(n3688) );
  OAI22_X1 U1364 ( .A1(n4584), .A2(n6370), .B1(n759), .B2(n267), .ZN(n3689) );
  OAI22_X1 U1365 ( .A1(n4552), .A2(n6373), .B1(n759), .B2(n269), .ZN(n3690) );
  OAI22_X1 U1366 ( .A1(n4520), .A2(n6374), .B1(n759), .B2(n271), .ZN(n3691) );
  OAI22_X1 U1367 ( .A1(n4488), .A2(n6377), .B1(n759), .B2(n273), .ZN(n3692) );
  OAI22_X1 U1368 ( .A1(n4456), .A2(n6378), .B1(n759), .B2(n275), .ZN(n3693) );
  OAI22_X1 U1369 ( .A1(n4424), .A2(n6381), .B1(n759), .B2(n277), .ZN(n3694) );
  OAI22_X1 U1370 ( .A1(n4392), .A2(n6384), .B1(n759), .B2(n279), .ZN(n3695) );
  OAI22_X1 U1371 ( .A1(n4360), .A2(n6383), .B1(n759), .B2(n281), .ZN(n3696) );
  OAI22_X1 U1372 ( .A1(n4328), .A2(n6391), .B1(n759), .B2(n283), .ZN(n3697) );
  OAI211_X1 U1374 ( .C1(n5623), .C2(n5351), .A(n771), .B(n772), .ZN(n768) );
  AOI222_X1 U1375 ( .A1(n718), .A2(n773), .B1(D_DATA_INBUS[20]), .B2(n720), 
        .C1(D_DATA_INBUS[4]), .C2(n721), .ZN(n772) );
  INV_X1 U1376 ( .A(n5697), .ZN(n773) );
  AOI22_X1 U1377 ( .A1(n722), .A2(n5698), .B1(n5695), .B2(n723), .ZN(n771) );
  OAI22_X1 U1378 ( .A1(n5351), .A2(\UUT/Mcontrol/N22 ), .B1(n758), .B2(n7394), 
        .ZN(n3698) );
  INV_X1 U1379 ( .A(n769), .ZN(n758) );
  OAI211_X1 U1380 ( .C1(n6106), .C2(n287), .A(n774), .B(n775), .ZN(n769) );
  AOI222_X1 U1381 ( .A1(\UUT/Mpath/the_mult/x_mult_out[4] ), .A2(n6357), .B1(
        n320), .B2(n776), .C1(n291), .C2(n777), .ZN(n775) );
  INV_X1 U1382 ( .A(n5596), .ZN(n777) );
  AOI22_X1 U1384 ( .A1(n6397), .A2(n778), .B1(n324), .B2(n6107), .ZN(n774) );
  INV_X1 U1385 ( .A(n5537), .ZN(n778) );
  OAI22_X1 U1386 ( .A1(n779), .A2(n556), .B1(n297), .B2(n2696), .ZN(n3699) );
  INV_X1 U1387 ( .A(\UUT/Mcontrol/Program_counter/N10 ), .ZN(n779) );
  OAI221_X1 U1388 ( .B1(n7233), .B2(n80), .C1(n51), .C2(n81), .A(n781), .ZN(
        n3700) );
  NAND2_X1 U1389 ( .A1(n7066), .A2(n6340), .ZN(n781) );
  OAI222_X1 U1390 ( .A1(n51), .A2(n94), .B1(n7233), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N78 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3701) );
  INV_X1 U1391 ( .A(n782), .ZN(n51) );
  OAI222_X1 U1392 ( .A1(n783), .A2(n99), .B1(n784), .B2(n101), .C1(n5353), 
        .C2(n102), .ZN(n782) );
  OAI221_X1 U1393 ( .B1(n103), .B2(n785), .C1(n5597), .C2(n105), .A(n786), 
        .ZN(n3702) );
  AOI22_X1 U1394 ( .A1(n107), .A2(n787), .B1(\UUT/Mpath/the_mult/Mad_out [35]), 
        .B2(n109), .ZN(n786) );
  OAI221_X1 U1395 ( .B1(n115), .B2(n788), .C1(n5539), .C2(n117), .A(n789), 
        .ZN(n3703) );
  AOI22_X1 U1396 ( .A1(n119), .A2(n787), .B1(\UUT/Mpath/the_mult/Mad_out [3]), 
        .B2(n121), .ZN(n789) );
  OAI22_X1 U1398 ( .A1(n7382), .A2(n790), .B1(n5540), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3704) );
  OAI221_X1 U1399 ( .B1(n791), .B2(n124), .C1(n125), .C2(n790), .A(n792), .ZN(
        n3705) );
  AOI22_X1 U1400 ( .A1(n127), .A2(n793), .B1(n129), .B2(n794), .ZN(n792) );
  INV_X1 U1401 ( .A(\UUT/Mpath/the_mult/x_operand1[3] ), .ZN(n790) );
  OAI221_X1 U1402 ( .B1(n791), .B2(n218), .C1(\UUT/Mpath/the_alu/N77 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n795), .ZN(n3706) );
  AOI22_X1 U1403 ( .A1(n220), .A2(n793), .B1(n221), .B2(n794), .ZN(n795) );
  OAI22_X1 U1404 ( .A1(n5289), .A2(n6393), .B1(n784), .B2(n223), .ZN(n3707) );
  OAI22_X1 U1405 ( .A1(n5257), .A2(n6396), .B1(n784), .B2(n225), .ZN(n3708) );
  OAI22_X1 U1406 ( .A1(n5225), .A2(n6387), .B1(n784), .B2(n227), .ZN(n3709) );
  OAI22_X1 U1407 ( .A1(n5193), .A2(n6395), .B1(n784), .B2(n229), .ZN(n3710) );
  OAI22_X1 U1408 ( .A1(n5161), .A2(n6390), .B1(n784), .B2(n231), .ZN(n3711) );
  OAI22_X1 U1409 ( .A1(n5129), .A2(n6385), .B1(n784), .B2(n233), .ZN(n3712) );
  OAI22_X1 U1410 ( .A1(n5097), .A2(n6389), .B1(n784), .B2(n235), .ZN(n3713) );
  OAI22_X1 U1411 ( .A1(n5065), .A2(n6382), .B1(n784), .B2(n237), .ZN(n3714) );
  OAI22_X1 U1412 ( .A1(n5033), .A2(n6380), .B1(n784), .B2(n239), .ZN(n3715) );
  OAI22_X1 U1413 ( .A1(n5001), .A2(n6379), .B1(n784), .B2(n241), .ZN(n3716) );
  OAI22_X1 U1414 ( .A1(n4969), .A2(n6376), .B1(n784), .B2(n243), .ZN(n3717) );
  OAI22_X1 U1415 ( .A1(n4937), .A2(n6375), .B1(n784), .B2(n245), .ZN(n3718) );
  OAI22_X1 U1416 ( .A1(n4905), .A2(n6372), .B1(n784), .B2(n247), .ZN(n3719) );
  OAI22_X1 U1417 ( .A1(n4873), .A2(n6371), .B1(n784), .B2(n249), .ZN(n3720) );
  OAI22_X1 U1418 ( .A1(n4841), .A2(n6368), .B1(n784), .B2(n251), .ZN(n3721) );
  OAI22_X1 U1419 ( .A1(n4809), .A2(n6367), .B1(n784), .B2(n253), .ZN(n3722) );
  OAI22_X1 U1420 ( .A1(n4777), .A2(n6364), .B1(n784), .B2(n255), .ZN(n3723) );
  OAI22_X1 U1421 ( .A1(n4745), .A2(n6362), .B1(n784), .B2(n257), .ZN(n3724) );
  OAI22_X1 U1422 ( .A1(n4713), .A2(n6361), .B1(n784), .B2(n259), .ZN(n3725) );
  OAI22_X1 U1423 ( .A1(n4681), .A2(n6365), .B1(n784), .B2(n261), .ZN(n3726) );
  OAI22_X1 U1424 ( .A1(n4649), .A2(n6366), .B1(n784), .B2(n263), .ZN(n3727) );
  OAI22_X1 U1425 ( .A1(n4617), .A2(n6369), .B1(n784), .B2(n265), .ZN(n3728) );
  OAI22_X1 U1426 ( .A1(n4585), .A2(n6370), .B1(n784), .B2(n267), .ZN(n3729) );
  OAI22_X1 U1427 ( .A1(n4553), .A2(n6373), .B1(n784), .B2(n269), .ZN(n3730) );
  OAI22_X1 U1428 ( .A1(n4521), .A2(n6374), .B1(n784), .B2(n271), .ZN(n3731) );
  OAI22_X1 U1429 ( .A1(n4489), .A2(n6377), .B1(n784), .B2(n273), .ZN(n3732) );
  OAI22_X1 U1430 ( .A1(n4457), .A2(n6378), .B1(n784), .B2(n275), .ZN(n3733) );
  OAI22_X1 U1431 ( .A1(n4425), .A2(n6381), .B1(n784), .B2(n277), .ZN(n3734) );
  OAI22_X1 U1432 ( .A1(n4393), .A2(n6384), .B1(n784), .B2(n279), .ZN(n3735) );
  OAI22_X1 U1433 ( .A1(n4361), .A2(n6383), .B1(n784), .B2(n281), .ZN(n3736) );
  OAI22_X1 U1434 ( .A1(n4329), .A2(n6391), .B1(n784), .B2(n283), .ZN(n3737) );
  OAI211_X1 U1436 ( .C1(n5623), .C2(n5354), .A(n796), .B(n797), .ZN(n793) );
  AOI222_X1 U1437 ( .A1(n718), .A2(n798), .B1(D_DATA_INBUS[19]), .B2(n720), 
        .C1(D_DATA_INBUS[3]), .C2(n721), .ZN(n797) );
  INV_X1 U1438 ( .A(n5707), .ZN(n798) );
  AOI22_X1 U1439 ( .A1(n722), .A2(n5708), .B1(n5705), .B2(n723), .ZN(n796) );
  OAI22_X1 U1440 ( .A1(n5354), .A2(\UUT/Mcontrol/N22 ), .B1(n783), .B2(n7394), 
        .ZN(n3738) );
  INV_X1 U1441 ( .A(n794), .ZN(n783) );
  OAI211_X1 U1442 ( .C1(n6108), .C2(n287), .A(n799), .B(n800), .ZN(n794) );
  AOI222_X1 U1443 ( .A1(\UUT/Mpath/the_mult/x_mult_out[3] ), .A2(n6357), .B1(
        n320), .B2(n801), .C1(n291), .C2(n802), .ZN(n800) );
  INV_X1 U1444 ( .A(n5597), .ZN(n802) );
  AOI22_X1 U1446 ( .A1(n6397), .A2(n803), .B1(n324), .B2(n6109), .ZN(n799) );
  INV_X1 U1447 ( .A(n5539), .ZN(n803) );
  OAI22_X1 U1448 ( .A1(n804), .A2(n556), .B1(n297), .B2(n2699), .ZN(n3739) );
  INV_X1 U1449 ( .A(\UUT/Mcontrol/Program_counter/N8 ), .ZN(n804) );
  OAI221_X1 U1450 ( .B1(n805), .B2(n80), .C1(n50), .C2(n81), .A(n806), .ZN(
        n3740) );
  NAND2_X1 U1451 ( .A1(\UUT/Mpath/the_mult/x_operand2 [2]), .A2(n6340), .ZN(
        n806) );
  INV_X1 U1453 ( .A(n807), .ZN(n50) );
  OAI222_X1 U1454 ( .A1(n808), .A2(n99), .B1(n809), .B2(n101), .C1(n5362), 
        .C2(n102), .ZN(n807) );
  OAI221_X1 U1455 ( .B1(n103), .B2(n810), .C1(n5600), .C2(n105), .A(n811), 
        .ZN(n3742) );
  AOI22_X1 U1456 ( .A1(n107), .A2(n812), .B1(\UUT/Mpath/the_mult/Mad_out [34]), 
        .B2(n109), .ZN(n811) );
  OAI221_X1 U1457 ( .B1(n115), .B2(n813), .C1(n5545), .C2(n117), .A(n814), 
        .ZN(n3743) );
  AOI22_X1 U1458 ( .A1(n119), .A2(n812), .B1(\UUT/Mpath/the_mult/Mad_out [2]), 
        .B2(n121), .ZN(n814) );
  OAI22_X1 U1460 ( .A1(n7384), .A2(n815), .B1(n5546), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3744) );
  OAI221_X1 U1461 ( .B1(n816), .B2(n124), .C1(n125), .C2(n815), .A(n817), .ZN(
        n3745) );
  AOI22_X1 U1462 ( .A1(n127), .A2(n818), .B1(n129), .B2(n819), .ZN(n817) );
  INV_X1 U1463 ( .A(\UUT/Mpath/the_mult/x_operand1[2] ), .ZN(n815) );
  OAI221_X1 U1464 ( .B1(n816), .B2(n218), .C1(\UUT/Mpath/the_alu/N79 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n820), .ZN(n3746) );
  AOI22_X1 U1465 ( .A1(n220), .A2(n818), .B1(n221), .B2(n819), .ZN(n820) );
  OAI22_X1 U1466 ( .A1(n5292), .A2(n6393), .B1(n809), .B2(n223), .ZN(n3747) );
  OAI22_X1 U1467 ( .A1(n5260), .A2(n6396), .B1(n809), .B2(n225), .ZN(n3748) );
  OAI22_X1 U1468 ( .A1(n5228), .A2(n6387), .B1(n809), .B2(n227), .ZN(n3749) );
  OAI22_X1 U1469 ( .A1(n5196), .A2(n6395), .B1(n809), .B2(n229), .ZN(n3750) );
  OAI22_X1 U1470 ( .A1(n5164), .A2(n6390), .B1(n809), .B2(n231), .ZN(n3751) );
  OAI22_X1 U1471 ( .A1(n5132), .A2(n6385), .B1(n809), .B2(n233), .ZN(n3752) );
  OAI22_X1 U1472 ( .A1(n5100), .A2(n6389), .B1(n809), .B2(n235), .ZN(n3753) );
  OAI22_X1 U1473 ( .A1(n5068), .A2(n6382), .B1(n809), .B2(n237), .ZN(n3754) );
  OAI22_X1 U1474 ( .A1(n5036), .A2(n6380), .B1(n809), .B2(n239), .ZN(n3755) );
  OAI22_X1 U1475 ( .A1(n5004), .A2(n6379), .B1(n809), .B2(n241), .ZN(n3756) );
  OAI22_X1 U1476 ( .A1(n4972), .A2(n6376), .B1(n809), .B2(n243), .ZN(n3757) );
  OAI22_X1 U1477 ( .A1(n4940), .A2(n6375), .B1(n809), .B2(n245), .ZN(n3758) );
  OAI22_X1 U1478 ( .A1(n4908), .A2(n6372), .B1(n809), .B2(n247), .ZN(n3759) );
  OAI22_X1 U1479 ( .A1(n4876), .A2(n6371), .B1(n809), .B2(n249), .ZN(n3760) );
  OAI22_X1 U1480 ( .A1(n4844), .A2(n6368), .B1(n809), .B2(n251), .ZN(n3761) );
  OAI22_X1 U1481 ( .A1(n4812), .A2(n6367), .B1(n809), .B2(n253), .ZN(n3762) );
  OAI22_X1 U1482 ( .A1(n4780), .A2(n6364), .B1(n809), .B2(n255), .ZN(n3763) );
  OAI22_X1 U1483 ( .A1(n4748), .A2(n6362), .B1(n809), .B2(n257), .ZN(n3764) );
  OAI22_X1 U1484 ( .A1(n4716), .A2(n6361), .B1(n809), .B2(n259), .ZN(n3765) );
  OAI22_X1 U1485 ( .A1(n4684), .A2(n6365), .B1(n809), .B2(n261), .ZN(n3766) );
  OAI22_X1 U1486 ( .A1(n4652), .A2(n6366), .B1(n809), .B2(n263), .ZN(n3767) );
  OAI22_X1 U1487 ( .A1(n4620), .A2(n6369), .B1(n809), .B2(n265), .ZN(n3768) );
  OAI22_X1 U1488 ( .A1(n4588), .A2(n6370), .B1(n809), .B2(n267), .ZN(n3769) );
  OAI22_X1 U1489 ( .A1(n4556), .A2(n6373), .B1(n809), .B2(n269), .ZN(n3770) );
  OAI22_X1 U1490 ( .A1(n4524), .A2(n6374), .B1(n809), .B2(n271), .ZN(n3771) );
  OAI22_X1 U1491 ( .A1(n4492), .A2(n6377), .B1(n809), .B2(n273), .ZN(n3772) );
  OAI22_X1 U1492 ( .A1(n4460), .A2(n6378), .B1(n809), .B2(n275), .ZN(n3773) );
  OAI22_X1 U1493 ( .A1(n4428), .A2(n6381), .B1(n809), .B2(n277), .ZN(n3774) );
  OAI22_X1 U1494 ( .A1(n4396), .A2(n6384), .B1(n809), .B2(n279), .ZN(n3775) );
  OAI22_X1 U1495 ( .A1(n4364), .A2(n6383), .B1(n809), .B2(n281), .ZN(n3776) );
  OAI22_X1 U1496 ( .A1(n4332), .A2(n6391), .B1(n809), .B2(n283), .ZN(n3777) );
  OAI211_X1 U1498 ( .C1(n5623), .C2(n5363), .A(n821), .B(n822), .ZN(n818) );
  AOI222_X1 U1499 ( .A1(n718), .A2(n823), .B1(D_DATA_INBUS[18]), .B2(n720), 
        .C1(D_DATA_INBUS[2]), .C2(n721), .ZN(n822) );
  NOR2_X1 U1500 ( .A1(n824), .A2(n825), .ZN(n721) );
  AOI22_X1 U1501 ( .A1(\UUT/Mpath/the_memhandle/N39 ), .A2(n826), .B1(n5663), 
        .B2(n5856), .ZN(n824) );
  AND2_X1 U1502 ( .A1(n723), .A2(n5664), .ZN(n720) );
  INV_X1 U1503 ( .A(n5728), .ZN(n823) );
  AND2_X1 U1504 ( .A1(n722), .A2(\UUT/Mpath/the_memhandle/N36 ), .ZN(n718) );
  AOI22_X1 U1505 ( .A1(n722), .A2(n5729), .B1(n5726), .B2(n723), .ZN(n821) );
  INV_X1 U1506 ( .A(n692), .ZN(n723) );
  INV_X1 U1507 ( .A(n827), .ZN(n722) );
  OAI22_X1 U1508 ( .A1(n5363), .A2(\UUT/Mcontrol/N22 ), .B1(n808), .B2(n7394), 
        .ZN(n3778) );
  INV_X1 U1509 ( .A(n819), .ZN(n808) );
  OAI211_X1 U1510 ( .C1(n6112), .C2(n287), .A(n828), .B(n829), .ZN(n819) );
  AOI222_X1 U1511 ( .A1(\UUT/Mpath/the_mult/x_mult_out[2] ), .A2(n6357), .B1(
        n320), .B2(n830), .C1(n291), .C2(n831), .ZN(n829) );
  INV_X1 U1512 ( .A(n5600), .ZN(n831) );
  AOI22_X1 U1514 ( .A1(n6397), .A2(n832), .B1(n324), .B2(n6113), .ZN(n828) );
  INV_X1 U1515 ( .A(n5545), .ZN(n832) );
  OAI221_X1 U1516 ( .B1(n833), .B2(n80), .C1(n49), .C2(n81), .A(n834), .ZN(
        n3779) );
  NAND2_X1 U1517 ( .A1(\UUT/Mpath/the_mult/x_operand2 [1]), .A2(n6340), .ZN(
        n834) );
  NAND2_X1 U1518 ( .A1(n125), .A2(n835), .ZN(n81) );
  OR2_X1 U1519 ( .A1(n6340), .A2(n835), .ZN(n80) );
  AOI222_X1 U1521 ( .A1(n6867), .A2(\UUT/jar_in [1]), .B1(n300), .B2(
        \UUT/branch_rega [1]), .C1(\UUT/Mcontrol/Nextpc_decoding/Bta [1]), 
        .C2(n301), .ZN(n836) );
  OAI221_X1 U1522 ( .B1(n103), .B2(n837), .C1(n5622), .C2(n105), .A(n838), 
        .ZN(n3781) );
  AOI22_X1 U1523 ( .A1(n107), .A2(n839), .B1(\UUT/Mpath/the_mult/Mad_out [32]), 
        .B2(n109), .ZN(n838) );
  OAI221_X1 U1524 ( .B1(n115), .B2(n840), .C1(n5589), .C2(n117), .A(n841), 
        .ZN(n3782) );
  AOI22_X1 U1525 ( .A1(n119), .A2(n839), .B1(\UUT/Mpath/the_mult/Mad_out [0]), 
        .B2(n121), .ZN(n841) );
  OAI22_X1 U1527 ( .A1(n7382), .A2(n842), .B1(n5590), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3783) );
  OAI221_X1 U1528 ( .B1(n5324), .B2(n124), .C1(n125), .C2(n842), .A(n843), 
        .ZN(n3784) );
  AOI22_X1 U1529 ( .A1(n127), .A2(n844), .B1(n129), .B2(n845), .ZN(n843) );
  INV_X1 U1530 ( .A(\UUT/Mpath/the_mult/x_operand1[0] ), .ZN(n842) );
  OAI221_X1 U1531 ( .B1(n5324), .B2(n218), .C1(\UUT/Mpath/the_alu/N83 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n846), .ZN(n3785) );
  AOI22_X1 U1532 ( .A1(n220), .A2(n844), .B1(n221), .B2(n845), .ZN(n846) );
  OAI22_X1 U1533 ( .A1(n5314), .A2(n6393), .B1(n847), .B2(n223), .ZN(n3786) );
  OAI22_X1 U1534 ( .A1(n5282), .A2(n6396), .B1(n847), .B2(n225), .ZN(n3787) );
  OAI22_X1 U1535 ( .A1(n5250), .A2(n6387), .B1(n847), .B2(n227), .ZN(n3788) );
  OAI22_X1 U1536 ( .A1(n5218), .A2(n6395), .B1(n847), .B2(n229), .ZN(n3789) );
  OAI22_X1 U1537 ( .A1(n5186), .A2(n6390), .B1(n847), .B2(n231), .ZN(n3790) );
  OAI22_X1 U1538 ( .A1(n5154), .A2(n6385), .B1(n847), .B2(n233), .ZN(n3791) );
  OAI22_X1 U1539 ( .A1(n5122), .A2(n6389), .B1(n847), .B2(n235), .ZN(n3792) );
  OAI22_X1 U1540 ( .A1(n5090), .A2(n6382), .B1(n847), .B2(n237), .ZN(n3793) );
  OAI22_X1 U1541 ( .A1(n5058), .A2(n6380), .B1(n847), .B2(n239), .ZN(n3794) );
  OAI22_X1 U1542 ( .A1(n5026), .A2(n6379), .B1(n847), .B2(n241), .ZN(n3795) );
  OAI22_X1 U1543 ( .A1(n4994), .A2(n6376), .B1(n847), .B2(n243), .ZN(n3796) );
  OAI22_X1 U1544 ( .A1(n4962), .A2(n6375), .B1(n847), .B2(n245), .ZN(n3797) );
  OAI22_X1 U1545 ( .A1(n4930), .A2(n6372), .B1(n847), .B2(n247), .ZN(n3798) );
  OAI22_X1 U1546 ( .A1(n4898), .A2(n6371), .B1(n847), .B2(n249), .ZN(n3799) );
  OAI22_X1 U1547 ( .A1(n4866), .A2(n6368), .B1(n847), .B2(n251), .ZN(n3800) );
  OAI22_X1 U1548 ( .A1(n4834), .A2(n6367), .B1(n847), .B2(n253), .ZN(n3801) );
  OAI22_X1 U1549 ( .A1(n4802), .A2(n6364), .B1(n847), .B2(n255), .ZN(n3802) );
  OAI22_X1 U1550 ( .A1(n4770), .A2(n6362), .B1(n847), .B2(n257), .ZN(n3803) );
  OAI22_X1 U1551 ( .A1(n4738), .A2(n6361), .B1(n847), .B2(n259), .ZN(n3804) );
  OAI22_X1 U1552 ( .A1(n4706), .A2(n6365), .B1(n847), .B2(n261), .ZN(n3805) );
  OAI22_X1 U1553 ( .A1(n4674), .A2(n6366), .B1(n847), .B2(n263), .ZN(n3806) );
  OAI22_X1 U1554 ( .A1(n4642), .A2(n6369), .B1(n847), .B2(n265), .ZN(n3807) );
  OAI22_X1 U1555 ( .A1(n4610), .A2(n6370), .B1(n847), .B2(n267), .ZN(n3808) );
  OAI22_X1 U1556 ( .A1(n4578), .A2(n6373), .B1(n847), .B2(n269), .ZN(n3809) );
  OAI22_X1 U1557 ( .A1(n4546), .A2(n6374), .B1(n847), .B2(n271), .ZN(n3810) );
  OAI22_X1 U1558 ( .A1(n4514), .A2(n6377), .B1(n847), .B2(n273), .ZN(n3811) );
  OAI22_X1 U1559 ( .A1(n4482), .A2(n6378), .B1(n847), .B2(n275), .ZN(n3812) );
  OAI22_X1 U1560 ( .A1(n4450), .A2(n6381), .B1(n847), .B2(n277), .ZN(n3813) );
  OAI22_X1 U1561 ( .A1(n4418), .A2(n6384), .B1(n847), .B2(n279), .ZN(n3814) );
  OAI22_X1 U1562 ( .A1(n4386), .A2(n6383), .B1(n847), .B2(n281), .ZN(n3815) );
  OAI22_X1 U1563 ( .A1(n4354), .A2(n6391), .B1(n847), .B2(n283), .ZN(n3816) );
  OAI221_X1 U1564 ( .B1(n103), .B2(n848), .C1(n5611), .C2(n105), .A(n849), 
        .ZN(n3817) );
  AOI22_X1 U1565 ( .A1(n107), .A2(n850), .B1(\UUT/Mpath/the_mult/Mad_out [33]), 
        .B2(n109), .ZN(n849) );
  OAI221_X1 U1566 ( .B1(n115), .B2(n851), .C1(n5567), .C2(n117), .A(n852), 
        .ZN(n3818) );
  AOI22_X1 U1567 ( .A1(n119), .A2(n850), .B1(\UUT/Mpath/the_mult/Mad_out [1]), 
        .B2(n121), .ZN(n852) );
  OAI22_X1 U1569 ( .A1(n7383), .A2(n853), .B1(n5568), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3819) );
  OAI221_X1 U1570 ( .B1(n854), .B2(n124), .C1(n125), .C2(n853), .A(n855), .ZN(
        n3820) );
  AOI22_X1 U1571 ( .A1(n127), .A2(n856), .B1(n129), .B2(n857), .ZN(n855) );
  INV_X1 U1572 ( .A(\UUT/Mpath/the_mult/x_operand1[1] ), .ZN(n853) );
  OAI221_X1 U1573 ( .B1(n854), .B2(n218), .C1(\UUT/Mpath/the_alu/N81 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n858), .ZN(n3821) );
  AOI22_X1 U1574 ( .A1(n220), .A2(n856), .B1(n221), .B2(n857), .ZN(n858) );
  OAI22_X1 U1575 ( .A1(n5303), .A2(n6393), .B1(n859), .B2(n223), .ZN(n3822) );
  OAI22_X1 U1576 ( .A1(n5271), .A2(n6396), .B1(n859), .B2(n225), .ZN(n3823) );
  OAI22_X1 U1577 ( .A1(n5239), .A2(n6387), .B1(n859), .B2(n227), .ZN(n3824) );
  OAI22_X1 U1578 ( .A1(n5207), .A2(n6395), .B1(n859), .B2(n229), .ZN(n3825) );
  OAI22_X1 U1579 ( .A1(n5175), .A2(n6390), .B1(n859), .B2(n231), .ZN(n3826) );
  OAI22_X1 U1580 ( .A1(n5143), .A2(n6385), .B1(n859), .B2(n233), .ZN(n3827) );
  OAI22_X1 U1581 ( .A1(n5111), .A2(n6389), .B1(n859), .B2(n235), .ZN(n3828) );
  OAI22_X1 U1582 ( .A1(n5079), .A2(n6382), .B1(n859), .B2(n237), .ZN(n3829) );
  OAI22_X1 U1583 ( .A1(n5047), .A2(n6380), .B1(n859), .B2(n239), .ZN(n3830) );
  OAI22_X1 U1584 ( .A1(n5015), .A2(n6379), .B1(n859), .B2(n241), .ZN(n3831) );
  OAI22_X1 U1585 ( .A1(n4983), .A2(n6376), .B1(n859), .B2(n243), .ZN(n3832) );
  OAI22_X1 U1586 ( .A1(n4951), .A2(n6375), .B1(n859), .B2(n245), .ZN(n3833) );
  OAI22_X1 U1587 ( .A1(n4919), .A2(n6372), .B1(n859), .B2(n247), .ZN(n3834) );
  OAI22_X1 U1588 ( .A1(n4887), .A2(n6371), .B1(n859), .B2(n249), .ZN(n3835) );
  OAI22_X1 U1589 ( .A1(n4855), .A2(n6368), .B1(n859), .B2(n251), .ZN(n3836) );
  OAI22_X1 U1590 ( .A1(n4823), .A2(n6367), .B1(n859), .B2(n253), .ZN(n3837) );
  OAI22_X1 U1591 ( .A1(n4791), .A2(n6364), .B1(n859), .B2(n255), .ZN(n3838) );
  OAI22_X1 U1592 ( .A1(n4759), .A2(n6362), .B1(n859), .B2(n257), .ZN(n3839) );
  OAI22_X1 U1593 ( .A1(n4727), .A2(n6361), .B1(n859), .B2(n259), .ZN(n3840) );
  OAI22_X1 U1594 ( .A1(n4695), .A2(n6365), .B1(n859), .B2(n261), .ZN(n3841) );
  OAI22_X1 U1595 ( .A1(n4663), .A2(n6366), .B1(n859), .B2(n263), .ZN(n3842) );
  OAI22_X1 U1596 ( .A1(n4631), .A2(n6369), .B1(n859), .B2(n265), .ZN(n3843) );
  OAI22_X1 U1597 ( .A1(n4599), .A2(n6370), .B1(n859), .B2(n267), .ZN(n3844) );
  OAI22_X1 U1598 ( .A1(n4567), .A2(n6373), .B1(n859), .B2(n269), .ZN(n3845) );
  OAI22_X1 U1599 ( .A1(n4535), .A2(n6374), .B1(n859), .B2(n271), .ZN(n3846) );
  OAI22_X1 U1600 ( .A1(n4503), .A2(n6377), .B1(n859), .B2(n273), .ZN(n3847) );
  OAI22_X1 U1601 ( .A1(n4471), .A2(n6378), .B1(n859), .B2(n275), .ZN(n3848) );
  OAI22_X1 U1602 ( .A1(n4439), .A2(n6381), .B1(n859), .B2(n277), .ZN(n3849) );
  OAI22_X1 U1603 ( .A1(n4407), .A2(n6384), .B1(n859), .B2(n279), .ZN(n3850) );
  OAI22_X1 U1604 ( .A1(n4375), .A2(n6383), .B1(n859), .B2(n281), .ZN(n3851) );
  OAI22_X1 U1605 ( .A1(n4343), .A2(n6391), .B1(n859), .B2(n283), .ZN(n3852) );
  OAI221_X1 U1606 ( .B1(n103), .B2(n860), .C1(n5607), .C2(n105), .A(n861), 
        .ZN(n3853) );
  AOI22_X1 U1607 ( .A1(n107), .A2(n862), .B1(\UUT/Mpath/the_mult/Mad_out [55]), 
        .B2(n109), .ZN(n861) );
  OAI221_X1 U1608 ( .B1(n115), .B2(n863), .C1(n5559), .C2(n117), .A(n864), 
        .ZN(n3854) );
  AOI22_X1 U1609 ( .A1(n119), .A2(n862), .B1(\UUT/Mpath/the_mult/Mad_out [23]), 
        .B2(n121), .ZN(n864) );
  OAI22_X1 U1611 ( .A1(n7382), .A2(n865), .B1(n5560), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n3855) );
  OAI221_X1 U1612 ( .B1(n866), .B2(n124), .C1(n125), .C2(n865), .A(n867), .ZN(
        n3856) );
  AOI22_X1 U1613 ( .A1(n127), .A2(n868), .B1(n129), .B2(n869), .ZN(n867) );
  INV_X1 U1614 ( .A(\UUT/Mpath/the_mult/x_operand1[23] ), .ZN(n865) );
  OAI221_X1 U1615 ( .B1(n866), .B2(n218), .C1(\UUT/Mpath/the_alu/N37 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n870), .ZN(n3857) );
  AOI22_X1 U1616 ( .A1(n220), .A2(n868), .B1(n221), .B2(n869), .ZN(n870) );
  OAI22_X1 U1617 ( .A1(n5299), .A2(n6393), .B1(n871), .B2(n223), .ZN(n3858) );
  OAI22_X1 U1618 ( .A1(n5267), .A2(n6396), .B1(n871), .B2(n225), .ZN(n3859) );
  OAI22_X1 U1619 ( .A1(n5235), .A2(n6387), .B1(n871), .B2(n227), .ZN(n3860) );
  OAI22_X1 U1620 ( .A1(n5203), .A2(n6395), .B1(n871), .B2(n229), .ZN(n3861) );
  OAI22_X1 U1621 ( .A1(n5171), .A2(n6390), .B1(n871), .B2(n231), .ZN(n3862) );
  OAI22_X1 U1622 ( .A1(n5139), .A2(n6385), .B1(n871), .B2(n233), .ZN(n3863) );
  OAI22_X1 U1623 ( .A1(n5107), .A2(n6389), .B1(n871), .B2(n235), .ZN(n3864) );
  OAI22_X1 U1624 ( .A1(n5075), .A2(n6382), .B1(n871), .B2(n237), .ZN(n3865) );
  OAI22_X1 U1625 ( .A1(n5043), .A2(n6380), .B1(n871), .B2(n239), .ZN(n3866) );
  OAI22_X1 U1626 ( .A1(n5011), .A2(n6379), .B1(n871), .B2(n241), .ZN(n3867) );
  OAI22_X1 U1627 ( .A1(n4979), .A2(n6376), .B1(n871), .B2(n243), .ZN(n3868) );
  OAI22_X1 U1628 ( .A1(n4947), .A2(n6375), .B1(n871), .B2(n245), .ZN(n3869) );
  OAI22_X1 U1629 ( .A1(n4915), .A2(n6372), .B1(n871), .B2(n247), .ZN(n3870) );
  OAI22_X1 U1630 ( .A1(n4883), .A2(n6371), .B1(n871), .B2(n249), .ZN(n3871) );
  OAI22_X1 U1631 ( .A1(n4851), .A2(n6368), .B1(n871), .B2(n251), .ZN(n3872) );
  OAI22_X1 U1632 ( .A1(n4819), .A2(n6367), .B1(n871), .B2(n253), .ZN(n3873) );
  OAI22_X1 U1633 ( .A1(n4787), .A2(n6364), .B1(n871), .B2(n255), .ZN(n3874) );
  OAI22_X1 U1634 ( .A1(n4755), .A2(n6362), .B1(n871), .B2(n257), .ZN(n3875) );
  OAI22_X1 U1635 ( .A1(n4723), .A2(n6361), .B1(n871), .B2(n259), .ZN(n3876) );
  OAI22_X1 U1636 ( .A1(n4691), .A2(n6365), .B1(n871), .B2(n261), .ZN(n3877) );
  OAI22_X1 U1637 ( .A1(n4659), .A2(n6366), .B1(n871), .B2(n263), .ZN(n3878) );
  OAI22_X1 U1638 ( .A1(n4627), .A2(n6369), .B1(n871), .B2(n265), .ZN(n3879) );
  OAI22_X1 U1639 ( .A1(n4595), .A2(n6370), .B1(n871), .B2(n267), .ZN(n3880) );
  OAI22_X1 U1640 ( .A1(n4563), .A2(n6373), .B1(n871), .B2(n269), .ZN(n3881) );
  OAI22_X1 U1641 ( .A1(n4531), .A2(n6374), .B1(n871), .B2(n271), .ZN(n3882) );
  OAI22_X1 U1642 ( .A1(n4499), .A2(n6377), .B1(n871), .B2(n273), .ZN(n3883) );
  OAI22_X1 U1643 ( .A1(n4467), .A2(n6378), .B1(n871), .B2(n275), .ZN(n3884) );
  OAI22_X1 U1644 ( .A1(n4435), .A2(n6381), .B1(n871), .B2(n277), .ZN(n3885) );
  OAI22_X1 U1645 ( .A1(n4403), .A2(n6384), .B1(n871), .B2(n279), .ZN(n3886) );
  OAI22_X1 U1646 ( .A1(n4371), .A2(n6383), .B1(n871), .B2(n281), .ZN(n3887) );
  OAI22_X1 U1647 ( .A1(n4339), .A2(n6391), .B1(n871), .B2(n283), .ZN(n3888) );
  OAI22_X1 U1648 ( .A1(n5297), .A2(n6393), .B1(n185), .B2(n223), .ZN(n3889) );
  OAI22_X1 U1649 ( .A1(n5265), .A2(n6396), .B1(n185), .B2(n225), .ZN(n3890) );
  OAI22_X1 U1650 ( .A1(n5233), .A2(n6387), .B1(n185), .B2(n227), .ZN(n3891) );
  OAI22_X1 U1651 ( .A1(n5201), .A2(n6395), .B1(n185), .B2(n229), .ZN(n3892) );
  OAI22_X1 U1652 ( .A1(n5169), .A2(n6390), .B1(n185), .B2(n231), .ZN(n3893) );
  OAI22_X1 U1653 ( .A1(n5137), .A2(n6385), .B1(n185), .B2(n233), .ZN(n3894) );
  OAI22_X1 U1654 ( .A1(n5105), .A2(n6389), .B1(n185), .B2(n235), .ZN(n3895) );
  OAI22_X1 U1655 ( .A1(n5073), .A2(n6382), .B1(n185), .B2(n237), .ZN(n3896) );
  OAI22_X1 U1656 ( .A1(n5041), .A2(n6380), .B1(n185), .B2(n239), .ZN(n3897) );
  OAI22_X1 U1657 ( .A1(n5009), .A2(n6379), .B1(n185), .B2(n241), .ZN(n3898) );
  OAI22_X1 U1658 ( .A1(n4977), .A2(n6376), .B1(n185), .B2(n243), .ZN(n3899) );
  OAI22_X1 U1659 ( .A1(n4945), .A2(n6375), .B1(n185), .B2(n245), .ZN(n3900) );
  OAI22_X1 U1660 ( .A1(n4913), .A2(n6372), .B1(n185), .B2(n247), .ZN(n3901) );
  OAI22_X1 U1661 ( .A1(n4881), .A2(n6371), .B1(n185), .B2(n249), .ZN(n3902) );
  OAI22_X1 U1662 ( .A1(n4849), .A2(n6368), .B1(n185), .B2(n251), .ZN(n3903) );
  OAI22_X1 U1663 ( .A1(n4817), .A2(n6367), .B1(n185), .B2(n253), .ZN(n3904) );
  OAI22_X1 U1664 ( .A1(n4785), .A2(n6364), .B1(n185), .B2(n255), .ZN(n3905) );
  OAI22_X1 U1665 ( .A1(n4753), .A2(n6362), .B1(n185), .B2(n257), .ZN(n3906) );
  OAI22_X1 U1666 ( .A1(n4721), .A2(n6361), .B1(n185), .B2(n259), .ZN(n3907) );
  OAI22_X1 U1667 ( .A1(n4689), .A2(n6365), .B1(n185), .B2(n261), .ZN(n3908) );
  OAI22_X1 U1668 ( .A1(n4657), .A2(n6366), .B1(n185), .B2(n263), .ZN(n3909) );
  OAI22_X1 U1669 ( .A1(n4625), .A2(n6369), .B1(n185), .B2(n265), .ZN(n3910) );
  OAI22_X1 U1670 ( .A1(n4593), .A2(n6370), .B1(n185), .B2(n267), .ZN(n3911) );
  OAI22_X1 U1671 ( .A1(n4561), .A2(n6373), .B1(n185), .B2(n269), .ZN(n3912) );
  OAI22_X1 U1672 ( .A1(n4529), .A2(n6374), .B1(n185), .B2(n271), .ZN(n3913) );
  OAI22_X1 U1673 ( .A1(n4497), .A2(n6377), .B1(n185), .B2(n273), .ZN(n3914) );
  OAI22_X1 U1674 ( .A1(n4465), .A2(n6378), .B1(n185), .B2(n275), .ZN(n3915) );
  OAI22_X1 U1675 ( .A1(n4433), .A2(n6381), .B1(n185), .B2(n277), .ZN(n3916) );
  OAI22_X1 U1676 ( .A1(n4401), .A2(n6384), .B1(n185), .B2(n279), .ZN(n3917) );
  OAI22_X1 U1677 ( .A1(n4369), .A2(n6383), .B1(n185), .B2(n281), .ZN(n3918) );
  OAI22_X1 U1678 ( .A1(n4337), .A2(n6391), .B1(n185), .B2(n283), .ZN(n3919) );
  OAI22_X1 U1680 ( .A1(n5296), .A2(n6393), .B1(n169), .B2(n223), .ZN(n3920) );
  OAI22_X1 U1681 ( .A1(n5264), .A2(n6396), .B1(n169), .B2(n225), .ZN(n3921) );
  OAI22_X1 U1682 ( .A1(n5232), .A2(n6387), .B1(n169), .B2(n227), .ZN(n3922) );
  OAI22_X1 U1683 ( .A1(n5200), .A2(n6395), .B1(n169), .B2(n229), .ZN(n3923) );
  OAI22_X1 U1684 ( .A1(n5168), .A2(n6390), .B1(n169), .B2(n231), .ZN(n3924) );
  OAI22_X1 U1685 ( .A1(n5136), .A2(n6385), .B1(n169), .B2(n233), .ZN(n3925) );
  OAI22_X1 U1686 ( .A1(n5104), .A2(n6389), .B1(n169), .B2(n235), .ZN(n3926) );
  OAI22_X1 U1687 ( .A1(n5072), .A2(n6382), .B1(n169), .B2(n237), .ZN(n3927) );
  OAI22_X1 U1688 ( .A1(n5040), .A2(n6380), .B1(n169), .B2(n239), .ZN(n3928) );
  OAI22_X1 U1689 ( .A1(n5008), .A2(n6379), .B1(n169), .B2(n241), .ZN(n3929) );
  OAI22_X1 U1690 ( .A1(n4976), .A2(n6376), .B1(n169), .B2(n243), .ZN(n3930) );
  OAI22_X1 U1691 ( .A1(n4944), .A2(n6375), .B1(n169), .B2(n245), .ZN(n3931) );
  OAI22_X1 U1692 ( .A1(n4912), .A2(n6372), .B1(n169), .B2(n247), .ZN(n3932) );
  OAI22_X1 U1693 ( .A1(n4880), .A2(n6371), .B1(n169), .B2(n249), .ZN(n3933) );
  OAI22_X1 U1694 ( .A1(n4848), .A2(n6368), .B1(n169), .B2(n251), .ZN(n3934) );
  OAI22_X1 U1695 ( .A1(n4816), .A2(n6367), .B1(n169), .B2(n253), .ZN(n3935) );
  OAI22_X1 U1696 ( .A1(n4784), .A2(n6364), .B1(n169), .B2(n255), .ZN(n3936) );
  OAI22_X1 U1697 ( .A1(n4752), .A2(n6362), .B1(n169), .B2(n257), .ZN(n3937) );
  OAI22_X1 U1698 ( .A1(n4720), .A2(n6361), .B1(n169), .B2(n259), .ZN(n3938) );
  OAI22_X1 U1699 ( .A1(n4688), .A2(n6365), .B1(n169), .B2(n261), .ZN(n3939) );
  OAI22_X1 U1700 ( .A1(n4656), .A2(n6366), .B1(n169), .B2(n263), .ZN(n3940) );
  OAI22_X1 U1701 ( .A1(n4624), .A2(n6369), .B1(n169), .B2(n265), .ZN(n3941) );
  OAI22_X1 U1702 ( .A1(n4592), .A2(n6370), .B1(n169), .B2(n267), .ZN(n3942) );
  OAI22_X1 U1703 ( .A1(n4560), .A2(n6373), .B1(n169), .B2(n269), .ZN(n3943) );
  OAI22_X1 U1704 ( .A1(n4528), .A2(n6374), .B1(n169), .B2(n271), .ZN(n3944) );
  OAI22_X1 U1705 ( .A1(n4496), .A2(n6377), .B1(n169), .B2(n273), .ZN(n3945) );
  OAI22_X1 U1706 ( .A1(n4464), .A2(n6378), .B1(n169), .B2(n275), .ZN(n3946) );
  OAI22_X1 U1707 ( .A1(n4432), .A2(n6381), .B1(n169), .B2(n277), .ZN(n3947) );
  OAI22_X1 U1708 ( .A1(n4400), .A2(n6384), .B1(n169), .B2(n279), .ZN(n3948) );
  OAI22_X1 U1709 ( .A1(n4368), .A2(n6383), .B1(n169), .B2(n281), .ZN(n3949) );
  OAI22_X1 U1710 ( .A1(n4336), .A2(n6391), .B1(n169), .B2(n283), .ZN(n3950) );
  OAI22_X1 U1712 ( .A1(n5295), .A2(n6393), .B1(n152), .B2(n223), .ZN(n3951) );
  OAI22_X1 U1713 ( .A1(n5263), .A2(n6396), .B1(n152), .B2(n225), .ZN(n3952) );
  OAI22_X1 U1714 ( .A1(n5231), .A2(n6387), .B1(n152), .B2(n227), .ZN(n3953) );
  OAI22_X1 U1715 ( .A1(n5199), .A2(n6395), .B1(n152), .B2(n229), .ZN(n3954) );
  OAI22_X1 U1716 ( .A1(n5167), .A2(n6390), .B1(n152), .B2(n231), .ZN(n3955) );
  OAI22_X1 U1717 ( .A1(n5135), .A2(n6385), .B1(n152), .B2(n233), .ZN(n3956) );
  OAI22_X1 U1718 ( .A1(n5103), .A2(n6389), .B1(n152), .B2(n235), .ZN(n3957) );
  OAI22_X1 U1719 ( .A1(n5071), .A2(n6382), .B1(n152), .B2(n237), .ZN(n3958) );
  OAI22_X1 U1720 ( .A1(n5039), .A2(n6380), .B1(n152), .B2(n239), .ZN(n3959) );
  OAI22_X1 U1721 ( .A1(n5007), .A2(n6379), .B1(n152), .B2(n241), .ZN(n3960) );
  OAI22_X1 U1722 ( .A1(n4975), .A2(n6376), .B1(n152), .B2(n243), .ZN(n3961) );
  OAI22_X1 U1723 ( .A1(n4943), .A2(n6375), .B1(n152), .B2(n245), .ZN(n3962) );
  OAI22_X1 U1724 ( .A1(n4911), .A2(n6372), .B1(n152), .B2(n247), .ZN(n3963) );
  OAI22_X1 U1725 ( .A1(n4879), .A2(n6371), .B1(n152), .B2(n249), .ZN(n3964) );
  OAI22_X1 U1726 ( .A1(n4847), .A2(n6368), .B1(n152), .B2(n251), .ZN(n3965) );
  OAI22_X1 U1727 ( .A1(n4815), .A2(n6367), .B1(n152), .B2(n253), .ZN(n3966) );
  OAI22_X1 U1728 ( .A1(n4783), .A2(n6364), .B1(n152), .B2(n255), .ZN(n3967) );
  OAI22_X1 U1729 ( .A1(n4751), .A2(n6362), .B1(n152), .B2(n257), .ZN(n3968) );
  OAI22_X1 U1730 ( .A1(n4719), .A2(n6361), .B1(n152), .B2(n259), .ZN(n3969) );
  OAI22_X1 U1731 ( .A1(n4687), .A2(n6365), .B1(n152), .B2(n261), .ZN(n3970) );
  OAI22_X1 U1732 ( .A1(n4655), .A2(n6366), .B1(n152), .B2(n263), .ZN(n3971) );
  OAI22_X1 U1733 ( .A1(n4623), .A2(n6369), .B1(n152), .B2(n265), .ZN(n3972) );
  OAI22_X1 U1734 ( .A1(n4591), .A2(n6370), .B1(n152), .B2(n267), .ZN(n3973) );
  OAI22_X1 U1735 ( .A1(n4559), .A2(n6373), .B1(n152), .B2(n269), .ZN(n3974) );
  OAI22_X1 U1736 ( .A1(n4527), .A2(n6374), .B1(n152), .B2(n271), .ZN(n3975) );
  OAI22_X1 U1737 ( .A1(n4495), .A2(n6377), .B1(n152), .B2(n273), .ZN(n3976) );
  OAI22_X1 U1738 ( .A1(n4463), .A2(n6378), .B1(n152), .B2(n275), .ZN(n3977) );
  OAI22_X1 U1739 ( .A1(n4431), .A2(n6381), .B1(n152), .B2(n277), .ZN(n3978) );
  OAI22_X1 U1740 ( .A1(n4399), .A2(n6384), .B1(n152), .B2(n279), .ZN(n3979) );
  OAI22_X1 U1741 ( .A1(n4367), .A2(n6383), .B1(n152), .B2(n281), .ZN(n3980) );
  OAI22_X1 U1742 ( .A1(n4335), .A2(n6391), .B1(n152), .B2(n283), .ZN(n3981) );
  OAI22_X1 U1744 ( .A1(n5294), .A2(n6393), .B1(n135), .B2(n223), .ZN(n3982) );
  OAI22_X1 U1745 ( .A1(n5262), .A2(n6396), .B1(n135), .B2(n225), .ZN(n3983) );
  OAI22_X1 U1746 ( .A1(n5230), .A2(n6387), .B1(n135), .B2(n227), .ZN(n3984) );
  OAI22_X1 U1747 ( .A1(n5198), .A2(n6395), .B1(n135), .B2(n229), .ZN(n3985) );
  OAI22_X1 U1748 ( .A1(n5166), .A2(n6390), .B1(n135), .B2(n231), .ZN(n3986) );
  OAI22_X1 U1749 ( .A1(n5134), .A2(n6385), .B1(n135), .B2(n233), .ZN(n3987) );
  OAI22_X1 U1750 ( .A1(n5102), .A2(n6389), .B1(n135), .B2(n235), .ZN(n3988) );
  OAI22_X1 U1751 ( .A1(n5070), .A2(n6382), .B1(n135), .B2(n237), .ZN(n3989) );
  OAI22_X1 U1752 ( .A1(n5038), .A2(n6380), .B1(n135), .B2(n239), .ZN(n3990) );
  OAI22_X1 U1753 ( .A1(n5006), .A2(n6379), .B1(n135), .B2(n241), .ZN(n3991) );
  OAI22_X1 U1754 ( .A1(n4974), .A2(n6376), .B1(n135), .B2(n243), .ZN(n3992) );
  OAI22_X1 U1755 ( .A1(n4942), .A2(n6375), .B1(n135), .B2(n245), .ZN(n3993) );
  OAI22_X1 U1756 ( .A1(n4910), .A2(n6372), .B1(n135), .B2(n247), .ZN(n3994) );
  OAI22_X1 U1757 ( .A1(n4878), .A2(n6371), .B1(n135), .B2(n249), .ZN(n3995) );
  OAI22_X1 U1758 ( .A1(n4846), .A2(n6368), .B1(n135), .B2(n251), .ZN(n3996) );
  OAI22_X1 U1759 ( .A1(n4814), .A2(n6367), .B1(n135), .B2(n253), .ZN(n3997) );
  OAI22_X1 U1760 ( .A1(n4782), .A2(n6364), .B1(n135), .B2(n255), .ZN(n3998) );
  OAI22_X1 U1761 ( .A1(n4750), .A2(n6362), .B1(n135), .B2(n257), .ZN(n3999) );
  OAI22_X1 U1762 ( .A1(n4718), .A2(n6361), .B1(n135), .B2(n259), .ZN(n4000) );
  OAI22_X1 U1763 ( .A1(n4686), .A2(n6365), .B1(n135), .B2(n261), .ZN(n4001) );
  OAI22_X1 U1764 ( .A1(n4654), .A2(n6366), .B1(n135), .B2(n263), .ZN(n4002) );
  OAI22_X1 U1765 ( .A1(n4622), .A2(n6369), .B1(n135), .B2(n265), .ZN(n4003) );
  OAI22_X1 U1766 ( .A1(n4590), .A2(n6370), .B1(n135), .B2(n267), .ZN(n4004) );
  OAI22_X1 U1767 ( .A1(n4558), .A2(n6373), .B1(n135), .B2(n269), .ZN(n4005) );
  OAI22_X1 U1768 ( .A1(n4526), .A2(n6374), .B1(n135), .B2(n271), .ZN(n4006) );
  OAI22_X1 U1769 ( .A1(n4494), .A2(n6377), .B1(n135), .B2(n273), .ZN(n4007) );
  OAI22_X1 U1770 ( .A1(n4462), .A2(n6378), .B1(n135), .B2(n275), .ZN(n4008) );
  OAI22_X1 U1771 ( .A1(n4430), .A2(n6381), .B1(n135), .B2(n277), .ZN(n4009) );
  OAI22_X1 U1772 ( .A1(n4398), .A2(n6384), .B1(n135), .B2(n279), .ZN(n4010) );
  OAI22_X1 U1773 ( .A1(n4366), .A2(n6383), .B1(n135), .B2(n281), .ZN(n4011) );
  OAI22_X1 U1774 ( .A1(n4334), .A2(n6391), .B1(n135), .B2(n283), .ZN(n4012) );
  OAI22_X1 U1776 ( .A1(n5293), .A2(n6393), .B1(n114), .B2(n223), .ZN(n4013) );
  OAI22_X1 U1777 ( .A1(n5261), .A2(n6396), .B1(n114), .B2(n225), .ZN(n4014) );
  OAI22_X1 U1778 ( .A1(n5229), .A2(n6387), .B1(n114), .B2(n227), .ZN(n4015) );
  OAI22_X1 U1779 ( .A1(n5197), .A2(n6395), .B1(n114), .B2(n229), .ZN(n4016) );
  OAI22_X1 U1780 ( .A1(n5165), .A2(n6390), .B1(n114), .B2(n231), .ZN(n4017) );
  OAI22_X1 U1781 ( .A1(n5133), .A2(n6385), .B1(n114), .B2(n233), .ZN(n4018) );
  OAI22_X1 U1782 ( .A1(n5101), .A2(n6389), .B1(n114), .B2(n235), .ZN(n4019) );
  OAI22_X1 U1783 ( .A1(n5069), .A2(n6382), .B1(n114), .B2(n237), .ZN(n4020) );
  OAI22_X1 U1784 ( .A1(n5037), .A2(n6380), .B1(n114), .B2(n239), .ZN(n4021) );
  OAI22_X1 U1785 ( .A1(n5005), .A2(n6379), .B1(n114), .B2(n241), .ZN(n4022) );
  OAI22_X1 U1786 ( .A1(n4973), .A2(n6376), .B1(n114), .B2(n243), .ZN(n4023) );
  OAI22_X1 U1787 ( .A1(n4941), .A2(n6375), .B1(n114), .B2(n245), .ZN(n4024) );
  OAI22_X1 U1788 ( .A1(n4909), .A2(n6372), .B1(n114), .B2(n247), .ZN(n4025) );
  OAI22_X1 U1789 ( .A1(n4877), .A2(n6371), .B1(n114), .B2(n249), .ZN(n4026) );
  OAI22_X1 U1790 ( .A1(n4845), .A2(n6368), .B1(n114), .B2(n251), .ZN(n4027) );
  OAI22_X1 U1791 ( .A1(n4813), .A2(n6367), .B1(n114), .B2(n253), .ZN(n4028) );
  OAI22_X1 U1792 ( .A1(n4781), .A2(n6364), .B1(n114), .B2(n255), .ZN(n4029) );
  OAI22_X1 U1793 ( .A1(n4749), .A2(n6362), .B1(n114), .B2(n257), .ZN(n4030) );
  OAI22_X1 U1794 ( .A1(n4717), .A2(n6361), .B1(n114), .B2(n259), .ZN(n4031) );
  OAI22_X1 U1795 ( .A1(n4685), .A2(n6365), .B1(n114), .B2(n261), .ZN(n4032) );
  OAI22_X1 U1796 ( .A1(n4653), .A2(n6366), .B1(n114), .B2(n263), .ZN(n4033) );
  OAI22_X1 U1797 ( .A1(n4621), .A2(n6369), .B1(n114), .B2(n265), .ZN(n4034) );
  OAI22_X1 U1798 ( .A1(n4589), .A2(n6370), .B1(n114), .B2(n267), .ZN(n4035) );
  OAI22_X1 U1799 ( .A1(n4557), .A2(n6373), .B1(n114), .B2(n269), .ZN(n4036) );
  OAI22_X1 U1800 ( .A1(n4525), .A2(n6374), .B1(n114), .B2(n271), .ZN(n4037) );
  OAI22_X1 U1801 ( .A1(n4493), .A2(n6377), .B1(n114), .B2(n273), .ZN(n4038) );
  OAI22_X1 U1802 ( .A1(n4461), .A2(n6378), .B1(n114), .B2(n275), .ZN(n4039) );
  OAI22_X1 U1803 ( .A1(n4429), .A2(n6381), .B1(n114), .B2(n277), .ZN(n4040) );
  OAI22_X1 U1804 ( .A1(n4397), .A2(n6384), .B1(n114), .B2(n279), .ZN(n4041) );
  OAI22_X1 U1805 ( .A1(n4365), .A2(n6383), .B1(n114), .B2(n281), .ZN(n4042) );
  OAI22_X1 U1806 ( .A1(n4333), .A2(n6391), .B1(n114), .B2(n283), .ZN(n4043) );
  OAI22_X1 U1808 ( .A1(n5291), .A2(n6393), .B1(n100), .B2(n223), .ZN(n4044) );
  OAI22_X1 U1809 ( .A1(n5259), .A2(n6396), .B1(n100), .B2(n225), .ZN(n4045) );
  OAI22_X1 U1810 ( .A1(n5227), .A2(n6387), .B1(n100), .B2(n227), .ZN(n4046) );
  OAI22_X1 U1811 ( .A1(n5195), .A2(n6395), .B1(n100), .B2(n229), .ZN(n4047) );
  OAI22_X1 U1812 ( .A1(n5163), .A2(n6390), .B1(n100), .B2(n231), .ZN(n4048) );
  OAI22_X1 U1813 ( .A1(n5131), .A2(n6385), .B1(n100), .B2(n233), .ZN(n4049) );
  OAI22_X1 U1814 ( .A1(n5099), .A2(n6389), .B1(n100), .B2(n235), .ZN(n4050) );
  OAI22_X1 U1815 ( .A1(n5067), .A2(n6382), .B1(n100), .B2(n237), .ZN(n4051) );
  OAI22_X1 U1816 ( .A1(n5035), .A2(n6380), .B1(n100), .B2(n239), .ZN(n4052) );
  OAI22_X1 U1817 ( .A1(n5003), .A2(n6379), .B1(n100), .B2(n241), .ZN(n4053) );
  OAI22_X1 U1818 ( .A1(n4971), .A2(n6376), .B1(n100), .B2(n243), .ZN(n4054) );
  OAI22_X1 U1819 ( .A1(n4939), .A2(n6375), .B1(n100), .B2(n245), .ZN(n4055) );
  OAI22_X1 U1820 ( .A1(n4907), .A2(n6372), .B1(n100), .B2(n247), .ZN(n4056) );
  OAI22_X1 U1821 ( .A1(n4875), .A2(n6371), .B1(n100), .B2(n249), .ZN(n4057) );
  OAI22_X1 U1822 ( .A1(n4843), .A2(n6368), .B1(n100), .B2(n251), .ZN(n4058) );
  OAI22_X1 U1823 ( .A1(n4811), .A2(n6367), .B1(n100), .B2(n253), .ZN(n4059) );
  OAI22_X1 U1824 ( .A1(n4779), .A2(n6364), .B1(n100), .B2(n255), .ZN(n4060) );
  OAI22_X1 U1825 ( .A1(n4747), .A2(n6362), .B1(n100), .B2(n257), .ZN(n4061) );
  OAI22_X1 U1826 ( .A1(n4715), .A2(n6361), .B1(n100), .B2(n259), .ZN(n4062) );
  OAI22_X1 U1827 ( .A1(n4683), .A2(n6365), .B1(n100), .B2(n261), .ZN(n4063) );
  OAI22_X1 U1828 ( .A1(n4651), .A2(n6366), .B1(n100), .B2(n263), .ZN(n4064) );
  OAI22_X1 U1829 ( .A1(n4619), .A2(n6369), .B1(n100), .B2(n265), .ZN(n4065) );
  OAI22_X1 U1830 ( .A1(n4587), .A2(n6370), .B1(n100), .B2(n267), .ZN(n4066) );
  OAI22_X1 U1831 ( .A1(n4555), .A2(n6373), .B1(n100), .B2(n269), .ZN(n4067) );
  OAI22_X1 U1832 ( .A1(n4523), .A2(n6374), .B1(n100), .B2(n271), .ZN(n4068) );
  OAI22_X1 U1833 ( .A1(n4491), .A2(n6377), .B1(n100), .B2(n273), .ZN(n4069) );
  OAI22_X1 U1834 ( .A1(n4459), .A2(n6378), .B1(n100), .B2(n275), .ZN(n4070) );
  OAI22_X1 U1835 ( .A1(n4427), .A2(n6381), .B1(n100), .B2(n277), .ZN(n4071) );
  OAI22_X1 U1836 ( .A1(n4395), .A2(n6384), .B1(n100), .B2(n279), .ZN(n4072) );
  OAI22_X1 U1837 ( .A1(n4363), .A2(n6383), .B1(n100), .B2(n281), .ZN(n4073) );
  OAI22_X1 U1838 ( .A1(n4331), .A2(n6391), .B1(n100), .B2(n283), .ZN(n4074) );
  OAI221_X1 U1840 ( .B1(n115), .B2(n873), .C1(n5541), .C2(n117), .A(n874), 
        .ZN(n4075) );
  AOI22_X1 U1841 ( .A1(n119), .A2(n108), .B1(\UUT/Mpath/the_mult/Mad_out [31]), 
        .B2(n121), .ZN(n874) );
  OAI22_X1 U1843 ( .A1(n7382), .A2(n875), .B1(n5542), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4076) );
  OAI221_X1 U1844 ( .B1(n5316), .B2(n124), .C1(n125), .C2(n875), .A(n876), 
        .ZN(n4077) );
  AOI22_X1 U1845 ( .A1(n127), .A2(n877), .B1(n129), .B2(n878), .ZN(n876) );
  INV_X1 U1846 ( .A(\UUT/Mpath/the_mult/x_operand1[31] ), .ZN(n875) );
  OAI221_X1 U1847 ( .B1(n5316), .B2(n218), .C1(\UUT/Mpath/the_alu/N21 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n879), .ZN(n4078) );
  AOI22_X1 U1848 ( .A1(n220), .A2(n877), .B1(n221), .B2(n878), .ZN(n879) );
  OAI22_X1 U1849 ( .A1(n5290), .A2(n6393), .B1(n880), .B2(n223), .ZN(n4079) );
  OAI22_X1 U1852 ( .A1(n5258), .A2(n224), .B1(n880), .B2(n225), .ZN(n4080) );
  NOR3_X1 U1854 ( .A1(\UUT/regfile/N336 ), .A2(n7391), .A3(n882), .ZN(n224) );
  OAI22_X1 U1855 ( .A1(n5226), .A2(n6387), .B1(n880), .B2(n227), .ZN(n4081) );
  OAI22_X1 U1858 ( .A1(n5194), .A2(n6395), .B1(n880), .B2(n229), .ZN(n4082) );
  OAI22_X1 U1861 ( .A1(n5162), .A2(n230), .B1(n880), .B2(n231), .ZN(n4083) );
  NOR3_X1 U1863 ( .A1(\UUT/regfile/N354 ), .A2(n7391), .A3(n881), .ZN(n230) );
  OAI22_X1 U1864 ( .A1(n5130), .A2(n232), .B1(n880), .B2(n233), .ZN(n4084) );
  NOR3_X1 U1866 ( .A1(\UUT/regfile/N360 ), .A2(n7391), .A3(n882), .ZN(n232) );
  OAI22_X1 U1867 ( .A1(n5098), .A2(n6389), .B1(n880), .B2(n235), .ZN(n4085) );
  OAI22_X1 U1870 ( .A1(n5066), .A2(n236), .B1(n880), .B2(n237), .ZN(n4086) );
  NOR3_X1 U1872 ( .A1(\UUT/regfile/N373 ), .A2(n7391), .A3(n884), .ZN(n236) );
  OAI22_X1 U1873 ( .A1(n5034), .A2(n238), .B1(n880), .B2(n239), .ZN(n4087) );
  NOR3_X1 U1875 ( .A1(\UUT/regfile/N379 ), .A2(n7392), .A3(n881), .ZN(n238) );
  OAI22_X1 U1876 ( .A1(n5002), .A2(n240), .B1(n880), .B2(n241), .ZN(n4088) );
  NOR3_X1 U1878 ( .A1(\UUT/regfile/N385 ), .A2(n7392), .A3(n882), .ZN(n240) );
  OAI22_X1 U1879 ( .A1(n4970), .A2(n242), .B1(n880), .B2(n243), .ZN(n4089) );
  NOR3_X1 U1881 ( .A1(\UUT/regfile/N273 ), .A2(n7392), .A3(n884), .ZN(n242) );
  OAI22_X1 U1882 ( .A1(n4938), .A2(n244), .B1(n880), .B2(n245), .ZN(n4090) );
  NOR3_X1 U1884 ( .A1(\UUT/regfile/N391 ), .A2(n7392), .A3(n883), .ZN(n244) );
  OAI22_X1 U1885 ( .A1(n4906), .A2(n246), .B1(n880), .B2(n247), .ZN(n4091) );
  NOR3_X1 U1887 ( .A1(\UUT/regfile/N397 ), .A2(n7392), .A3(n884), .ZN(n246) );
  OAI22_X1 U1888 ( .A1(n4874), .A2(n248), .B1(n880), .B2(n249), .ZN(n4092) );
  NOR3_X1 U1890 ( .A1(\UUT/regfile/N403 ), .A2(n7392), .A3(n881), .ZN(n248) );
  OAI22_X1 U1891 ( .A1(n4842), .A2(n250), .B1(n880), .B2(n251), .ZN(n4093) );
  NOR3_X1 U1893 ( .A1(\UUT/regfile/N409 ), .A2(n7392), .A3(n882), .ZN(n250) );
  OAI22_X1 U1894 ( .A1(n4810), .A2(n252), .B1(n880), .B2(n253), .ZN(n4094) );
  NOR3_X1 U1896 ( .A1(\UUT/regfile/N415 ), .A2(n7392), .A3(n883), .ZN(n252) );
  OAI22_X1 U1897 ( .A1(n4778), .A2(n6364), .B1(n880), .B2(n255), .ZN(n4095) );
  OAI22_X1 U1900 ( .A1(n4746), .A2(n256), .B1(n880), .B2(n257), .ZN(n4096) );
  NOR3_X1 U1902 ( .A1(\UUT/regfile/N427 ), .A2(n7392), .A3(n881), .ZN(n256) );
  OAI22_X1 U1903 ( .A1(n4714), .A2(n6361), .B1(n880), .B2(n259), .ZN(n4097) );
  OAI22_X1 U1906 ( .A1(n4682), .A2(n260), .B1(n880), .B2(n261), .ZN(n4098) );
  NOR3_X1 U1908 ( .A1(\UUT/regfile/N439 ), .A2(n7392), .A3(n883), .ZN(n260) );
  OAI22_X1 U1909 ( .A1(n4650), .A2(n262), .B1(n880), .B2(n263), .ZN(n4099) );
  NOR3_X1 U1911 ( .A1(\UUT/regfile/N445 ), .A2(n7393), .A3(n884), .ZN(n262) );
  OAI22_X1 U1912 ( .A1(n4618), .A2(n264), .B1(n880), .B2(n265), .ZN(n4100) );
  NOR3_X1 U1914 ( .A1(\UUT/regfile/N280 ), .A2(n7393), .A3(n881), .ZN(n264) );
  OAI22_X1 U1915 ( .A1(n4586), .A2(n266), .B1(n880), .B2(n267), .ZN(n4101) );
  NOR3_X1 U1917 ( .A1(\UUT/regfile/N451 ), .A2(n7393), .A3(n881), .ZN(n266) );
  OAI22_X1 U1918 ( .A1(n4554), .A2(n268), .B1(n880), .B2(n269), .ZN(n4102) );
  NOR3_X1 U1920 ( .A1(\UUT/regfile/N457 ), .A2(n7393), .A3(n882), .ZN(n268) );
  OAI22_X1 U1921 ( .A1(n4522), .A2(n270), .B1(n880), .B2(n271), .ZN(n4103) );
  NOR3_X1 U1923 ( .A1(\UUT/regfile/N286 ), .A2(n7393), .A3(n882), .ZN(n270) );
  OAI22_X1 U1924 ( .A1(n4490), .A2(n272), .B1(n880), .B2(n273), .ZN(n4104) );
  NOR3_X1 U1926 ( .A1(\UUT/regfile/N293 ), .A2(n7393), .A3(n883), .ZN(n272) );
  OAI22_X1 U1927 ( .A1(n4458), .A2(n274), .B1(n880), .B2(n275), .ZN(n4105) );
  NOR3_X1 U1929 ( .A1(\UUT/regfile/N299 ), .A2(n7393), .A3(n884), .ZN(n274) );
  OAI22_X1 U1930 ( .A1(n4426), .A2(n276), .B1(n880), .B2(n277), .ZN(n4106) );
  NOR3_X1 U1932 ( .A1(\UUT/regfile/N305 ), .A2(n7393), .A3(n881), .ZN(n276) );
  NAND2_X1 U1933 ( .A1(\UUT/rd_addr [1]), .A2(n885), .ZN(n881) );
  OAI22_X1 U1934 ( .A1(n4394), .A2(n278), .B1(n880), .B2(n279), .ZN(n4107) );
  NOR3_X1 U1936 ( .A1(\UUT/regfile/N311 ), .A2(n7393), .A3(n882), .ZN(n278) );
  NAND2_X1 U1937 ( .A1(n886), .A2(\UUT/rd_addr [1]), .ZN(n882) );
  OAI22_X1 U1938 ( .A1(n4362), .A2(n280), .B1(n880), .B2(n281), .ZN(n4108) );
  NOR3_X1 U1940 ( .A1(\UUT/regfile/N318 ), .A2(n7393), .A3(n883), .ZN(n280) );
  NAND2_X1 U1941 ( .A1(n887), .A2(n885), .ZN(n883) );
  OAI22_X1 U1942 ( .A1(n4330), .A2(n282), .B1(n880), .B2(n283), .ZN(n4109) );
  NOR3_X1 U1944 ( .A1(\UUT/regfile/N324 ), .A2(n7393), .A3(n884), .ZN(n282) );
  NAND2_X1 U1945 ( .A1(n886), .A2(n887), .ZN(n884) );
  INV_X1 U1946 ( .A(\UUT/rd_addr [1]), .ZN(n887) );
  INV_X1 U1947 ( .A(n885), .ZN(n886) );
  NAND2_X1 U1948 ( .A1(\UUT/Mcontrol/m_sampled_xrd[0] ), .A2(n5315), .ZN(n885)
         );
  OAI22_X1 U1949 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mpath/the_memhandle/N239 ), .B1(n888), .B2(n7394), .ZN(n4110) );
  INV_X1 U1950 ( .A(\UUT/daddr_out [1]), .ZN(n888) );
  OAI222_X1 U1951 ( .A1(n49), .A2(n94), .B1(n833), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N82 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n4111) );
  INV_X1 U1952 ( .A(\UUT/break_code[1] ), .ZN(n833) );
  INV_X1 U1953 ( .A(n889), .ZN(n49) );
  OAI222_X1 U1954 ( .A1(n890), .A2(n99), .B1(n859), .B2(n101), .C1(n5395), 
        .C2(n102), .ZN(n889) );
  OAI222_X1 U1956 ( .A1(n891), .A2(n692), .B1(n892), .B2(n827), .C1(n5623), 
        .C2(n5396), .ZN(n856) );
  AOI221_X1 U1957 ( .B1(\UUT/Mpath/the_memhandle/N36 ), .B2(n893), .C1(
        \UUT/Mpath/the_memhandle/N38 ), .C2(n643), .A(n5800), .ZN(n892) );
  INV_X1 U1958 ( .A(n5798), .ZN(n643) );
  INV_X1 U1959 ( .A(n5799), .ZN(n893) );
  AOI221_X1 U1960 ( .B1(D_DATA_INBUS[1]), .B2(n5663), .C1(D_DATA_INBUS[17]), 
        .C2(n5664), .A(n5797), .ZN(n891) );
  OAI22_X1 U1961 ( .A1(n5396), .A2(\UUT/Mcontrol/N22 ), .B1(n890), .B2(n7394), 
        .ZN(n4112) );
  INV_X1 U1962 ( .A(n857), .ZN(n890) );
  OAI211_X1 U1963 ( .C1(n5958), .C2(n287), .A(n894), .B(n895), .ZN(n857) );
  AOI222_X1 U1964 ( .A1(\UUT/Mpath/the_mult/x_mult_out[1] ), .A2(n6357), .B1(
        n320), .B2(n896), .C1(n291), .C2(n897), .ZN(n895) );
  INV_X1 U1965 ( .A(n5611), .ZN(n897) );
  AOI22_X1 U1967 ( .A1(n6397), .A2(n898), .B1(n324), .B2(\UUT/daddr_out [1]), 
        .ZN(n894) );
  INV_X1 U1968 ( .A(n5567), .ZN(n898) );
  OAI221_X1 U1969 ( .B1(n5322), .B2(n218), .C1(\UUT/Mpath/the_alu/N33 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n899), .ZN(n4113) );
  AOI22_X1 U1970 ( .A1(n220), .A2(n193), .B1(n221), .B2(n194), .ZN(n899) );
  OAI221_X1 U1971 ( .B1(n5799), .B2(n284), .C1(n5623), .C2(n5378), .A(n285), 
        .ZN(n193) );
  OAI22_X1 U1972 ( .A1(n5378), .A2(\UUT/Mcontrol/N22 ), .B1(n184), .B2(n7394), 
        .ZN(n4114) );
  OAI221_X1 U1974 ( .B1(n5508), .B2(n286), .C1(n5507), .C2(n287), .A(n900), 
        .ZN(n194) );
  INV_X1 U1976 ( .A(n5605), .ZN(n902) );
  INV_X1 U1977 ( .A(n5555), .ZN(n901) );
  OAI221_X1 U1978 ( .B1(n5321), .B2(n218), .C1(\UUT/Mpath/the_alu/N31 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n903), .ZN(n4115) );
  AOI22_X1 U1979 ( .A1(n220), .A2(n177), .B1(n221), .B2(n178), .ZN(n903) );
  OAI221_X1 U1980 ( .B1(n5728), .B2(n284), .C1(n5623), .C2(n5375), .A(n285), 
        .ZN(n177) );
  OAI22_X1 U1981 ( .A1(n5375), .A2(\UUT/Mcontrol/N22 ), .B1(n168), .B2(n7394), 
        .ZN(n4116) );
  INV_X1 U1985 ( .A(n5604), .ZN(n906) );
  INV_X1 U1986 ( .A(n5553), .ZN(n905) );
  OAI221_X1 U1987 ( .B1(n5320), .B2(n218), .C1(\UUT/Mpath/the_alu/N29 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n907), .ZN(n4117) );
  AOI22_X1 U1988 ( .A1(n220), .A2(n160), .B1(n221), .B2(n161), .ZN(n907) );
  OAI221_X1 U1989 ( .B1(n5707), .B2(n284), .C1(n5623), .C2(n5372), .A(n285), 
        .ZN(n160) );
  OAI22_X1 U1990 ( .A1(n5372), .A2(\UUT/Mcontrol/N22 ), .B1(n151), .B2(n7394), 
        .ZN(n4118) );
  INV_X1 U1994 ( .A(n5603), .ZN(n910) );
  INV_X1 U1995 ( .A(n5551), .ZN(n909) );
  OAI221_X1 U1996 ( .B1(n5319), .B2(n218), .C1(\UUT/Mpath/the_alu/N27 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n911), .ZN(n4119) );
  AOI22_X1 U1997 ( .A1(n220), .A2(n143), .B1(n221), .B2(n144), .ZN(n911) );
  OAI221_X1 U1998 ( .B1(n5697), .B2(n284), .C1(n5623), .C2(n5369), .A(n285), 
        .ZN(n143) );
  OAI22_X1 U1999 ( .A1(n5369), .A2(\UUT/Mcontrol/N22 ), .B1(n134), .B2(n7394), 
        .ZN(n4120) );
  INV_X1 U2003 ( .A(n5602), .ZN(n914) );
  INV_X1 U2004 ( .A(n5549), .ZN(n913) );
  OAI221_X1 U2005 ( .B1(n5318), .B2(n218), .C1(\UUT/Mpath/the_alu/N25 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n915), .ZN(n4121) );
  AOI22_X1 U2006 ( .A1(n220), .A2(n128), .B1(n221), .B2(n130), .ZN(n915) );
  OAI221_X1 U2007 ( .B1(n5687), .B2(n284), .C1(n5623), .C2(n5366), .A(n285), 
        .ZN(n128) );
  OAI22_X1 U2008 ( .A1(n5366), .A2(\UUT/Mcontrol/N22 ), .B1(n113), .B2(n7395), 
        .ZN(n4122) );
  OAI221_X1 U2010 ( .B1(n5476), .B2(n286), .C1(n5475), .C2(n287), .A(n916), 
        .ZN(n130) );
  INV_X1 U2012 ( .A(n5601), .ZN(n918) );
  INV_X1 U2013 ( .A(n5547), .ZN(n917) );
  OAI221_X1 U2014 ( .B1(n103), .B2(n919), .C1(n5601), .C2(n105), .A(n920), 
        .ZN(n4123) );
  AOI22_X1 U2015 ( .A1(n107), .A2(n120), .B1(\UUT/Mpath/the_mult/Mad_out [61]), 
        .B2(n109), .ZN(n920) );
  OAI221_X1 U2017 ( .B1(n115), .B2(n921), .C1(n5543), .C2(n117), .A(n922), 
        .ZN(n4124) );
  AOI22_X1 U2018 ( .A1(n119), .A2(n923), .B1(\UUT/Mpath/the_mult/Mad_out [30]), 
        .B2(n121), .ZN(n922) );
  NOR2_X1 U2020 ( .A1(n926), .A2(n927), .ZN(n925) );
  INV_X1 U2022 ( .A(\UUT/Mpath/the_mult/N255 ), .ZN(n926) );
  NAND3_X1 U2024 ( .A1(n924), .A2(n927), .A3(\UUT/Mpath/the_mult/N255 ), .ZN(
        n929) );
  INV_X1 U2025 ( .A(\UUT/Mpath/the_mult/N312 ), .ZN(n927) );
  INV_X1 U2026 ( .A(\UUT/Mpath/the_mult/N311 ), .ZN(n924) );
  OAI221_X1 U2028 ( .B1(n103), .B2(n930), .C1(n5599), .C2(n105), .A(n931), 
        .ZN(n4125) );
  AOI22_X1 U2029 ( .A1(n107), .A2(n923), .B1(\UUT/Mpath/the_mult/Mad_out [62]), 
        .B2(n109), .ZN(n931) );
  NOR2_X1 U2031 ( .A1(n934), .A2(n935), .ZN(n933) );
  INV_X1 U2034 ( .A(\UUT/Mpath/the_mult/N285 ), .ZN(n934) );
  NAND3_X1 U2036 ( .A1(n932), .A2(n935), .A3(\UUT/Mpath/the_mult/N285 ), .ZN(
        n936) );
  INV_X1 U2037 ( .A(\UUT/Mpath/the_mult/N314 ), .ZN(n935) );
  INV_X1 U2038 ( .A(\UUT/Mpath/the_mult/N313 ), .ZN(n932) );
  AND2_X1 U2040 ( .A1(n5315), .A2(\UUT/Mcontrol/N22 ), .ZN(n928) );
  OAI22_X1 U2041 ( .A1(n7383), .A2(n937), .B1(n5544), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4126) );
  OAI221_X1 U2042 ( .B1(n5317), .B2(n6350), .C1(n125), .C2(n937), .A(n938), 
        .ZN(n4127) );
  AOI22_X1 U2043 ( .A1(n127), .A2(n872), .B1(n129), .B2(n939), .ZN(n938) );
  INV_X1 U2046 ( .A(\UUT/Mpath/the_mult/x_operand1[30] ), .ZN(n937) );
  NAND2_X1 U2047 ( .A1(n125), .A2(n940), .ZN(n124) );
  OAI221_X1 U2050 ( .B1(n5317), .B2(n218), .C1(\UUT/Mpath/the_alu/N23 ), .C2(
        \UUT/Mcontrol/N22 ), .A(n941), .ZN(n4128) );
  AOI22_X1 U2051 ( .A1(n220), .A2(n872), .B1(n221), .B2(n939), .ZN(n941) );
  OAI221_X1 U2053 ( .B1(n5677), .B2(n284), .C1(n5623), .C2(n5360), .A(n285), 
        .ZN(n872) );
  OAI22_X1 U2056 ( .A1(n5360), .A2(\UUT/Mcontrol/N22 ), .B1(n98), .B2(n7395), 
        .ZN(n4129) );
  INV_X1 U2057 ( .A(n939), .ZN(n98) );
  INV_X1 U2060 ( .A(n5599), .ZN(n944) );
  INV_X1 U2061 ( .A(n5543), .ZN(n943) );
  OAI222_X1 U2062 ( .A1(n87), .A2(n7398), .B1(n86), .B2(n94), .C1(
        \UUT/Mpath/the_alu/N22 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n4130) );
  AND3_X1 U2063 ( .A1(n945), .A2(n150), .A3(n204), .ZN(n87) );
  AOI21_X1 U2064 ( .B1(n5752), .B2(n205), .A(n456), .ZN(n204) );
  NAND2_X1 U2065 ( .A1(n5751), .A2(n205), .ZN(n150) );
  NOR2_X1 U2066 ( .A1(n203), .A2(n946), .ZN(n205) );
  INV_X1 U2067 ( .A(n198), .ZN(n203) );
  NAND3_X1 U2068 ( .A1(n946), .A2(\UUT/Mcontrol/d_sampled_finstr [15]), .A3(
        n198), .ZN(n945) );
  NOR2_X1 U2069 ( .A1(n835), .A2(n947), .ZN(n198) );
  OAI22_X1 U2070 ( .A1(n5357), .A2(\UUT/Mcontrol/N22 ), .B1(n948), .B2(n7395), 
        .ZN(n4131) );
  OAI222_X1 U2071 ( .A1(n71), .A2(n94), .B1(n84), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N38 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n4132) );
  INV_X1 U2072 ( .A(n949), .ZN(n71) );
  OAI222_X1 U2073 ( .A1(n950), .A2(n99), .B1(n871), .B2(n101), .C1(n5383), 
        .C2(n102), .ZN(n949) );
  OAI221_X1 U2075 ( .B1(n951), .B2(n284), .C1(n5623), .C2(n5384), .A(n285), 
        .ZN(n868) );
  INV_X1 U2076 ( .A(D_DATA_INBUS[23]), .ZN(n951) );
  OAI22_X1 U2077 ( .A1(n5384), .A2(\UUT/Mcontrol/N22 ), .B1(n950), .B2(n7395), 
        .ZN(n4133) );
  INV_X1 U2078 ( .A(n869), .ZN(n950) );
  OAI211_X1 U2079 ( .C1(n5969), .C2(n287), .A(n952), .B(n953), .ZN(n869) );
  AOI222_X1 U2080 ( .A1(\UUT/Mpath/the_mult/x_mult_out[23] ), .A2(n6357), .B1(
        n320), .B2(n954), .C1(n291), .C2(n955), .ZN(n953) );
  INV_X1 U2081 ( .A(n5607), .ZN(n955) );
  AOI22_X1 U2083 ( .A1(n6397), .A2(n956), .B1(n324), .B2(n6114), .ZN(n952) );
  INV_X1 U2084 ( .A(n5559), .ZN(n956) );
  OAI22_X1 U2085 ( .A1(n7383), .A2(n957), .B1(n5968), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4134) );
  INV_X1 U2086 ( .A(\UUT/jar_in [23]), .ZN(n957) );
  OAI22_X1 U2087 ( .A1(n7383), .A2(n958), .B1(n5979), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4135) );
  INV_X1 U2088 ( .A(\UUT/jar_in [22]), .ZN(n958) );
  OAI22_X1 U2089 ( .A1(n7383), .A2(n959), .B1(n5989), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4136) );
  INV_X1 U2090 ( .A(\UUT/jar_in [21]), .ZN(n959) );
  OAI22_X1 U2091 ( .A1(n7384), .A2(n960), .B1(n5999), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4137) );
  INV_X1 U2092 ( .A(\UUT/jar_in [20]), .ZN(n960) );
  OAI22_X1 U2093 ( .A1(n7383), .A2(n961), .B1(n6012), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4138) );
  INV_X1 U2094 ( .A(\UUT/jar_in [19]), .ZN(n961) );
  OAI22_X1 U2095 ( .A1(n7384), .A2(n962), .B1(n6025), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4139) );
  INV_X1 U2096 ( .A(\UUT/jar_in [18]), .ZN(n962) );
  OAI22_X1 U2097 ( .A1(n7384), .A2(n963), .B1(n6046), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4140) );
  INV_X1 U2098 ( .A(\UUT/jar_in [17]), .ZN(n963) );
  OAI22_X1 U2099 ( .A1(n7384), .A2(n964), .B1(n6058), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4141) );
  INV_X1 U2100 ( .A(\UUT/jar_in [16]), .ZN(n964) );
  OAI22_X1 U2101 ( .A1(n7384), .A2(n965), .B1(n6069), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4142) );
  INV_X1 U2102 ( .A(\UUT/jar_in [15]), .ZN(n965) );
  OAI22_X1 U2103 ( .A1(n7384), .A2(n966), .B1(n6083), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4143) );
  INV_X1 U2104 ( .A(\UUT/jar_in [14]), .ZN(n966) );
  OAI22_X1 U2105 ( .A1(n7384), .A2(n967), .B1(n6093), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4144) );
  INV_X1 U2106 ( .A(\UUT/jar_in [13]), .ZN(n967) );
  OAI22_X1 U2107 ( .A1(n7384), .A2(n968), .B1(n6223), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4145) );
  OAI22_X1 U2108 ( .A1(n7384), .A2(n969), .B1(n6232), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4146) );
  OAI22_X1 U2109 ( .A1(n7384), .A2(n970), .B1(n6241), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4147) );
  OAI22_X1 U2110 ( .A1(n7386), .A2(n971), .B1(n6143), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4148) );
  OAI22_X1 U2111 ( .A1(n7385), .A2(n972), .B1(n6152), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4149) );
  OAI22_X1 U2112 ( .A1(n7384), .A2(n973), .B1(n6161), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4150) );
  OAI22_X1 U2113 ( .A1(n7385), .A2(n974), .B1(n6170), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4151) );
  OAI22_X1 U2114 ( .A1(n7385), .A2(n975), .B1(n6179), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4152) );
  OAI22_X1 U2115 ( .A1(n7385), .A2(n976), .B1(n6188), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4153) );
  OAI22_X1 U2116 ( .A1(n7385), .A2(n977), .B1(n6200), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4154) );
  OAI22_X1 U2117 ( .A1(n7385), .A2(n978), .B1(n6211), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4155) );
  OAI22_X1 U2118 ( .A1(n7385), .A2(n979), .B1(n5957), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4156) );
  INV_X1 U2119 ( .A(\UUT/jar_in [1]), .ZN(n979) );
  OAI221_X1 U2120 ( .B1(n79), .B2(n296), .C1(n297), .C2(n2709), .A(n980), .ZN(
        n4157) );
  AOI22_X1 U2121 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [0]), .A2(n301), .B1(
        \UUT/jar_in [0]), .B2(n6867), .ZN(n980) );
  OAI22_X1 U2122 ( .A1(n7385), .A2(n981), .B1(n5524), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4158) );
  INV_X1 U2123 ( .A(\UUT/jar_in [0]), .ZN(n981) );
  NAND2_X1 U2129 ( .A1(n985), .A2(n297), .ZN(n296) );
  OAI22_X1 U2130 ( .A1(n986), .A2(n556), .B1(n297), .B2(n2711), .ZN(n4160) );
  INV_X1 U2131 ( .A(\UUT/Mcontrol/Program_counter/N24 ), .ZN(n986) );
  OAI22_X1 U2132 ( .A1(\UUT/Mpath/the_memhandle/N240 ), .A2(\UUT/Mcontrol/N22 ), .B1(n987), .B2(n7395), .ZN(n4161) );
  INV_X1 U2133 ( .A(\UUT/daddr_out [0]), .ZN(n987) );
  OAI222_X1 U2134 ( .A1(n47), .A2(n94), .B1(n79), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N84 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n4162) );
  INV_X1 U2135 ( .A(n457), .ZN(n302) );
  NOR2_X1 U2136 ( .A1(n835), .A2(n7393), .ZN(n457) );
  INV_X1 U2137 ( .A(n6966), .ZN(n79) );
  OAI21_X1 U2139 ( .B1(n6131), .B2(n6071), .A(n5900), .ZN(n835) );
  INV_X1 U2140 ( .A(n988), .ZN(n47) );
  OAI222_X1 U2141 ( .A1(n989), .A2(n5332), .B1(n847), .B2(n101), .C1(n5428), 
        .C2(n102), .ZN(n988) );
  OAI222_X1 U2143 ( .A1(n990), .A2(n692), .B1(n991), .B2(n827), .C1(n5623), 
        .C2(n5429), .ZN(n844) );
  NAND2_X1 U2144 ( .A1(n5623), .A2(n826), .ZN(n827) );
  INV_X1 U2145 ( .A(n5856), .ZN(n826) );
  AOI221_X1 U2146 ( .B1(\UUT/Mpath/the_memhandle/N36 ), .B2(n992), .C1(
        \UUT/Mpath/the_memhandle/N38 ), .C2(n667), .A(n5872), .ZN(n991) );
  INV_X1 U2147 ( .A(n5869), .ZN(n667) );
  INV_X1 U2148 ( .A(n5870), .ZN(n992) );
  NAND2_X1 U2149 ( .A1(n5856), .A2(n5623), .ZN(n692) );
  AOI221_X1 U2150 ( .B1(n5664), .B2(D_DATA_INBUS[16]), .C1(n5663), .C2(
        D_DATA_INBUS[0]), .A(n5868), .ZN(n990) );
  OAI22_X1 U2151 ( .A1(n5429), .A2(\UUT/Mcontrol/N22 ), .B1(n989), .B2(n7395), 
        .ZN(n4163) );
  INV_X1 U2152 ( .A(n845), .ZN(n989) );
  OAI211_X1 U2153 ( .C1(n5526), .C2(n287), .A(n993), .B(n994), .ZN(n845) );
  AOI222_X1 U2154 ( .A1(\UUT/Mpath/the_mult/x_mult_out[0] ), .A2(n6357), .B1(
        n320), .B2(n995), .C1(n291), .C2(n996), .ZN(n994) );
  INV_X1 U2155 ( .A(n5622), .ZN(n996) );
  AOI22_X1 U2158 ( .A1(n6397), .A2(n999), .B1(n324), .B2(\UUT/daddr_out [0]), 
        .ZN(n993) );
  INV_X1 U2159 ( .A(n286), .ZN(n324) );
  INV_X1 U2160 ( .A(n5589), .ZN(n999) );
  OAI22_X1 U2161 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mpath/N111 ), .B1(n7226), 
        .B2(n1000), .ZN(n4164) );
  OAI221_X1 U2162 ( .B1(n5329), .B2(n1001), .C1(\UUT/Mpath/the_alu/N467 ), 
        .C2(\UUT/Mcontrol/N22 ), .A(n1002), .ZN(n4165) );
  NAND3_X1 U2163 ( .A1(n1003), .A2(\UUT/Mcontrol/N22 ), .A3(n1004), .ZN(n1002)
         );
  AOI21_X1 U2164 ( .B1(n7175), .B2(n1005), .A(n1007), .ZN(n1004) );
  INV_X1 U2165 ( .A(n7081), .ZN(n1007) );
  OAI22_X1 U2166 ( .A1(n1008), .A2(n556), .B1(n297), .B2(n2712), .ZN(n4166) );
  INV_X1 U2167 ( .A(\UUT/Mcontrol/Program_counter/N22 ), .ZN(n1008) );
  OAI22_X1 U2168 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mpath/the_memhandle/N236 ), .B1(n6287), .B2(n7396), .ZN(n4167) );
  OAI22_X1 U2169 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mpath/the_memhandle/N238 ), .B1(n1009), .B2(n7396), .ZN(n4168) );
  INV_X1 U2170 ( .A(dmem_ishalf), .ZN(n1009) );
  OAI22_X1 U2171 ( .A1(n5623), .A2(\UUT/Mcontrol/N22 ), .B1(n1010), .B2(n7396), 
        .ZN(n4169) );
  INV_X1 U2172 ( .A(dmem_read), .ZN(n1010) );
  OAI21_X1 U2173 ( .B1(\UUT/Mcontrol/N22 ), .B2(\UUT/Mpath/the_memhandle/N235 ), .A(n1011), .ZN(n4170) );
  OAI21_X1 U2174 ( .B1(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), .B2(
        \UUT/x_we ), .A(\UUT/Mcontrol/N22 ), .ZN(n1011) );
  OAI22_X1 U2175 ( .A1(n7386), .A2(n1012), .B1(n5315), .B2(\UUT/Mcontrol/N22 ), 
        .ZN(n4171) );
  OAI22_X1 U2176 ( .A1(n7386), .A2(\UUT/Mcontrol/N19 ), .B1(\UUT/Mcontrol/N22 ), .B2(n1012), .ZN(n4172) );
  OAI22_X1 U2177 ( .A1(n7386), .A2(n1014), .B1(\UUT/Mcontrol/N22 ), .B2(n2713), 
        .ZN(n4173) );
  OAI221_X1 U2178 ( .B1(n5775), .B2(n1015), .C1(\UUT/Mcontrol/N22 ), .C2(n1014), .A(n1016), .ZN(n4174) );
  AOI221_X1 U2179 ( .B1(n1017), .B2(\UUT/Mcontrol/d_sampled_finstr [12]), .C1(
        n1018), .C2(\UUT/Mcontrol/d_sampled_finstr [17]), .A(n1019), .ZN(n1016) );
  OAI22_X1 U2181 ( .A1(n7386), .A2(n1020), .B1(\UUT/Mcontrol/N22 ), .B2(n2715), 
        .ZN(n4175) );
  OAI221_X1 U2182 ( .B1(n5768), .B2(n1015), .C1(\UUT/Mcontrol/N22 ), .C2(n1020), .A(n1021), .ZN(n4176) );
  AOI221_X1 U2183 ( .B1(n1017), .B2(\UUT/Mcontrol/d_sampled_finstr [13]), .C1(
        n1018), .C2(\UUT/Mcontrol/d_sampled_finstr [18]), .A(n1019), .ZN(n1021) );
  OAI22_X1 U2185 ( .A1(n7386), .A2(n1022), .B1(\UUT/Mcontrol/N22 ), .B2(n2717), 
        .ZN(n4177) );
  OAI221_X1 U2186 ( .B1(n5760), .B2(n1015), .C1(\UUT/Mcontrol/N22 ), .C2(n1022), .A(n1023), .ZN(n4178) );
  AOI221_X1 U2187 ( .B1(n1017), .B2(\UUT/Mcontrol/d_sampled_finstr [14]), .C1(
        n1018), .C2(\UUT/Mcontrol/d_sampled_finstr [19]), .A(n1019), .ZN(n1023) );
  OAI22_X1 U2189 ( .A1(n7386), .A2(n1024), .B1(\UUT/Mcontrol/N22 ), .B2(n2719), 
        .ZN(n4179) );
  OAI221_X1 U2190 ( .B1(n5753), .B2(n1015), .C1(\UUT/Mcontrol/N22 ), .C2(n1024), .A(n1025), .ZN(n4180) );
  AOI221_X1 U2191 ( .B1(n1017), .B2(\UUT/Mcontrol/d_sampled_finstr [15]), .C1(
        n1018), .C2(\UUT/Mcontrol/d_sampled_finstr [20]), .A(n1019), .ZN(n1025) );
  NOR2_X1 U2193 ( .A1(n1026), .A2(n1027), .ZN(n4181) );
  AOI22_X1 U2194 ( .A1(\UUT/shift_op [0]), .A2(n7382), .B1(\UUT/Mcontrol/N22 ), 
        .B2(\UUT/Mcontrol/d_sampled_finstr [0]), .ZN(n1027) );
  OAI22_X1 U2195 ( .A1(n7386), .A2(n1028), .B1(\UUT/Mcontrol/N22 ), .B2(
        \UUT/Mpath/the_mult/N231 ), .ZN(n4182) );
  OAI22_X1 U2196 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1028), .B1(n1029), .B2(n7396), 
        .ZN(n4183) );
  INV_X1 U2197 ( .A(\UUT/Mpath/the_mult/x_mul_command[0] ), .ZN(n1028) );
  OAI22_X1 U2198 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mcontrol/st_logic/N34 ), 
        .B1(n1029), .B2(n7396), .ZN(n4184) );
  INV_X1 U2199 ( .A(\UUT/d_mul_command [0]), .ZN(n1029) );
  OAI21_X1 U2200 ( .B1(n5330), .B2(n297), .A(n1030), .ZN(n4185) );
  NAND2_X1 U2201 ( .A1(I_DATA_INBUS[0]), .A2(n297), .ZN(n1030) );
  NOR2_X1 U2202 ( .A1(n1026), .A2(n1031), .ZN(n4186) );
  AOI22_X1 U2203 ( .A1(\UUT/shift_op [1]), .A2(n7382), .B1(\UUT/Mcontrol/N22 ), 
        .B2(\UUT/Mcontrol/d_sampled_finstr [1]), .ZN(n1031) );
  OAI22_X1 U2204 ( .A1(n7387), .A2(n1032), .B1(\UUT/Mcontrol/N22 ), .B2(
        \UUT/Mpath/the_mult/N230 ), .ZN(n4187) );
  OAI22_X1 U2205 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1032), .B1(n1033), .B2(n7396), 
        .ZN(n4188) );
  OAI22_X1 U2207 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mcontrol/st_logic/N27 ), 
        .B1(n1033), .B2(n7397), .ZN(n4189) );
  INV_X1 U2208 ( .A(\UUT/d_mul_command [1]), .ZN(n1033) );
  OAI21_X1 U2209 ( .B1(n5329), .B2(n297), .A(n1034), .ZN(n4190) );
  NAND2_X1 U2210 ( .A1(I_DATA_INBUS[1]), .A2(n297), .ZN(n1034) );
  OAI221_X1 U2211 ( .B1(n7210), .B2(n1001), .C1(\UUT/Mcontrol/N22 ), .C2(n2724), .A(n1035), .ZN(n4191) );
  NOR2_X1 U2212 ( .A1(n1026), .A2(n1036), .ZN(n4192) );
  AOI22_X1 U2213 ( .A1(\UUT/shift_op [2]), .A2(n7382), .B1(\UUT/Mcontrol/N22 ), 
        .B2(\UUT/Mcontrol/d_sampled_finstr [2]), .ZN(n1036) );
  AND2_X1 U2214 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1037), .ZN(n1026) );
  OAI211_X1 U2215 ( .C1(n7100), .C2(n1038), .A(n7049), .B(n1039), .ZN(n1037)
         );
  OAI22_X1 U2216 ( .A1(n7387), .A2(n1040), .B1(\UUT/Mcontrol/N22 ), .B2(
        \UUT/Mpath/the_mult/N244 ), .ZN(n4193) );
  OAI22_X1 U2217 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1040), .B1(n1041), .B2(n7397), 
        .ZN(n4194) );
  OAI22_X1 U2219 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mcontrol/st_logic/N26 ), 
        .B1(n1041), .B2(n7397), .ZN(n4195) );
  INV_X1 U2220 ( .A(\UUT/d_mul_command [2]), .ZN(n1041) );
  OAI21_X1 U2221 ( .B1(n7210), .B2(n297), .A(n1042), .ZN(n4196) );
  NAND2_X1 U2222 ( .A1(I_DATA_INBUS[2]), .A2(n297), .ZN(n1042) );
  OAI221_X1 U2223 ( .B1(n5327), .B2(n1001), .C1(\UUT/Mcontrol/N22 ), .C2(n2727), .A(n1035), .ZN(n4197) );
  NAND3_X1 U2224 ( .A1(n1039), .A2(n1043), .A3(\UUT/Mcontrol/N22 ), .ZN(n1035)
         );
  OAI22_X1 U2225 ( .A1(n7387), .A2(n1044), .B1(\UUT/Mcontrol/N22 ), .B2(
        \UUT/Mpath/the_mult/N229 ), .ZN(n4198) );
  OAI22_X1 U2226 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1044), .B1(n1045), .B2(n7397), 
        .ZN(n4199) );
  INV_X1 U2227 ( .A(\UUT/Mpath/the_mult/x_mul_command[3] ), .ZN(n1044) );
  OAI22_X1 U2228 ( .A1(\UUT/Mcontrol/N22 ), .A2(n2728), .B1(n1045), .B2(n7397), 
        .ZN(n4200) );
  INV_X1 U2229 ( .A(\UUT/d_mul_command [3]), .ZN(n1045) );
  OAI21_X1 U2230 ( .B1(n5327), .B2(n297), .A(n1046), .ZN(n4201) );
  NAND2_X1 U2231 ( .A1(I_DATA_INBUS[3]), .A2(n297), .ZN(n1046) );
  OAI221_X1 U2232 ( .B1(n7221), .B2(n1001), .C1(\UUT/Mpath/the_alu/N453 ), 
        .C2(\UUT/Mcontrol/N22 ), .A(n1047), .ZN(n4202) );
  NAND4_X1 U2233 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1048), .A3(n1049), .A4(n5900), 
        .ZN(n1047) );
  NAND3_X1 U2234 ( .A1(n5944), .A2(n1050), .A3(n1051), .ZN(n1049) );
  OAI22_X1 U2235 ( .A1(n7387), .A2(n1052), .B1(\UUT/Mcontrol/N22 ), .B2(n2730), 
        .ZN(n4203) );
  OAI22_X1 U2236 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1052), .B1(n7391), .B2(n1053), 
        .ZN(n4204) );
  OAI22_X1 U2238 ( .A1(\UUT/Mcontrol/N22 ), .A2(n2732), .B1(n7391), .B2(n1053), 
        .ZN(n4205) );
  OAI21_X1 U2239 ( .B1(n7221), .B2(n297), .A(n1054), .ZN(n4206) );
  NAND2_X1 U2240 ( .A1(I_DATA_INBUS[4]), .A2(n297), .ZN(n1054) );
  OAI22_X1 U2241 ( .A1(\UUT/Mpath/the_alu/N466 ), .A2(\UUT/Mcontrol/N22 ), 
        .B1(n1055), .B2(n7397), .ZN(n4207) );
  AOI22_X1 U2242 ( .A1(n7098), .A2(n1057), .B1(
        \UUT/Mcontrol/d_sampled_finstr [5]), .B2(n1058), .ZN(n1055) );
  NAND2_X1 U2243 ( .A1(n1005), .A2(n1059), .ZN(n1057) );
  INV_X1 U2244 ( .A(n1043), .ZN(n1005) );
  OAI21_X1 U2245 ( .B1(n5946), .B2(n5944), .A(n1050), .ZN(n1043) );
  OAI22_X1 U2246 ( .A1(n7387), .A2(n1060), .B1(\UUT/Mcontrol/N22 ), .B2(n2734), 
        .ZN(n4208) );
  OAI22_X1 U2247 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1060), .B1(n7390), .B2(n1061), 
        .ZN(n4209) );
  OAI22_X1 U2249 ( .A1(\UUT/Mcontrol/N22 ), .A2(n2736), .B1(n7391), .B2(n1061), 
        .ZN(n4210) );
  OAI21_X1 U2250 ( .B1(n7203), .B2(n297), .A(n1062), .ZN(n4211) );
  NAND2_X1 U2251 ( .A1(I_DATA_INBUS[5]), .A2(n297), .ZN(n1062) );
  OAI21_X1 U2252 ( .B1(n6035), .B2(n297), .A(n1063), .ZN(n4212) );
  NAND2_X1 U2253 ( .A1(I_DATA_INBUS[6]), .A2(n297), .ZN(n1063) );
  OAI21_X1 U2254 ( .B1(n5971), .B2(n297), .A(n1064), .ZN(n4213) );
  NAND2_X1 U2255 ( .A1(I_DATA_INBUS[7]), .A2(n297), .ZN(n1064) );
  OAI21_X1 U2256 ( .B1(n5776), .B2(n297), .A(n1065), .ZN(n4214) );
  NAND2_X1 U2257 ( .A1(I_DATA_INBUS[8]), .A2(n297), .ZN(n1065) );
  OAI21_X1 U2258 ( .B1(n5769), .B2(n297), .A(n1066), .ZN(n4215) );
  NAND2_X1 U2259 ( .A1(I_DATA_INBUS[9]), .A2(n297), .ZN(n1066) );
  OAI21_X1 U2260 ( .B1(n5762), .B2(n297), .A(n1067), .ZN(n4216) );
  NAND2_X1 U2261 ( .A1(I_DATA_INBUS[10]), .A2(n297), .ZN(n1067) );
  OAI21_X1 U2262 ( .B1(n5906), .B2(n297), .A(n1068), .ZN(n4217) );
  NAND2_X1 U2263 ( .A1(I_DATA_INBUS[11]), .A2(n297), .ZN(n1068) );
  OAI21_X1 U2264 ( .B1(n5905), .B2(n297), .A(n1069), .ZN(n4218) );
  NAND2_X1 U2265 ( .A1(I_DATA_INBUS[12]), .A2(n297), .ZN(n1069) );
  OAI21_X1 U2266 ( .B1(n5903), .B2(n297), .A(n1070), .ZN(n4219) );
  NAND2_X1 U2267 ( .A1(I_DATA_INBUS[13]), .A2(n297), .ZN(n1070) );
  OAI21_X1 U2268 ( .B1(n5902), .B2(n297), .A(n1071), .ZN(n4220) );
  NAND2_X1 U2269 ( .A1(I_DATA_INBUS[14]), .A2(n297), .ZN(n1071) );
  OAI21_X1 U2270 ( .B1(n5720), .B2(n297), .A(n1072), .ZN(n4221) );
  NAND2_X1 U2271 ( .A1(I_DATA_INBUS[15]), .A2(n297), .ZN(n1072) );
  OAI21_X1 U2272 ( .B1(n5897), .B2(n297), .A(n1073), .ZN(n4222) );
  NAND2_X1 U2273 ( .A1(I_DATA_INBUS[16]), .A2(n297), .ZN(n1073) );
  OAI21_X1 U2274 ( .B1(n5904), .B2(n297), .A(n1074), .ZN(n4223) );
  NAND2_X1 U2275 ( .A1(I_DATA_INBUS[17]), .A2(n297), .ZN(n1074) );
  OAI21_X1 U2276 ( .B1(n5896), .B2(n297), .A(n1075), .ZN(n4224) );
  NAND2_X1 U2277 ( .A1(I_DATA_INBUS[18]), .A2(n297), .ZN(n1075) );
  OAI21_X1 U2278 ( .B1(n5901), .B2(n297), .A(n1076), .ZN(n4225) );
  NAND2_X1 U2279 ( .A1(I_DATA_INBUS[19]), .A2(n297), .ZN(n1076) );
  OAI21_X1 U2280 ( .B1(n5899), .B2(n297), .A(n1077), .ZN(n4226) );
  NAND2_X1 U2281 ( .A1(I_DATA_INBUS[20]), .A2(n297), .ZN(n1077) );
  OAI21_X1 U2282 ( .B1(n5907), .B2(n297), .A(n1078), .ZN(n4227) );
  NAND2_X1 U2283 ( .A1(I_DATA_INBUS[21]), .A2(n297), .ZN(n1078) );
  OAI21_X1 U2284 ( .B1(n5775), .B2(n297), .A(n1079), .ZN(n4228) );
  NAND2_X1 U2285 ( .A1(I_DATA_INBUS[22]), .A2(n297), .ZN(n1079) );
  OAI21_X1 U2286 ( .B1(n5768), .B2(n297), .A(n1080), .ZN(n4229) );
  NAND2_X1 U2287 ( .A1(I_DATA_INBUS[23]), .A2(n297), .ZN(n1080) );
  OAI21_X1 U2288 ( .B1(n5760), .B2(n297), .A(n1081), .ZN(n4230) );
  NAND2_X1 U2289 ( .A1(I_DATA_INBUS[24]), .A2(n297), .ZN(n1081) );
  OAI21_X1 U2290 ( .B1(n5753), .B2(n297), .A(n1082), .ZN(n4231) );
  NAND2_X1 U2291 ( .A1(I_DATA_INBUS[25]), .A2(n297), .ZN(n1082) );
  OAI21_X1 U2292 ( .B1(\UUT/Mcontrol/N22 ), .B2(n1083), .A(n1084), .ZN(n4232)
         );
  OAI21_X1 U2293 ( .B1(n1085), .B2(n1086), .A(\UUT/Mcontrol/N22 ), .ZN(n1084)
         );
  INV_X1 U2294 ( .A(n1087), .ZN(n1086) );
  NOR3_X1 U2295 ( .A1(n1088), .A2(n7041), .A3(n7075), .ZN(n1085) );
  OAI221_X1 U2296 ( .B1(n1089), .B2(n7398), .C1(\UUT/Mcontrol/N22 ), .C2(n1090), .A(n1091), .ZN(n4233) );
  AOI21_X1 U2297 ( .B1(n1092), .B2(n7101), .A(n6872), .ZN(n1089) );
  OAI21_X1 U2298 ( .B1(n7093), .B2(n1093), .A(n1094), .ZN(n1092) );
  NOR3_X1 U2299 ( .A1(n1088), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A3(n7075), .ZN(n1093) );
  INV_X1 U2300 ( .A(\UUT/Mcontrol/Operation_decoding32/N1987 ), .ZN(n1088) );
  OAI211_X1 U2301 ( .C1(\UUT/Mcontrol/N22 ), .C2(n1095), .A(n1096), .B(n1091), 
        .ZN(n4234) );
  NAND4_X1 U2302 ( .A1(n6988), .A2(\UUT/Mcontrol/N22 ), .A3(n7101), .A4(n6875), 
        .ZN(n1096) );
  OAI22_X1 U2303 ( .A1(\UUT/Mcontrol/N22 ), .A2(n2761), .B1(n1098), .B2(n7397), 
        .ZN(n4235) );
  OAI211_X1 U2304 ( .C1(\UUT/Mcontrol/N22 ), .C2(n1099), .A(n1100), .B(n1091), 
        .ZN(n4236) );
  NAND2_X1 U2305 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1101), .ZN(n1091) );
  OR3_X1 U2306 ( .A1(n1102), .A2(n1103), .A3(n7398), .ZN(n1100) );
  AOI21_X1 U2307 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2005 ), .B2(
        \UUT/Mcontrol/Operation_decoding32/N2017 ), .A(
        \UUT/Mcontrol/d_instr [26]), .ZN(n1102) );
  OAI22_X1 U2309 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1104), .B1(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .B2(n1000), .ZN(n4237) );
  INV_X1 U2310 ( .A(\UUT/exe_outsel [0]), .ZN(n1104) );
  OAI22_X1 U2311 ( .A1(\UUT/Mcontrol/N22 ), .A2(\UUT/Mpath/N116 ), .B1(n7191), 
        .B2(n1000), .ZN(n4238) );
  NAND2_X1 U2312 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1105), .ZN(n1000) );
  NAND4_X1 U2313 ( .A1(n7095), .A2(n7098), .A3(n1050), .A4(n1059), .ZN(n1105)
         );
  OAI21_X1 U2314 ( .B1(n297), .B2(n6997), .A(n1106), .ZN(n4239) );
  NAND2_X1 U2315 ( .A1(I_DATA_INBUS[26]), .A2(n297), .ZN(n1106) );
  OAI21_X1 U2316 ( .B1(n297), .B2(n2764), .A(n1107), .ZN(n4240) );
  NAND2_X1 U2317 ( .A1(I_DATA_INBUS[27]), .A2(n297), .ZN(n1107) );
  OAI21_X1 U2318 ( .B1(n297), .B2(n2765), .A(n1108), .ZN(n4241) );
  NAND2_X1 U2319 ( .A1(I_DATA_INBUS[28]), .A2(n297), .ZN(n1108) );
  OAI21_X1 U2320 ( .B1(\UUT/Mcontrol/Operation_decoding32/N1877 ), .B2(n297), 
        .A(n1109), .ZN(n4242) );
  NAND2_X1 U2321 ( .A1(I_DATA_INBUS[29]), .A2(n297), .ZN(n1109) );
  OAI21_X1 U2322 ( .B1(n7191), .B2(n297), .A(n1110), .ZN(n4243) );
  NAND2_X1 U2323 ( .A1(I_DATA_INBUS[30]), .A2(n297), .ZN(n1110) );
  OAI22_X1 U2324 ( .A1(n7388), .A2(n1111), .B1(\UUT/Mcontrol/N22 ), .B2(n1112), 
        .ZN(n4244) );
  OAI221_X1 U2326 ( .B1(n5907), .B2(n1015), .C1(\UUT/Mcontrol/N22 ), .C2(n1111), .A(n1113), .ZN(n4245) );
  AOI221_X1 U2327 ( .B1(n1017), .B2(\UUT/Mcontrol/d_sampled_finstr [11]), .C1(
        n1018), .C2(\UUT/Mcontrol/d_sampled_finstr [16]), .A(n1019), .ZN(n1113) );
  NOR4_X1 U2328 ( .A1(n1114), .A2(n5909), .A3(n5908), .A4(n7180), .ZN(n1019)
         );
  AND2_X1 U2329 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1115), .ZN(n1018) );
  OAI21_X1 U2330 ( .B1(n1116), .B2(n1117), .A(n1118), .ZN(n1115) );
  OAI21_X1 U2331 ( .B1(n1119), .B2(n1120), .A(n6868), .ZN(n1118) );
  NAND3_X1 U2333 ( .A1(n5911), .A2(n7101), .A3(n7145), .ZN(n1123) );
  NAND2_X1 U2334 ( .A1(n6879), .A2(n451), .ZN(n1121) );
  AOI21_X1 U2335 ( .B1(n1125), .B2(n6868), .A(n7397), .ZN(n1017) );
  OR3_X1 U2336 ( .A1(n1117), .A2(n1050), .A3(n7204), .ZN(n1125) );
  INV_X1 U2337 ( .A(n1003), .ZN(n1117) );
  NAND3_X1 U2339 ( .A1(n5914), .A2(n1126), .A3(n1127), .ZN(n1015) );
  NOR3_X1 U2340 ( .A1(n1128), .A2(n7117), .A3(n5937), .ZN(n1127) );
  INV_X1 U2341 ( .A(n1114), .ZN(n1126) );
  NAND3_X1 U2342 ( .A1(n1003), .A2(\UUT/Mcontrol/N22 ), .A3(n1122), .ZN(n1114)
         );
  NOR3_X1 U2343 ( .A1(n6872), .A2(n7179), .A3(n6827), .ZN(n1122) );
  NOR3_X1 U2344 ( .A1(n1119), .A2(n1058), .A3(n1120), .ZN(n1003) );
  INV_X1 U2345 ( .A(n5945), .ZN(n1120) );
  OAI21_X1 U2346 ( .B1(n7227), .B2(n297), .A(n1129), .ZN(n4246) );
  NAND2_X1 U2347 ( .A1(I_DATA_INBUS[31]), .A2(n297), .ZN(n1129) );
  OAI221_X1 U2351 ( .B1(n5330), .B2(n1001), .C1(\UUT/Mpath/the_alu/N468 ), 
        .C2(\UUT/Mcontrol/N22 ), .A(n1130), .ZN(n4247) );
  NAND3_X1 U2352 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1131), .A3(n1132), .ZN(n1130)
         );
  NAND3_X1 U2353 ( .A1(n1133), .A2(n7013), .A3(n1135), .ZN(n1131) );
  OAI21_X1 U2354 ( .B1(n7130), .B2(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
        .A(n1136), .ZN(n1135) );
  OAI21_X1 U2355 ( .B1(n7081), .B2(n7169), .A(n7127), .ZN(n1136) );
  NAND3_X1 U2356 ( .A1(n1137), .A2(\UUT/Mcontrol/Operation_decoding32/N2060 ), 
        .A3(n5947), .ZN(n1133) );
  INV_X1 U2357 ( .A(n1138), .ZN(n1137) );
  AOI21_X1 U2358 ( .B1(\UUT/Mcontrol/Operation_decoding32/N2047 ), .B2(n7130), 
        .A(\UUT/Mcontrol/Operation_decoding32/N1922 ), .ZN(n1138) );
  NAND2_X1 U2359 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1058), .ZN(n1001) );
  OAI22_X1 U2360 ( .A1(n7388), .A2(n1139), .B1(\UUT/Mcontrol/N22 ), .B2(n840), 
        .ZN(n4248) );
  INV_X1 U2362 ( .A(\UUT/Mpath/the_mult/x_mult_out[0] ), .ZN(n1139) );
  OAI22_X1 U2363 ( .A1(n7388), .A2(n1140), .B1(\UUT/Mcontrol/N22 ), .B2(n851), 
        .ZN(n4249) );
  INV_X1 U2365 ( .A(\UUT/Mpath/the_mult/x_mult_out[1] ), .ZN(n1140) );
  OAI22_X1 U2366 ( .A1(n7388), .A2(n1141), .B1(\UUT/Mcontrol/N22 ), .B2(n813), 
        .ZN(n4250) );
  INV_X1 U2368 ( .A(\UUT/Mpath/the_mult/x_mult_out[2] ), .ZN(n1141) );
  OAI22_X1 U2369 ( .A1(n7388), .A2(n1142), .B1(\UUT/Mcontrol/N22 ), .B2(n788), 
        .ZN(n4251) );
  INV_X1 U2371 ( .A(\UUT/Mpath/the_mult/x_mult_out[3] ), .ZN(n1142) );
  OAI22_X1 U2372 ( .A1(n7387), .A2(n1143), .B1(\UUT/Mcontrol/N22 ), .B2(n763), 
        .ZN(n4252) );
  INV_X1 U2374 ( .A(\UUT/Mpath/the_mult/x_mult_out[4] ), .ZN(n1143) );
  OAI22_X1 U2375 ( .A1(n7389), .A2(n1144), .B1(\UUT/Mcontrol/N22 ), .B2(n738), 
        .ZN(n4253) );
  INV_X1 U2377 ( .A(\UUT/Mpath/the_mult/x_mult_out[5] ), .ZN(n1144) );
  OAI22_X1 U2378 ( .A1(n7388), .A2(n1145), .B1(\UUT/Mcontrol/N22 ), .B2(n708), 
        .ZN(n4254) );
  INV_X1 U2380 ( .A(\UUT/Mpath/the_mult/x_mult_out[6] ), .ZN(n1145) );
  OAI22_X1 U2381 ( .A1(n7389), .A2(n1146), .B1(\UUT/Mcontrol/N22 ), .B2(n683), 
        .ZN(n4255) );
  INV_X1 U2383 ( .A(\UUT/Mpath/the_mult/x_mult_out[7] ), .ZN(n1146) );
  OAI22_X1 U2384 ( .A1(n7389), .A2(n1147), .B1(\UUT/Mcontrol/N22 ), .B2(n659), 
        .ZN(n4256) );
  INV_X1 U2386 ( .A(\UUT/Mpath/the_mult/x_mult_out[8] ), .ZN(n1147) );
  OAI22_X1 U2387 ( .A1(n7388), .A2(n1148), .B1(\UUT/Mcontrol/N22 ), .B2(n635), 
        .ZN(n4257) );
  INV_X1 U2389 ( .A(\UUT/Mpath/the_mult/x_mult_out[9] ), .ZN(n1148) );
  OAI22_X1 U2390 ( .A1(n7389), .A2(n1149), .B1(\UUT/Mcontrol/N22 ), .B2(n612), 
        .ZN(n4258) );
  INV_X1 U2392 ( .A(\UUT/Mpath/the_mult/x_mult_out[10] ), .ZN(n1149) );
  OAI22_X1 U2393 ( .A1(n7389), .A2(n1150), .B1(\UUT/Mcontrol/N22 ), .B2(n589), 
        .ZN(n4259) );
  INV_X1 U2395 ( .A(\UUT/Mpath/the_mult/x_mult_out[11] ), .ZN(n1150) );
  OAI22_X1 U2396 ( .A1(n7389), .A2(n1151), .B1(\UUT/Mcontrol/N22 ), .B2(n565), 
        .ZN(n4260) );
  INV_X1 U2398 ( .A(\UUT/Mpath/the_mult/x_mult_out[12] ), .ZN(n1151) );
  OAI22_X1 U2399 ( .A1(n7389), .A2(n1152), .B1(\UUT/Mcontrol/N22 ), .B2(n540), 
        .ZN(n4261) );
  INV_X1 U2401 ( .A(\UUT/Mpath/the_mult/x_mult_out[13] ), .ZN(n1152) );
  OAI22_X1 U2402 ( .A1(n7389), .A2(n1153), .B1(\UUT/Mcontrol/N22 ), .B2(n516), 
        .ZN(n4262) );
  INV_X1 U2404 ( .A(\UUT/Mpath/the_mult/x_mult_out[14] ), .ZN(n1153) );
  OAI22_X1 U2405 ( .A1(n7389), .A2(n1154), .B1(\UUT/Mcontrol/N22 ), .B2(n489), 
        .ZN(n4263) );
  INV_X1 U2407 ( .A(\UUT/Mpath/the_mult/x_mult_out[15] ), .ZN(n1154) );
  OAI22_X1 U2408 ( .A1(n7390), .A2(n1155), .B1(\UUT/Mcontrol/N22 ), .B2(n461), 
        .ZN(n4264) );
  INV_X1 U2410 ( .A(\UUT/Mpath/the_mult/x_mult_out[16] ), .ZN(n1155) );
  OAI22_X1 U2411 ( .A1(n7389), .A2(n1156), .B1(\UUT/Mcontrol/N22 ), .B2(n432), 
        .ZN(n4265) );
  INV_X1 U2413 ( .A(\UUT/Mpath/the_mult/x_mult_out[17] ), .ZN(n1156) );
  OAI22_X1 U2414 ( .A1(n7389), .A2(n1157), .B1(\UUT/Mcontrol/N22 ), .B2(n408), 
        .ZN(n4266) );
  INV_X1 U2416 ( .A(\UUT/Mpath/the_mult/x_mult_out[18] ), .ZN(n1157) );
  OAI22_X1 U2417 ( .A1(n7390), .A2(n1158), .B1(\UUT/Mcontrol/N22 ), .B2(n384), 
        .ZN(n4267) );
  INV_X1 U2419 ( .A(\UUT/Mpath/the_mult/x_mult_out[19] ), .ZN(n1158) );
  OAI22_X1 U2420 ( .A1(n7390), .A2(n1159), .B1(\UUT/Mcontrol/N22 ), .B2(n357), 
        .ZN(n4268) );
  INV_X1 U2422 ( .A(\UUT/Mpath/the_mult/x_mult_out[20] ), .ZN(n1159) );
  OAI22_X1 U2423 ( .A1(n7390), .A2(n1160), .B1(\UUT/Mcontrol/N22 ), .B2(n334), 
        .ZN(n4269) );
  INV_X1 U2425 ( .A(\UUT/Mpath/the_mult/x_mult_out[21] ), .ZN(n1160) );
  OAI22_X1 U2426 ( .A1(n7390), .A2(n1161), .B1(\UUT/Mcontrol/N22 ), .B2(n309), 
        .ZN(n4270) );
  INV_X1 U2428 ( .A(\UUT/Mpath/the_mult/x_mult_out[22] ), .ZN(n1161) );
  OAI22_X1 U2429 ( .A1(n7389), .A2(n1162), .B1(\UUT/Mcontrol/N22 ), .B2(n863), 
        .ZN(n4271) );
  INV_X1 U2431 ( .A(\UUT/Mpath/the_mult/x_mult_out[23] ), .ZN(n1162) );
  OAI22_X1 U2432 ( .A1(n7390), .A2(n1163), .B1(\UUT/Mcontrol/N22 ), .B2(n212), 
        .ZN(n4272) );
  INV_X1 U2434 ( .A(\UUT/Mpath/the_mult/x_mult_out[24] ), .ZN(n1163) );
  OAI22_X1 U2435 ( .A1(n7390), .A2(n1164), .B1(\UUT/Mcontrol/N22 ), .B2(n189), 
        .ZN(n4273) );
  INV_X1 U2437 ( .A(\UUT/Mpath/the_mult/x_mult_out[25] ), .ZN(n1164) );
  OAI22_X1 U2438 ( .A1(n7390), .A2(n1165), .B1(\UUT/Mcontrol/N22 ), .B2(n173), 
        .ZN(n4274) );
  INV_X1 U2440 ( .A(\UUT/Mpath/the_mult/x_mult_out[26] ), .ZN(n1165) );
  OAI22_X1 U2441 ( .A1(n7390), .A2(n1166), .B1(\UUT/Mcontrol/N22 ), .B2(n156), 
        .ZN(n4275) );
  INV_X1 U2443 ( .A(\UUT/Mpath/the_mult/x_mult_out[27] ), .ZN(n1166) );
  OAI22_X1 U2444 ( .A1(n7390), .A2(n1167), .B1(\UUT/Mcontrol/N22 ), .B2(n139), 
        .ZN(n4276) );
  INV_X1 U2446 ( .A(\UUT/Mpath/the_mult/x_mult_out[28] ), .ZN(n1167) );
  OAI22_X1 U2447 ( .A1(n7390), .A2(n1168), .B1(\UUT/Mcontrol/N22 ), .B2(n116), 
        .ZN(n4277) );
  INV_X1 U2449 ( .A(\UUT/Mpath/the_mult/x_mult_out[29] ), .ZN(n1168) );
  OAI22_X1 U2450 ( .A1(n7388), .A2(n1169), .B1(\UUT/Mcontrol/N22 ), .B2(n921), 
        .ZN(n4278) );
  INV_X1 U2452 ( .A(n6835), .ZN(n1169) );
  OAI22_X1 U2453 ( .A1(n7382), .A2(n1170), .B1(\UUT/Mcontrol/N22 ), .B2(n873), 
        .ZN(n4279) );
  INV_X1 U2455 ( .A(n7155), .ZN(n1170) );
  INV_X1 U2456 ( .A(\UUT/Mcontrol/N22 ), .ZN(n122) );
  OAI21_X1 U2457 ( .B1(\UUT/Mcontrol/N22 ), .B2(n837), .A(n1171), .ZN(n4280)
         );
  NAND2_X1 U2458 ( .A1(\UUT/Mpath/the_mult/x_mult_out[32] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1171) );
  OAI21_X1 U2460 ( .B1(\UUT/Mcontrol/N22 ), .B2(n848), .A(n1172), .ZN(n4281)
         );
  NAND2_X1 U2461 ( .A1(\UUT/Mpath/the_mult/x_mult_out[33] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1172) );
  OAI21_X1 U2463 ( .B1(\UUT/Mcontrol/N22 ), .B2(n810), .A(n1173), .ZN(n4282)
         );
  NAND2_X1 U2464 ( .A1(\UUT/Mpath/the_mult/x_mult_out[34] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1173) );
  INV_X1 U2465 ( .A(\UUT/Mpath/the_mult/Mult_out[34] ), .ZN(n810) );
  OAI21_X1 U2466 ( .B1(\UUT/Mcontrol/N22 ), .B2(n785), .A(n1174), .ZN(n4283)
         );
  NAND2_X1 U2467 ( .A1(\UUT/Mpath/the_mult/x_mult_out[35] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1174) );
  INV_X1 U2468 ( .A(\UUT/Mpath/the_mult/Mult_out[35] ), .ZN(n785) );
  OAI21_X1 U2469 ( .B1(\UUT/Mcontrol/N22 ), .B2(n760), .A(n1175), .ZN(n4284)
         );
  NAND2_X1 U2470 ( .A1(\UUT/Mpath/the_mult/x_mult_out[36] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1175) );
  INV_X1 U2471 ( .A(\UUT/Mpath/the_mult/Mult_out[36] ), .ZN(n760) );
  OAI21_X1 U2472 ( .B1(\UUT/Mcontrol/N22 ), .B2(n735), .A(n1176), .ZN(n4285)
         );
  NAND2_X1 U2473 ( .A1(\UUT/Mpath/the_mult/x_mult_out[37] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1176) );
  INV_X1 U2474 ( .A(\UUT/Mpath/the_mult/Mult_out[37] ), .ZN(n735) );
  OAI21_X1 U2475 ( .B1(\UUT/Mcontrol/N22 ), .B2(n705), .A(n1177), .ZN(n4286)
         );
  NAND2_X1 U2476 ( .A1(\UUT/Mpath/the_mult/x_mult_out[38] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1177) );
  INV_X1 U2477 ( .A(\UUT/Mpath/the_mult/Mult_out[38] ), .ZN(n705) );
  OAI21_X1 U2478 ( .B1(\UUT/Mcontrol/N22 ), .B2(n680), .A(n1178), .ZN(n4287)
         );
  NAND2_X1 U2479 ( .A1(\UUT/Mpath/the_mult/x_mult_out[39] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1178) );
  INV_X1 U2480 ( .A(\UUT/Mpath/the_mult/Mult_out[39] ), .ZN(n680) );
  OAI21_X1 U2481 ( .B1(\UUT/Mcontrol/N22 ), .B2(n656), .A(n1179), .ZN(n4288)
         );
  NAND2_X1 U2482 ( .A1(\UUT/Mpath/the_mult/x_mult_out[40] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1179) );
  INV_X1 U2483 ( .A(\UUT/Mpath/the_mult/Mult_out[40] ), .ZN(n656) );
  OAI21_X1 U2484 ( .B1(\UUT/Mcontrol/N22 ), .B2(n632), .A(n1180), .ZN(n4289)
         );
  NAND2_X1 U2485 ( .A1(\UUT/Mpath/the_mult/x_mult_out[41] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1180) );
  INV_X1 U2486 ( .A(\UUT/Mpath/the_mult/Mult_out[41] ), .ZN(n632) );
  OAI21_X1 U2487 ( .B1(\UUT/Mcontrol/N22 ), .B2(n609), .A(n1181), .ZN(n4290)
         );
  NAND2_X1 U2488 ( .A1(\UUT/Mpath/the_mult/x_mult_out[42] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1181) );
  INV_X1 U2489 ( .A(\UUT/Mpath/the_mult/Mult_out[42] ), .ZN(n609) );
  OAI21_X1 U2490 ( .B1(\UUT/Mcontrol/N22 ), .B2(n586), .A(n1182), .ZN(n4291)
         );
  NAND2_X1 U2491 ( .A1(\UUT/Mpath/the_mult/x_mult_out[43] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1182) );
  INV_X1 U2492 ( .A(\UUT/Mpath/the_mult/Mult_out[43] ), .ZN(n586) );
  OAI21_X1 U2493 ( .B1(\UUT/Mcontrol/N22 ), .B2(n562), .A(n1183), .ZN(n4292)
         );
  NAND2_X1 U2494 ( .A1(\UUT/Mpath/the_mult/x_mult_out[44] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1183) );
  INV_X1 U2495 ( .A(\UUT/Mpath/the_mult/Mult_out[44] ), .ZN(n562) );
  OAI21_X1 U2496 ( .B1(\UUT/Mcontrol/N22 ), .B2(n537), .A(n1184), .ZN(n4293)
         );
  NAND2_X1 U2497 ( .A1(\UUT/Mpath/the_mult/x_mult_out[45] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1184) );
  INV_X1 U2498 ( .A(\UUT/Mpath/the_mult/Mult_out[45] ), .ZN(n537) );
  OAI21_X1 U2499 ( .B1(\UUT/Mcontrol/N22 ), .B2(n513), .A(n1185), .ZN(n4294)
         );
  NAND2_X1 U2500 ( .A1(\UUT/Mpath/the_mult/x_mult_out[46] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1185) );
  INV_X1 U2501 ( .A(\UUT/Mpath/the_mult/Mult_out[46] ), .ZN(n513) );
  OAI21_X1 U2502 ( .B1(\UUT/Mcontrol/N22 ), .B2(n486), .A(n1186), .ZN(n4295)
         );
  NAND2_X1 U2503 ( .A1(\UUT/Mpath/the_mult/x_mult_out[47] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1186) );
  INV_X1 U2504 ( .A(\UUT/Mpath/the_mult/Mult_out[47] ), .ZN(n486) );
  OAI21_X1 U2505 ( .B1(\UUT/Mcontrol/N22 ), .B2(n458), .A(n1187), .ZN(n4296)
         );
  NAND2_X1 U2506 ( .A1(\UUT/Mpath/the_mult/x_mult_out[48] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1187) );
  INV_X1 U2507 ( .A(\UUT/Mpath/the_mult/Mult_out[48] ), .ZN(n458) );
  OAI21_X1 U2508 ( .B1(\UUT/Mcontrol/N22 ), .B2(n429), .A(n1188), .ZN(n4297)
         );
  NAND2_X1 U2509 ( .A1(\UUT/Mpath/the_mult/x_mult_out[49] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1188) );
  INV_X1 U2510 ( .A(\UUT/Mpath/the_mult/Mult_out[49] ), .ZN(n429) );
  OAI21_X1 U2511 ( .B1(\UUT/Mcontrol/N22 ), .B2(n405), .A(n1189), .ZN(n4298)
         );
  NAND2_X1 U2512 ( .A1(\UUT/Mpath/the_mult/x_mult_out[50] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1189) );
  INV_X1 U2513 ( .A(\UUT/Mpath/the_mult/Mult_out[50] ), .ZN(n405) );
  OAI21_X1 U2514 ( .B1(\UUT/Mcontrol/N22 ), .B2(n381), .A(n1190), .ZN(n4299)
         );
  NAND2_X1 U2515 ( .A1(\UUT/Mpath/the_mult/x_mult_out[51] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1190) );
  INV_X1 U2516 ( .A(\UUT/Mpath/the_mult/Mult_out[51] ), .ZN(n381) );
  OAI21_X1 U2517 ( .B1(\UUT/Mcontrol/N22 ), .B2(n354), .A(n1191), .ZN(n4300)
         );
  NAND2_X1 U2518 ( .A1(\UUT/Mpath/the_mult/x_mult_out[52] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1191) );
  INV_X1 U2519 ( .A(\UUT/Mpath/the_mult/Mult_out[52] ), .ZN(n354) );
  OAI21_X1 U2520 ( .B1(\UUT/Mcontrol/N22 ), .B2(n331), .A(n1192), .ZN(n4301)
         );
  NAND2_X1 U2521 ( .A1(\UUT/Mpath/the_mult/x_mult_out[53] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1192) );
  INV_X1 U2522 ( .A(\UUT/Mpath/the_mult/Mult_out[53] ), .ZN(n331) );
  OAI21_X1 U2523 ( .B1(\UUT/Mcontrol/N22 ), .B2(n306), .A(n1193), .ZN(n4302)
         );
  NAND2_X1 U2524 ( .A1(\UUT/Mpath/the_mult/x_mult_out[54] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1193) );
  INV_X1 U2525 ( .A(\UUT/Mpath/the_mult/Mult_out[54] ), .ZN(n306) );
  OAI21_X1 U2526 ( .B1(\UUT/Mcontrol/N22 ), .B2(n860), .A(n1194), .ZN(n4303)
         );
  NAND2_X1 U2527 ( .A1(\UUT/Mpath/the_mult/x_mult_out[55] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1194) );
  INV_X1 U2528 ( .A(\UUT/Mpath/the_mult/Mult_out[55] ), .ZN(n860) );
  OAI21_X1 U2529 ( .B1(\UUT/Mcontrol/N22 ), .B2(n209), .A(n1195), .ZN(n4304)
         );
  NAND2_X1 U2530 ( .A1(\UUT/Mpath/the_mult/x_mult_out[56] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1195) );
  INV_X1 U2531 ( .A(\UUT/Mpath/the_mult/Mult_out[56] ), .ZN(n209) );
  OAI21_X1 U2532 ( .B1(\UUT/Mcontrol/N22 ), .B2(n186), .A(n1196), .ZN(n4305)
         );
  NAND2_X1 U2533 ( .A1(\UUT/Mpath/the_mult/x_mult_out[57] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1196) );
  INV_X1 U2534 ( .A(\UUT/Mpath/the_mult/Mult_out[57] ), .ZN(n186) );
  OAI21_X1 U2535 ( .B1(\UUT/Mcontrol/N22 ), .B2(n170), .A(n1197), .ZN(n4306)
         );
  NAND2_X1 U2536 ( .A1(\UUT/Mpath/the_mult/x_mult_out[58] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1197) );
  INV_X1 U2537 ( .A(\UUT/Mpath/the_mult/Mult_out[58] ), .ZN(n170) );
  OAI21_X1 U2538 ( .B1(\UUT/Mcontrol/N22 ), .B2(n153), .A(n1198), .ZN(n4307)
         );
  NAND2_X1 U2539 ( .A1(\UUT/Mpath/the_mult/x_mult_out[59] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1198) );
  INV_X1 U2540 ( .A(\UUT/Mpath/the_mult/Mult_out[59] ), .ZN(n153) );
  OAI21_X1 U2541 ( .B1(\UUT/Mcontrol/N22 ), .B2(n136), .A(n1199), .ZN(n4308)
         );
  NAND2_X1 U2542 ( .A1(\UUT/Mpath/the_mult/x_mult_out[60] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1199) );
  INV_X1 U2543 ( .A(\UUT/Mpath/the_mult/Mult_out[60] ), .ZN(n136) );
  OAI21_X1 U2544 ( .B1(\UUT/Mcontrol/N22 ), .B2(n919), .A(n1200), .ZN(n4309)
         );
  NAND2_X1 U2545 ( .A1(\UUT/Mpath/the_mult/x_mult_out[61] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1200) );
  INV_X1 U2546 ( .A(\UUT/Mpath/the_mult/Mult_out[61] ), .ZN(n919) );
  NAND2_X1 U2548 ( .A1(\UUT/Mpath/the_mult/x_mult_out[62] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1201) );
  INV_X1 U2549 ( .A(\UUT/Mpath/the_mult/Mult_out[62] ), .ZN(n930) );
  OAI21_X1 U2550 ( .B1(\UUT/Mcontrol/N22 ), .B2(n104), .A(n1202), .ZN(n4311)
         );
  NAND2_X1 U2551 ( .A1(\UUT/Mpath/the_mult/x_mult_out[63] ), .A2(
        \UUT/Mcontrol/N22 ), .ZN(n1202) );
  INV_X1 U2552 ( .A(\UUT/Mpath/the_mult/Mult_out[63] ), .ZN(n104) );
  OAI22_X1 U2553 ( .A1(n46), .A2(n2835), .B1(n48), .B2(n86), .ZN(n4312) );
  OAI222_X1 U2555 ( .A1(n880), .A2(n101), .B1(n948), .B2(n99), .C1(n5356), 
        .C2(n102), .ZN(n1203) );
  NOR3_X1 U2561 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n293) );
  INV_X1 U2562 ( .A(\UUT/Mpath/the_mult/N198 ), .ZN(n1207) );
  INV_X1 U2563 ( .A(n5598), .ZN(n1206) );
  INV_X1 U2565 ( .A(n5541), .ZN(n1205) );
  NOR3_X1 U2566 ( .A1(n1208), .A2(\UUT/Mpath/the_mult/N198 ), .A3(n1209), .ZN(
        n289) );
  INV_X1 U2567 ( .A(\UUT/Mpath/the_mult/N216 ), .ZN(n1209) );
  NAND2_X1 U2568 ( .A1(n287), .A2(n998), .ZN(n1208) );
  INV_X1 U2569 ( .A(\UUT/Mpath/N125 ), .ZN(n998) );
  NAND3_X1 U2570 ( .A1(\UUT/Mpath/N125 ), .A2(n287), .A3(\UUT/Mpath/N128 ), 
        .ZN(n286) );
  NOR2_X1 U2572 ( .A1(\UUT/exe_outsel [0]), .A2(\UUT/Mpath/N121 ), .ZN(n997)
         );
  OAI221_X1 U2575 ( .B1(n5668), .B2(n284), .C1(n5623), .C2(n5357), .A(n285), 
        .ZN(n877) );
  INV_X1 U2577 ( .A(n693), .ZN(n499) );
  NAND2_X1 U2578 ( .A1(n5626), .A2(n5623), .ZN(n693) );
  NOR4_X1 U2579 ( .A1(n5822), .A2(n5823), .A3(n825), .A4(n1211), .ZN(n1210) );
  INV_X1 U2580 ( .A(\UUT/Mpath/the_memhandle/N86 ), .ZN(n1211) );
  OR3_X1 U2581 ( .A1(n5823), .A2(n5825), .A3(n825), .ZN(n284) );
  INV_X1 U2582 ( .A(n5623), .ZN(n825) );
  AND4_X1 U2585 ( .A1(n1087), .A2(n1212), .A3(n6875), .A4(n1094), .ZN(n1098)
         );
  INV_X1 U2586 ( .A(n7012), .ZN(n1094) );
  NAND3_X1 U2587 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1981 ), .A2(n7021), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N1987 ), .ZN(n1212) );
  NOR4_X1 U2588 ( .A1(n1101), .A2(n6872), .A3(n1103), .A4(n7093), .ZN(n1087)
         );
  INV_X1 U2589 ( .A(n5920), .ZN(n1101) );
  INV_X1 U2590 ( .A(dmem_isbyte), .ZN(n6287) );
  NAND3_X1 U2591 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n6130) );
  AOI222_X1 U2592 ( .A1(\UUT/Mpath/the_alu/sum[10] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N147 ), .B2(n6834), .C1(n1218), .C2(n1219), .ZN(
        n1215) );
  AOI22_X1 U2594 ( .A1(\UUT/Mpath/the_alu/N211 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N179 ), .B2(n1221), .ZN(n1214) );
  AOI22_X1 U2595 ( .A1(\UUT/Mpath/the_alu/N115 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[10] ), .B2(n1223), .ZN(n1213) );
  AND2_X1 U2596 ( .A1(n1224), .A2(n1225), .ZN(n6129) );
  AOI222_X1 U2597 ( .A1(\UUT/Mpath/the_shift/sh_rol [10]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [10]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [10]), .C2(n1228), .ZN(n1225) );
  AOI22_X1 U2598 ( .A1(\UUT/Mpath/the_shift/sh_sra [10]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [10]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1224) );
  NAND3_X1 U2599 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n6128) );
  AOI222_X1 U2600 ( .A1(\UUT/Mpath/the_alu/sum[11] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N146 ), .B2(n6834), .C1(n1218), .C2(n1233), .ZN(
        n1232) );
  INV_X1 U2601 ( .A(\UUT/Mpath/the_alu/N61 ), .ZN(n1233) );
  AOI22_X1 U2602 ( .A1(\UUT/Mpath/the_alu/N210 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N178 ), .B2(n1221), .ZN(n1231) );
  AOI22_X1 U2603 ( .A1(\UUT/Mpath/the_alu/N114 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[11] ), .B2(n1223), .ZN(n1230) );
  AND2_X1 U2604 ( .A1(n1234), .A2(n1235), .ZN(n6127) );
  AOI222_X1 U2605 ( .A1(\UUT/Mpath/the_shift/sh_rol [11]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [11]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [11]), .C2(n1228), .ZN(n1235) );
  AOI22_X1 U2606 ( .A1(\UUT/Mpath/the_shift/sh_sra [11]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [11]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1234) );
  NAND3_X1 U2607 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n6126) );
  AOI222_X1 U2608 ( .A1(\UUT/Mpath/the_alu/sum[12] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N145 ), .B2(n6834), .C1(n1218), .C2(n1239), .ZN(
        n1238) );
  INV_X1 U2609 ( .A(\UUT/Mpath/the_alu/N59 ), .ZN(n1239) );
  AOI22_X1 U2610 ( .A1(\UUT/Mpath/the_alu/N209 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N177 ), .B2(n1221), .ZN(n1237) );
  AOI22_X1 U2611 ( .A1(\UUT/Mpath/the_alu/N113 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[12] ), .B2(n1223), .ZN(n1236) );
  AND2_X1 U2612 ( .A1(n1240), .A2(n1241), .ZN(n6125) );
  AOI222_X1 U2613 ( .A1(\UUT/Mpath/the_shift/sh_rol [12]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [12]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [12]), .C2(n1228), .ZN(n1241) );
  AOI22_X1 U2614 ( .A1(\UUT/Mpath/the_shift/sh_sra [12]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [12]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1240) );
  NAND3_X1 U2615 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n6124) );
  AOI222_X1 U2616 ( .A1(\UUT/Mpath/the_alu/sum[13] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N144 ), .B2(n6834), .C1(n1218), .C2(n1245), .ZN(
        n1244) );
  AOI22_X1 U2618 ( .A1(\UUT/Mpath/the_alu/N208 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N176 ), .B2(n1221), .ZN(n1243) );
  AOI22_X1 U2619 ( .A1(\UUT/Mpath/the_alu/N112 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[13] ), .B2(n1223), .ZN(n1242) );
  NAND3_X1 U2620 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n6123) );
  AOI222_X1 U2621 ( .A1(\UUT/Mpath/the_alu/sum[14] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N143 ), .B2(n6834), .C1(n1218), .C2(n1249), .ZN(
        n1248) );
  INV_X1 U2622 ( .A(\UUT/Mpath/the_alu/N55 ), .ZN(n1249) );
  AOI22_X1 U2623 ( .A1(\UUT/Mpath/the_alu/N207 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N175 ), .B2(n1221), .ZN(n1247) );
  AOI22_X1 U2624 ( .A1(\UUT/Mpath/the_alu/N111 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[14] ), .B2(n1223), .ZN(n1246) );
  NAND3_X1 U2625 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n6122) );
  AOI222_X1 U2626 ( .A1(\UUT/Mpath/the_alu/sum[15] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N142 ), .B2(n6834), .C1(n1218), .C2(n1253), .ZN(
        n1252) );
  INV_X1 U2627 ( .A(\UUT/Mpath/the_alu/N53 ), .ZN(n1253) );
  AOI22_X1 U2628 ( .A1(\UUT/Mpath/the_alu/N206 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N174 ), .B2(n1221), .ZN(n1251) );
  AOI22_X1 U2629 ( .A1(\UUT/Mpath/the_alu/N110 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[15] ), .B2(n1223), .ZN(n1250) );
  NAND3_X1 U2630 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n6121) );
  AOI222_X1 U2631 ( .A1(\UUT/Mpath/the_alu/sum[16] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N141 ), .B2(n6834), .C1(n1218), .C2(n1257), .ZN(
        n1256) );
  INV_X1 U2632 ( .A(\UUT/Mpath/the_alu/N51 ), .ZN(n1257) );
  AOI22_X1 U2633 ( .A1(\UUT/Mpath/the_alu/N205 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N173 ), .B2(n1221), .ZN(n1255) );
  AOI22_X1 U2634 ( .A1(\UUT/Mpath/the_alu/N109 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[16] ), .B2(n1223), .ZN(n1254) );
  NAND3_X1 U2635 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n6120) );
  AOI222_X1 U2636 ( .A1(\UUT/Mpath/the_alu/sum[17] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N140 ), .B2(n6834), .C1(n1218), .C2(n1261), .ZN(
        n1260) );
  AOI22_X1 U2638 ( .A1(\UUT/Mpath/the_alu/N204 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N172 ), .B2(n1221), .ZN(n1259) );
  AOI22_X1 U2639 ( .A1(\UUT/Mpath/the_alu/N108 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[17] ), .B2(n1223), .ZN(n1258) );
  NAND3_X1 U2640 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n6119) );
  AOI222_X1 U2641 ( .A1(\UUT/Mpath/the_alu/sum[18] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N139 ), .B2(n6834), .C1(n1218), .C2(n1265), .ZN(
        n1264) );
  AOI22_X1 U2643 ( .A1(\UUT/Mpath/the_alu/N203 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N171 ), .B2(n1221), .ZN(n1263) );
  AOI22_X1 U2644 ( .A1(\UUT/Mpath/the_alu/N107 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[18] ), .B2(n1223), .ZN(n1262) );
  NAND3_X1 U2645 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n6118) );
  AOI222_X1 U2646 ( .A1(\UUT/Mpath/the_alu/sum[19] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N138 ), .B2(n6834), .C1(n1218), .C2(n1269), .ZN(
        n1268) );
  INV_X1 U2647 ( .A(\UUT/Mpath/the_alu/N45 ), .ZN(n1269) );
  AOI22_X1 U2648 ( .A1(\UUT/Mpath/the_alu/N202 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N170 ), .B2(n1221), .ZN(n1267) );
  AOI22_X1 U2649 ( .A1(\UUT/Mpath/the_alu/N106 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[19] ), .B2(n1223), .ZN(n1266) );
  NAND3_X1 U2650 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n6117) );
  INV_X1 U2652 ( .A(\UUT/Mpath/the_alu/N43 ), .ZN(n1273) );
  AOI22_X1 U2653 ( .A1(\UUT/Mpath/the_alu/N201 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N169 ), .B2(n1221), .ZN(n1271) );
  AOI22_X1 U2654 ( .A1(\UUT/Mpath/the_alu/N105 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[20] ), .B2(n1223), .ZN(n1270) );
  NAND3_X1 U2655 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n6116) );
  AOI222_X1 U2656 ( .A1(\UUT/Mpath/the_alu/sum[21] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N136 ), .B2(n6834), .C1(n1218), .C2(n1277), .ZN(
        n1276) );
  INV_X1 U2657 ( .A(\UUT/Mpath/the_alu/N41 ), .ZN(n1277) );
  AOI22_X1 U2658 ( .A1(\UUT/Mpath/the_alu/N200 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N168 ), .B2(n1221), .ZN(n1275) );
  AOI22_X1 U2659 ( .A1(\UUT/Mpath/the_alu/N104 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[21] ), .B2(n1223), .ZN(n1274) );
  NAND3_X1 U2660 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n6115) );
  AOI222_X1 U2661 ( .A1(\UUT/Mpath/the_alu/sum[22] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N135 ), .B2(n6834), .C1(n1218), .C2(n1281), .ZN(
        n1280) );
  INV_X1 U2662 ( .A(\UUT/Mpath/the_alu/N39 ), .ZN(n1281) );
  AOI22_X1 U2663 ( .A1(\UUT/Mpath/the_alu/N199 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N167 ), .B2(n1221), .ZN(n1279) );
  AOI22_X1 U2664 ( .A1(\UUT/Mpath/the_alu/N103 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[22] ), .B2(n1223), .ZN(n1278) );
  NAND3_X1 U2665 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n6114) );
  AOI222_X1 U2666 ( .A1(\UUT/Mpath/the_alu/sum[23] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N134 ), .B2(n6834), .C1(n1218), .C2(n1285), .ZN(
        n1284) );
  INV_X1 U2667 ( .A(\UUT/Mpath/the_alu/N37 ), .ZN(n1285) );
  AOI22_X1 U2668 ( .A1(\UUT/Mpath/the_alu/N198 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N166 ), .B2(n1221), .ZN(n1283) );
  AOI22_X1 U2669 ( .A1(\UUT/Mpath/the_alu/N102 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[23] ), .B2(n1223), .ZN(n1282) );
  NAND3_X1 U2670 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n6113) );
  AOI222_X1 U2671 ( .A1(\UUT/Mpath/the_alu/sum[2] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N155 ), .B2(n6834), .C1(n1218), .C2(n1289), .ZN(
        n1288) );
  INV_X1 U2672 ( .A(\UUT/Mpath/the_alu/N79 ), .ZN(n1289) );
  AOI22_X1 U2673 ( .A1(\UUT/Mpath/the_alu/N219 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N187 ), .B2(n1221), .ZN(n1287) );
  AOI22_X1 U2674 ( .A1(\UUT/Mpath/the_alu/N123 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[2] ), .B2(n1223), .ZN(n1286) );
  AND2_X1 U2675 ( .A1(n1290), .A2(n1291), .ZN(n6112) );
  AOI222_X1 U2676 ( .A1(\UUT/Mpath/the_shift/sh_rol [2]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [2]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [2]), .C2(n1228), .ZN(n1291) );
  AOI22_X1 U2677 ( .A1(\UUT/Mpath/the_shift/sh_sra [2]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [2]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1290) );
  AOI22_X1 U2680 ( .A1(\UUT/Mpath/the_shift/sh_sra [31]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [31]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1292) );
  INV_X1 U2681 ( .A(n1294), .ZN(n6110) );
  OAI211_X1 U2682 ( .C1(\UUT/Mpath/the_alu/N21 ), .C2(n7215), .A(n1296), .B(
        n1297), .ZN(n1294) );
  AOI22_X1 U2683 ( .A1(\UUT/Mpath/the_alu/diff[31] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[31] ), .B2(n7213), .ZN(n1297) );
  AOI22_X1 U2684 ( .A1(\UUT/Mpath/the_alu/N22 ), .A2(n1298), .B1(n1299), .B2(
        n1300), .ZN(n1296) );
  INV_X1 U2685 ( .A(\UUT/Mpath/the_alu/N22 ), .ZN(n1300) );
  OAI221_X1 U2686 ( .B1(n1301), .B2(n1302), .C1(\UUT/Mpath/the_alu/N21 ), .C2(
        n1303), .A(n1304), .ZN(n1299) );
  OAI22_X1 U2687 ( .A1(\UUT/Mpath/the_alu/N21 ), .A2(n1301), .B1(n1305), .B2(
        n1302), .ZN(n1298) );
  INV_X1 U2688 ( .A(\UUT/Mpath/the_alu/N21 ), .ZN(n1302) );
  NAND3_X1 U2689 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n6109) );
  AOI222_X1 U2690 ( .A1(\UUT/Mpath/the_alu/sum[3] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N154 ), .B2(n6834), .C1(n1218), .C2(n1309), .ZN(
        n1308) );
  INV_X1 U2691 ( .A(\UUT/Mpath/the_alu/N77 ), .ZN(n1309) );
  AOI22_X1 U2692 ( .A1(\UUT/Mpath/the_alu/N218 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N186 ), .B2(n1221), .ZN(n1307) );
  AOI22_X1 U2693 ( .A1(\UUT/Mpath/the_alu/N122 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[3] ), .B2(n1223), .ZN(n1306) );
  AND2_X1 U2694 ( .A1(n1310), .A2(n1311), .ZN(n6108) );
  AOI222_X1 U2695 ( .A1(\UUT/Mpath/the_shift/sh_rol [3]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [3]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [3]), .C2(n1228), .ZN(n1311) );
  AOI22_X1 U2696 ( .A1(\UUT/Mpath/the_shift/sh_sra [3]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [3]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1310) );
  NAND3_X1 U2697 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n6107) );
  AOI222_X1 U2698 ( .A1(\UUT/Mpath/the_alu/sum[4] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N153 ), .B2(n6834), .C1(n1218), .C2(n1315), .ZN(
        n1314) );
  INV_X1 U2699 ( .A(\UUT/Mpath/the_alu/N75 ), .ZN(n1315) );
  AOI22_X1 U2700 ( .A1(\UUT/Mpath/the_alu/N217 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N185 ), .B2(n1221), .ZN(n1313) );
  AOI22_X1 U2701 ( .A1(\UUT/Mpath/the_alu/N121 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[4] ), .B2(n1223), .ZN(n1312) );
  AND2_X1 U2702 ( .A1(n1316), .A2(n1317), .ZN(n6106) );
  AOI222_X1 U2703 ( .A1(\UUT/Mpath/the_shift/sh_rol [4]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [4]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [4]), .C2(n1228), .ZN(n1317) );
  AOI22_X1 U2704 ( .A1(\UUT/Mpath/the_shift/sh_sra [4]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [4]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1316) );
  NAND3_X1 U2705 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n6105) );
  AOI222_X1 U2706 ( .A1(\UUT/Mpath/the_alu/sum[5] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N152 ), .B2(n6834), .C1(n1218), .C2(n1321), .ZN(
        n1320) );
  AOI22_X1 U2708 ( .A1(\UUT/Mpath/the_alu/N216 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N184 ), .B2(n1221), .ZN(n1319) );
  AOI22_X1 U2709 ( .A1(\UUT/Mpath/the_alu/N120 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[5] ), .B2(n1223), .ZN(n1318) );
  AND2_X1 U2710 ( .A1(n1322), .A2(n1323), .ZN(n6104) );
  AOI222_X1 U2711 ( .A1(\UUT/Mpath/the_shift/sh_rol [5]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [5]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [5]), .C2(n1228), .ZN(n1323) );
  AOI22_X1 U2712 ( .A1(\UUT/Mpath/the_shift/sh_sra [5]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [5]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1322) );
  NAND3_X1 U2713 ( .A1(n1324), .A2(n1325), .A3(n1326), .ZN(n6103) );
  AOI222_X1 U2714 ( .A1(\UUT/Mpath/the_alu/sum[6] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N151 ), .B2(n6834), .C1(n1218), .C2(n1327), .ZN(
        n1326) );
  INV_X1 U2715 ( .A(\UUT/Mpath/the_alu/N71 ), .ZN(n1327) );
  AOI22_X1 U2716 ( .A1(\UUT/Mpath/the_alu/N215 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N183 ), .B2(n1221), .ZN(n1325) );
  AOI22_X1 U2717 ( .A1(\UUT/Mpath/the_alu/N119 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[6] ), .B2(n1223), .ZN(n1324) );
  AND2_X1 U2718 ( .A1(n1328), .A2(n1329), .ZN(n6102) );
  AOI222_X1 U2719 ( .A1(\UUT/Mpath/the_shift/sh_rol [6]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [6]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [6]), .C2(n1228), .ZN(n1329) );
  AOI22_X1 U2720 ( .A1(\UUT/Mpath/the_shift/sh_sra [6]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [6]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1328) );
  NAND3_X1 U2721 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n6101) );
  AOI222_X1 U2722 ( .A1(\UUT/Mpath/the_alu/sum[7] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N150 ), .B2(n6834), .C1(n1218), .C2(n1333), .ZN(
        n1332) );
  INV_X1 U2723 ( .A(\UUT/Mpath/the_alu/N69 ), .ZN(n1333) );
  AOI22_X1 U2724 ( .A1(\UUT/Mpath/the_alu/N214 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N182 ), .B2(n1221), .ZN(n1331) );
  AOI22_X1 U2725 ( .A1(\UUT/Mpath/the_alu/N118 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[7] ), .B2(n1223), .ZN(n1330) );
  AOI222_X1 U2727 ( .A1(\UUT/Mpath/the_shift/sh_rol [7]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [7]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [7]), .C2(n1228), .ZN(n1335) );
  AOI22_X1 U2728 ( .A1(\UUT/Mpath/the_shift/sh_sra [7]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [7]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1334) );
  NAND3_X1 U2729 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n6099) );
  AOI222_X1 U2730 ( .A1(\UUT/Mpath/the_alu/sum[8] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N149 ), .B2(n6834), .C1(n1218), .C2(n1339), .ZN(
        n1338) );
  INV_X1 U2731 ( .A(\UUT/Mpath/the_alu/N67 ), .ZN(n1339) );
  AOI22_X1 U2732 ( .A1(\UUT/Mpath/the_alu/N213 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N181 ), .B2(n1221), .ZN(n1337) );
  AOI22_X1 U2733 ( .A1(\UUT/Mpath/the_alu/N117 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[8] ), .B2(n1223), .ZN(n1336) );
  AND2_X1 U2734 ( .A1(n1340), .A2(n1341), .ZN(n6098) );
  AOI222_X1 U2735 ( .A1(\UUT/Mpath/the_shift/sh_rol [8]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [8]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [8]), .C2(n1228), .ZN(n1341) );
  AOI22_X1 U2736 ( .A1(\UUT/Mpath/the_shift/sh_sra [8]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [8]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1340) );
  NAND3_X1 U2737 ( .A1(n1342), .A2(n1343), .A3(n1344), .ZN(n6097) );
  AOI222_X1 U2738 ( .A1(\UUT/Mpath/the_alu/sum[9] ), .A2(n7213), .B1(
        \UUT/Mpath/the_alu/N148 ), .B2(n6834), .C1(n1218), .C2(n1345), .ZN(
        n1344) );
  INV_X1 U2739 ( .A(\UUT/Mpath/the_alu/N65 ), .ZN(n1345) );
  AOI22_X1 U2740 ( .A1(\UUT/Mpath/the_alu/N212 ), .A2(n1220), .B1(
        \UUT/Mpath/the_alu/N180 ), .B2(n1221), .ZN(n1343) );
  AOI22_X1 U2743 ( .A1(\UUT/Mpath/the_alu/N116 ), .A2(n1222), .B1(
        \UUT/Mpath/the_alu/diff[9] ), .B2(n1223), .ZN(n1342) );
  INV_X1 U2744 ( .A(n1303), .ZN(n1222) );
  AND2_X1 U2745 ( .A1(n1346), .A2(n1347), .ZN(n6096) );
  AOI222_X1 U2746 ( .A1(\UUT/Mpath/the_shift/sh_rol [9]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [9]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [9]), .C2(n1228), .ZN(n1347) );
  AOI22_X1 U2747 ( .A1(\UUT/Mpath/the_shift/sh_sra [9]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [9]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1346) );
  AND2_X1 U2748 ( .A1(n1348), .A2(n1349), .ZN(n6094) );
  AOI222_X1 U2749 ( .A1(\UUT/Mpath/the_shift/sh_rol [13]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [13]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [13]), .C2(n1228), .ZN(n1349) );
  AOI22_X1 U2750 ( .A1(\UUT/Mpath/the_shift/sh_sra [13]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [13]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1348) );
  AND2_X1 U2751 ( .A1(n1350), .A2(n1351), .ZN(n6084) );
  AOI222_X1 U2752 ( .A1(\UUT/Mpath/the_shift/sh_rol [14]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [14]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [14]), .C2(n1228), .ZN(n1351) );
  AOI22_X1 U2753 ( .A1(\UUT/Mpath/the_shift/sh_sra [14]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [14]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1350) );
  AND2_X1 U2754 ( .A1(n1352), .A2(n1353), .ZN(n6070) );
  AOI222_X1 U2755 ( .A1(\UUT/Mpath/the_shift/sh_rol [15]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [15]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [15]), .C2(n1228), .ZN(n1353) );
  AOI22_X1 U2756 ( .A1(\UUT/Mpath/the_shift/sh_sra [15]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [15]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1352) );
  AND2_X1 U2757 ( .A1(n1354), .A2(n1355), .ZN(n6059) );
  AOI222_X1 U2758 ( .A1(\UUT/Mpath/the_shift/sh_rol [16]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [16]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [16]), .C2(n1228), .ZN(n1355) );
  AOI22_X1 U2759 ( .A1(\UUT/Mpath/the_shift/sh_sra [16]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [16]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1354) );
  AND2_X1 U2760 ( .A1(n1356), .A2(n1357), .ZN(n6047) );
  AOI222_X1 U2761 ( .A1(\UUT/Mpath/the_shift/sh_rol [17]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [17]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [17]), .C2(n1228), .ZN(n1357) );
  AOI22_X1 U2762 ( .A1(\UUT/Mpath/the_shift/sh_sra [17]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [17]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1356) );
  AND2_X1 U2763 ( .A1(n1358), .A2(n1359), .ZN(n6026) );
  AOI222_X1 U2764 ( .A1(\UUT/Mpath/the_shift/sh_rol [18]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [18]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [18]), .C2(n1228), .ZN(n1359) );
  AOI22_X1 U2765 ( .A1(\UUT/Mpath/the_shift/sh_sra [18]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [18]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1358) );
  AND2_X1 U2766 ( .A1(n1360), .A2(n1361), .ZN(n6013) );
  AOI222_X1 U2767 ( .A1(\UUT/Mpath/the_shift/sh_rol [19]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [19]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [19]), .C2(n1228), .ZN(n1361) );
  AOI22_X1 U2768 ( .A1(\UUT/Mpath/the_shift/sh_sra [19]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [19]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1360) );
  AND2_X1 U2769 ( .A1(n1362), .A2(n1363), .ZN(n6000) );
  AOI222_X1 U2770 ( .A1(\UUT/Mpath/the_shift/sh_rol [20]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [20]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [20]), .C2(n1228), .ZN(n1363) );
  AOI22_X1 U2771 ( .A1(\UUT/Mpath/the_shift/sh_sra [20]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [20]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1362) );
  AOI222_X1 U2773 ( .A1(\UUT/Mpath/the_shift/sh_rol [21]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [21]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [21]), .C2(n1228), .ZN(n1365) );
  AOI22_X1 U2774 ( .A1(\UUT/Mpath/the_shift/sh_sra [21]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [21]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1364) );
  AOI222_X1 U2776 ( .A1(\UUT/Mpath/the_shift/sh_rol [22]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [22]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [22]), .C2(n1228), .ZN(n1367) );
  AOI22_X1 U2777 ( .A1(\UUT/Mpath/the_shift/sh_sra [22]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [22]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1366) );
  AOI222_X1 U2779 ( .A1(\UUT/Mpath/the_shift/sh_rol [23]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [23]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [23]), .C2(n1228), .ZN(n1369) );
  AOI22_X1 U2780 ( .A1(\UUT/Mpath/the_shift/sh_sra [23]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [23]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1368) );
  AND2_X1 U2781 ( .A1(n1370), .A2(n1371), .ZN(n5958) );
  AOI222_X1 U2782 ( .A1(\UUT/Mpath/the_shift/sh_rol [1]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [1]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [1]), .C2(n1228), .ZN(n1371) );
  AOI22_X1 U2783 ( .A1(\UUT/Mpath/the_shift/sh_sra [1]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [1]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1370) );
  NOR4_X1 U2784 ( .A1(n1372), .A2(n1128), .A3(n5937), .A4(n7117), .ZN(n5946)
         );
  INV_X1 U2785 ( .A(n5917), .ZN(n1128) );
  INV_X1 U2786 ( .A(n7251), .ZN(n1372) );
  NAND3_X1 U2787 ( .A1(n7021), .A2(n6995), .A3(n451), .ZN(n5944) );
  OR2_X1 U2804 ( .A1(\UUT/Mpath/the_memhandle/N120 ), .A2(
        \UUT/Mpath/the_memhandle/N86 ), .ZN(n5825) );
  NAND2_X1 U2805 ( .A1(n5862), .A2(n5856), .ZN(n5823) );
  INV_X1 U2808 ( .A(n5752), .ZN(n5761) );
  NAND2_X1 U2810 ( .A1(n1374), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .ZN(n5754) );
  INV_X1 U2811 ( .A(n6004), .ZN(n1374) );
  AND2_X1 U2813 ( .A1(n1375), .A2(n1376), .ZN(n5526) );
  AOI222_X1 U2814 ( .A1(\UUT/Mpath/the_shift/sh_rol [0]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [0]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [0]), .C2(n1228), .ZN(n1376) );
  AOI22_X1 U2815 ( .A1(\UUT/Mpath/the_shift/sh_sra [0]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [0]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1375) );
  INV_X1 U2816 ( .A(n1377), .ZN(n5516) );
  OAI211_X1 U2817 ( .C1(\UUT/Mpath/the_alu/N35 ), .C2(n7215), .A(n1378), .B(
        n1379), .ZN(n1377) );
  AOI22_X1 U2818 ( .A1(\UUT/Mpath/the_alu/diff[24] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[24] ), .B2(n7213), .ZN(n1379) );
  AOI22_X1 U2819 ( .A1(\UUT/Mpath/the_alu/N36 ), .A2(n1380), .B1(n1381), .B2(
        n1382), .ZN(n1378) );
  INV_X1 U2820 ( .A(\UUT/Mpath/the_alu/N36 ), .ZN(n1382) );
  OAI221_X1 U2821 ( .B1(n1301), .B2(n1383), .C1(\UUT/Mpath/the_alu/N35 ), .C2(
        n1303), .A(n1304), .ZN(n1381) );
  OAI22_X1 U2822 ( .A1(\UUT/Mpath/the_alu/N35 ), .A2(n1301), .B1(n1305), .B2(
        n1383), .ZN(n1380) );
  INV_X1 U2823 ( .A(\UUT/Mpath/the_alu/N35 ), .ZN(n1383) );
  AND2_X1 U2824 ( .A1(n1384), .A2(n1385), .ZN(n5515) );
  AOI222_X1 U2825 ( .A1(\UUT/Mpath/the_shift/sh_rol [24]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [24]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [24]), .C2(n1228), .ZN(n1385) );
  AOI22_X1 U2826 ( .A1(\UUT/Mpath/the_shift/sh_sra [24]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [24]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1384) );
  INV_X1 U2827 ( .A(n1386), .ZN(n5508) );
  OAI211_X1 U2828 ( .C1(\UUT/Mpath/the_alu/N33 ), .C2(n7215), .A(n1387), .B(
        n1388), .ZN(n1386) );
  AOI22_X1 U2829 ( .A1(\UUT/Mpath/the_alu/diff[25] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[25] ), .B2(n7213), .ZN(n1388) );
  AOI22_X1 U2830 ( .A1(\UUT/Mpath/the_alu/N34 ), .A2(n1389), .B1(n1390), .B2(
        n1391), .ZN(n1387) );
  INV_X1 U2831 ( .A(\UUT/Mpath/the_alu/N34 ), .ZN(n1391) );
  OAI221_X1 U2832 ( .B1(n1301), .B2(n1392), .C1(\UUT/Mpath/the_alu/N33 ), .C2(
        n1303), .A(n1304), .ZN(n1390) );
  OAI22_X1 U2833 ( .A1(\UUT/Mpath/the_alu/N33 ), .A2(n1301), .B1(n1305), .B2(
        n1392), .ZN(n1389) );
  INV_X1 U2834 ( .A(\UUT/Mpath/the_alu/N33 ), .ZN(n1392) );
  AND2_X1 U2835 ( .A1(n1393), .A2(n1394), .ZN(n5507) );
  AOI222_X1 U2836 ( .A1(\UUT/Mpath/the_shift/sh_rol [25]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [25]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [25]), .C2(n1228), .ZN(n1394) );
  AOI22_X1 U2837 ( .A1(\UUT/Mpath/the_shift/sh_sra [25]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [25]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1393) );
  INV_X1 U2838 ( .A(n1395), .ZN(n5500) );
  OAI211_X1 U2839 ( .C1(\UUT/Mpath/the_alu/N31 ), .C2(n7215), .A(n1396), .B(
        n1397), .ZN(n1395) );
  AOI22_X1 U2840 ( .A1(\UUT/Mpath/the_alu/diff[26] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[26] ), .B2(n7213), .ZN(n1397) );
  AOI22_X1 U2841 ( .A1(\UUT/Mpath/the_alu/N32 ), .A2(n1398), .B1(n1399), .B2(
        n1400), .ZN(n1396) );
  INV_X1 U2842 ( .A(\UUT/Mpath/the_alu/N32 ), .ZN(n1400) );
  OAI221_X1 U2843 ( .B1(n1301), .B2(n1401), .C1(\UUT/Mpath/the_alu/N31 ), .C2(
        n1303), .A(n1304), .ZN(n1399) );
  OAI22_X1 U2844 ( .A1(\UUT/Mpath/the_alu/N31 ), .A2(n1301), .B1(n1305), .B2(
        n1401), .ZN(n1398) );
  INV_X1 U2845 ( .A(\UUT/Mpath/the_alu/N31 ), .ZN(n1401) );
  AND2_X1 U2846 ( .A1(n1402), .A2(n1403), .ZN(n5499) );
  AOI222_X1 U2847 ( .A1(\UUT/Mpath/the_shift/sh_rol [26]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [26]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [26]), .C2(n1228), .ZN(n1403) );
  AOI22_X1 U2848 ( .A1(\UUT/Mpath/the_shift/sh_sra [26]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [26]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1402) );
  INV_X1 U2849 ( .A(n1404), .ZN(n5492) );
  OAI211_X1 U2850 ( .C1(\UUT/Mpath/the_alu/N29 ), .C2(n7215), .A(n1405), .B(
        n1406), .ZN(n1404) );
  AOI22_X1 U2851 ( .A1(\UUT/Mpath/the_alu/diff[27] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[27] ), .B2(n7213), .ZN(n1406) );
  AOI22_X1 U2852 ( .A1(\UUT/Mpath/the_alu/N30 ), .A2(n1407), .B1(n1408), .B2(
        n1409), .ZN(n1405) );
  INV_X1 U2853 ( .A(\UUT/Mpath/the_alu/N30 ), .ZN(n1409) );
  OAI221_X1 U2854 ( .B1(n1301), .B2(n1410), .C1(\UUT/Mpath/the_alu/N29 ), .C2(
        n1303), .A(n1304), .ZN(n1408) );
  OAI22_X1 U2855 ( .A1(\UUT/Mpath/the_alu/N29 ), .A2(n1301), .B1(n1305), .B2(
        n1410), .ZN(n1407) );
  INV_X1 U2856 ( .A(\UUT/Mpath/the_alu/N29 ), .ZN(n1410) );
  AND2_X1 U2857 ( .A1(n1411), .A2(n1412), .ZN(n5491) );
  AOI222_X1 U2858 ( .A1(\UUT/Mpath/the_shift/sh_rol [27]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [27]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [27]), .C2(n1228), .ZN(n1412) );
  AOI22_X1 U2859 ( .A1(\UUT/Mpath/the_shift/sh_sra [27]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [27]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1411) );
  OAI211_X1 U2861 ( .C1(\UUT/Mpath/the_alu/N27 ), .C2(n7215), .A(n1414), .B(
        n1415), .ZN(n1413) );
  AOI22_X1 U2862 ( .A1(\UUT/Mpath/the_alu/diff[28] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[28] ), .B2(n7213), .ZN(n1415) );
  AOI22_X1 U2863 ( .A1(\UUT/Mpath/the_alu/N28 ), .A2(n1416), .B1(n1417), .B2(
        n1418), .ZN(n1414) );
  INV_X1 U2864 ( .A(\UUT/Mpath/the_alu/N28 ), .ZN(n1418) );
  OAI221_X1 U2865 ( .B1(n1301), .B2(n1419), .C1(\UUT/Mpath/the_alu/N27 ), .C2(
        n1303), .A(n1304), .ZN(n1417) );
  OAI22_X1 U2866 ( .A1(\UUT/Mpath/the_alu/N27 ), .A2(n1301), .B1(n1305), .B2(
        n1419), .ZN(n1416) );
  INV_X1 U2867 ( .A(\UUT/Mpath/the_alu/N27 ), .ZN(n1419) );
  AND2_X1 U2868 ( .A1(n1420), .A2(n1421), .ZN(n5483) );
  AOI222_X1 U2869 ( .A1(\UUT/Mpath/the_shift/sh_rol [28]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [28]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [28]), .C2(n1228), .ZN(n1421) );
  AOI22_X1 U2870 ( .A1(\UUT/Mpath/the_shift/sh_sra [28]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [28]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1420) );
  OAI211_X1 U2872 ( .C1(\UUT/Mpath/the_alu/N25 ), .C2(n7215), .A(n1423), .B(
        n1424), .ZN(n1422) );
  AOI22_X1 U2874 ( .A1(\UUT/Mpath/the_alu/N26 ), .A2(n1425), .B1(n1426), .B2(
        n1427), .ZN(n1423) );
  INV_X1 U2875 ( .A(\UUT/Mpath/the_alu/N26 ), .ZN(n1427) );
  OAI221_X1 U2876 ( .B1(n1301), .B2(n1428), .C1(\UUT/Mpath/the_alu/N25 ), .C2(
        n1303), .A(n1304), .ZN(n1426) );
  OAI22_X1 U2877 ( .A1(\UUT/Mpath/the_alu/N25 ), .A2(n1301), .B1(n1305), .B2(
        n1428), .ZN(n1425) );
  INV_X1 U2878 ( .A(\UUT/Mpath/the_alu/N25 ), .ZN(n1428) );
  AND2_X1 U2879 ( .A1(n1429), .A2(n1430), .ZN(n5475) );
  AOI222_X1 U2880 ( .A1(\UUT/Mpath/the_shift/sh_rol [29]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [29]), .B2(n6343), .C1(
        \UUT/Mpath/the_shift/sh_sll [29]), .C2(n1228), .ZN(n1430) );
  AOI22_X1 U2881 ( .A1(\UUT/Mpath/the_shift/sh_sra [29]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [29]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1429) );
  INV_X1 U2882 ( .A(n1431), .ZN(n5467) );
  OAI211_X1 U2883 ( .C1(\UUT/Mpath/the_alu/N23 ), .C2(n7215), .A(n1432), .B(
        n1433), .ZN(n1431) );
  AOI22_X1 U2885 ( .A1(\UUT/Mpath/the_alu/N24 ), .A2(n1434), .B1(n1435), .B2(
        n1436), .ZN(n1432) );
  INV_X1 U2886 ( .A(\UUT/Mpath/the_alu/N24 ), .ZN(n1436) );
  OAI221_X1 U2887 ( .B1(n1301), .B2(n1437), .C1(\UUT/Mpath/the_alu/N23 ), .C2(
        n1303), .A(n1304), .ZN(n1435) );
  OAI22_X1 U2888 ( .A1(\UUT/Mpath/the_alu/N23 ), .A2(n1301), .B1(n1305), .B2(
        n1437), .ZN(n1434) );
  INV_X1 U2889 ( .A(\UUT/Mpath/the_alu/N23 ), .ZN(n1437) );
  AOI222_X1 U2891 ( .A1(\UUT/Mpath/the_shift/sh_rol [30]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [30]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [30]), .C2(n1228), .ZN(n1439) );
  INV_X1 U2894 ( .A(\UUT/Mpath/the_shift/N111 ), .ZN(n1440) );
  INV_X1 U2896 ( .A(n6282), .ZN(n1441) );
  AOI22_X1 U2897 ( .A1(\UUT/Mpath/the_shift/sh_sra [30]), .A2(n1229), .B1(
        \UUT/Mpath/the_shift/sh_srl [30]), .B2(\UUT/Mpath/the_shift/N118 ), 
        .ZN(n1438) );
  INV_X1 U2899 ( .A(\UUT/Mpath/the_shift/N115 ), .ZN(n1442) );
  AND4_X1 U2900 ( .A1(n1443), .A2(n1444), .A3(n1445), .A4(n1446), .ZN(n5428)
         );
  NOR4_X1 U2901 ( .A1(n1447), .A2(n1448), .A3(n1449), .A4(n1450), .ZN(n1446)
         );
  NAND3_X1 U2902 ( .A1(n5889), .A2(n5885), .A3(n5894), .ZN(n1450) );
  OAI211_X1 U2903 ( .C1(n5656), .C2(n5314), .A(n5874), .B(n5881), .ZN(n1449)
         );
  OAI222_X1 U2904 ( .A1(n5654), .A2(n5186), .B1(n5655), .B2(n5154), .C1(n5657), 
        .C2(n5282), .ZN(n1448) );
  OAI221_X1 U2905 ( .B1(n6925), .B2(n5090), .C1(n6352), .C2(n5122), .A(n1451), 
        .ZN(n1447) );
  AOI22_X1 U2906 ( .A1(n1452), .A2(n1453), .B1(n1454), .B2(n1455), .ZN(n1451)
         );
  AOI211_X1 U2907 ( .C1(n1456), .C2(n1457), .A(n1458), .B(n1459), .ZN(n1445)
         );
  OAI22_X1 U2908 ( .A1(n5637), .A2(n4738), .B1(n5647), .B2(n4642), .ZN(n1459)
         );
  OAI222_X1 U2909 ( .A1(n5642), .A2(n4578), .B1(n5648), .B2(n4546), .C1(n6936), 
        .C2(n4610), .ZN(n1458) );
  AOI221_X1 U2910 ( .B1(n6348), .B2(n1461), .C1(n1462), .C2(n1463), .A(n1464), 
        .ZN(n1444) );
  OAI22_X1 U2911 ( .A1(n4386), .A2(n1465), .B1(n5218), .B2(n1466), .ZN(n1464)
         );
  AOI222_X1 U2913 ( .A1(n1467), .A2(n1468), .B1(n1469), .B2(n1470), .C1(n1471), 
        .C2(n1472), .ZN(n1443) );
  AND4_X1 U2914 ( .A1(n1473), .A2(n1474), .A3(n1475), .A4(n1476), .ZN(n5425)
         );
  NOR4_X1 U2915 ( .A1(n1477), .A2(n1478), .A3(n1479), .A4(n1480), .ZN(n1476)
         );
  NAND3_X1 U2916 ( .A1(n5866), .A2(n5865), .A3(n5867), .ZN(n1480) );
  OAI211_X1 U2917 ( .C1(n5656), .C2(n5313), .A(n5863), .B(n5864), .ZN(n1479)
         );
  OAI222_X1 U2918 ( .A1(n5654), .A2(n5185), .B1(n5655), .B2(n5153), .C1(n5657), 
        .C2(n5281), .ZN(n1478) );
  OAI221_X1 U2919 ( .B1(n6925), .B2(n5089), .C1(n6353), .C2(n5121), .A(n1481), 
        .ZN(n1477) );
  AOI22_X1 U2920 ( .A1(n1482), .A2(n1453), .B1(n1483), .B2(n1455), .ZN(n1481)
         );
  AOI211_X1 U2921 ( .C1(n1484), .C2(n1457), .A(n1485), .B(n1486), .ZN(n1475)
         );
  OAI22_X1 U2922 ( .A1(n5637), .A2(n4737), .B1(n5647), .B2(n4641), .ZN(n1486)
         );
  OAI222_X1 U2923 ( .A1(n5642), .A2(n4577), .B1(n5648), .B2(n4545), .C1(n6936), 
        .C2(n4609), .ZN(n1485) );
  AOI221_X1 U2924 ( .B1(n6349), .B2(n1487), .C1(n1462), .C2(n1488), .A(n1489), 
        .ZN(n1474) );
  OAI22_X1 U2925 ( .A1(n4385), .A2(n1465), .B1(n5217), .B2(n1466), .ZN(n1489)
         );
  AOI222_X1 U2927 ( .A1(n1490), .A2(n1468), .B1(n1469), .B2(n1491), .C1(n1492), 
        .C2(n1472), .ZN(n1473) );
  AND4_X1 U2928 ( .A1(n1493), .A2(n1494), .A3(n1495), .A4(n1496), .ZN(n5422)
         );
  NOR4_X1 U2929 ( .A1(n1497), .A2(n1498), .A3(n1499), .A4(n1500), .ZN(n1496)
         );
  NAND3_X1 U2930 ( .A1(n5854), .A2(n5853), .A3(n5855), .ZN(n1500) );
  OAI211_X1 U2931 ( .C1(n5656), .C2(n5312), .A(n5851), .B(n5852), .ZN(n1499)
         );
  OAI222_X1 U2932 ( .A1(n5654), .A2(n5184), .B1(n5655), .B2(n5152), .C1(n5657), 
        .C2(n5280), .ZN(n1498) );
  OAI221_X1 U2933 ( .B1(n6925), .B2(n5088), .C1(n6353), .C2(n5120), .A(n1501), 
        .ZN(n1497) );
  AOI22_X1 U2934 ( .A1(n1502), .A2(n1453), .B1(n1503), .B2(n1455), .ZN(n1501)
         );
  AOI211_X1 U2935 ( .C1(n1504), .C2(n1457), .A(n1505), .B(n1506), .ZN(n1495)
         );
  OAI22_X1 U2936 ( .A1(n5637), .A2(n4736), .B1(n5647), .B2(n4640), .ZN(n1506)
         );
  OAI222_X1 U2937 ( .A1(n5642), .A2(n4576), .B1(n5648), .B2(n4544), .C1(n6936), 
        .C2(n4608), .ZN(n1505) );
  AOI221_X1 U2938 ( .B1(n6349), .B2(n1507), .C1(n1462), .C2(n1508), .A(n1509), 
        .ZN(n1494) );
  OAI22_X1 U2939 ( .A1(n4384), .A2(n1465), .B1(n5216), .B2(n1466), .ZN(n1509)
         );
  AOI222_X1 U2941 ( .A1(n1510), .A2(n1468), .B1(n1469), .B2(n1511), .C1(n1512), 
        .C2(n1472), .ZN(n1493) );
  AND4_X1 U2942 ( .A1(n1513), .A2(n1514), .A3(n1515), .A4(n1516), .ZN(n5419)
         );
  NOR4_X1 U2943 ( .A1(n1517), .A2(n1518), .A3(n1519), .A4(n1520), .ZN(n1516)
         );
  NAND3_X1 U2944 ( .A1(n5849), .A2(n5848), .A3(n5850), .ZN(n1520) );
  OAI211_X1 U2945 ( .C1(n5656), .C2(n5311), .A(n5846), .B(n5847), .ZN(n1519)
         );
  OAI222_X1 U2946 ( .A1(n5654), .A2(n5183), .B1(n5655), .B2(n5151), .C1(n5657), 
        .C2(n5279), .ZN(n1518) );
  OAI221_X1 U2947 ( .B1(n6925), .B2(n5087), .C1(n6353), .C2(n5119), .A(n1521), 
        .ZN(n1517) );
  AOI22_X1 U2948 ( .A1(n1522), .A2(n1453), .B1(n1523), .B2(n1455), .ZN(n1521)
         );
  AOI211_X1 U2949 ( .C1(n1524), .C2(n1457), .A(n1525), .B(n1526), .ZN(n1515)
         );
  OAI22_X1 U2950 ( .A1(n5637), .A2(n4735), .B1(n5647), .B2(n4639), .ZN(n1526)
         );
  OAI222_X1 U2951 ( .A1(n5642), .A2(n4575), .B1(n5648), .B2(n4543), .C1(n6936), 
        .C2(n4607), .ZN(n1525) );
  AOI221_X1 U2952 ( .B1(n6349), .B2(n1527), .C1(n1462), .C2(n1528), .A(n1529), 
        .ZN(n1514) );
  OAI22_X1 U2953 ( .A1(n4383), .A2(n1465), .B1(n5215), .B2(n1466), .ZN(n1529)
         );
  AOI222_X1 U2955 ( .A1(n1530), .A2(n1468), .B1(n1469), .B2(n1531), .C1(n1532), 
        .C2(n1472), .ZN(n1513) );
  AND4_X1 U2956 ( .A1(n1533), .A2(n1534), .A3(n1535), .A4(n1536), .ZN(n5416)
         );
  NOR4_X1 U2957 ( .A1(n1537), .A2(n1538), .A3(n1539), .A4(n1540), .ZN(n1536)
         );
  NAND3_X1 U2958 ( .A1(n5844), .A2(n5843), .A3(n5845), .ZN(n1540) );
  OAI211_X1 U2959 ( .C1(n5656), .C2(n5310), .A(n5841), .B(n5842), .ZN(n1539)
         );
  OAI222_X1 U2960 ( .A1(n5654), .A2(n5182), .B1(n5655), .B2(n5150), .C1(n5657), 
        .C2(n5278), .ZN(n1538) );
  OAI221_X1 U2961 ( .B1(n6925), .B2(n5086), .C1(n6352), .C2(n5118), .A(n1541), 
        .ZN(n1537) );
  AOI22_X1 U2962 ( .A1(n1542), .A2(n1453), .B1(n1543), .B2(n1455), .ZN(n1541)
         );
  AOI211_X1 U2963 ( .C1(n1544), .C2(n1457), .A(n1545), .B(n1546), .ZN(n1535)
         );
  OAI22_X1 U2964 ( .A1(n5637), .A2(n4734), .B1(n5647), .B2(n4638), .ZN(n1546)
         );
  OAI222_X1 U2965 ( .A1(n5642), .A2(n4574), .B1(n5648), .B2(n4542), .C1(n6936), 
        .C2(n4606), .ZN(n1545) );
  AOI221_X1 U2966 ( .B1(n6348), .B2(n1547), .C1(n1462), .C2(n1548), .A(n1549), 
        .ZN(n1534) );
  OAI22_X1 U2967 ( .A1(n4382), .A2(n1465), .B1(n5214), .B2(n1466), .ZN(n1549)
         );
  AOI222_X1 U2969 ( .A1(n1550), .A2(n1468), .B1(n1469), .B2(n1551), .C1(n1552), 
        .C2(n1472), .ZN(n1533) );
  AND4_X1 U2970 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .ZN(n5413)
         );
  NOR4_X1 U2971 ( .A1(n1557), .A2(n1558), .A3(n1559), .A4(n1560), .ZN(n1556)
         );
  NAND3_X1 U2972 ( .A1(n5839), .A2(n5838), .A3(n5840), .ZN(n1560) );
  OAI211_X1 U2973 ( .C1(n5656), .C2(n5309), .A(n5836), .B(n5837), .ZN(n1559)
         );
  OAI222_X1 U2974 ( .A1(n5654), .A2(n5181), .B1(n5655), .B2(n5149), .C1(n5657), 
        .C2(n5277), .ZN(n1558) );
  OAI221_X1 U2975 ( .B1(n6925), .B2(n5085), .C1(n6352), .C2(n5117), .A(n1561), 
        .ZN(n1557) );
  AOI22_X1 U2976 ( .A1(n1562), .A2(n1453), .B1(n1563), .B2(n1455), .ZN(n1561)
         );
  AOI211_X1 U2977 ( .C1(n1564), .C2(n1457), .A(n1565), .B(n1566), .ZN(n1555)
         );
  OAI22_X1 U2978 ( .A1(n5637), .A2(n4733), .B1(n5647), .B2(n4637), .ZN(n1566)
         );
  OAI222_X1 U2979 ( .A1(n5642), .A2(n4573), .B1(n5648), .B2(n4541), .C1(n6936), 
        .C2(n4605), .ZN(n1565) );
  AOI221_X1 U2980 ( .B1(n6349), .B2(n1567), .C1(n1462), .C2(n1568), .A(n1569), 
        .ZN(n1554) );
  OAI22_X1 U2981 ( .A1(n4381), .A2(n1465), .B1(n5213), .B2(n1466), .ZN(n1569)
         );
  AOI222_X1 U2983 ( .A1(n1570), .A2(n1468), .B1(n1469), .B2(n1571), .C1(n1572), 
        .C2(n1472), .ZN(n1553) );
  AND4_X1 U2984 ( .A1(n1573), .A2(n1574), .A3(n1575), .A4(n1576), .ZN(n5410)
         );
  NOR4_X1 U2985 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .ZN(n1576)
         );
  NAND3_X1 U2986 ( .A1(n5834), .A2(n5833), .A3(n5835), .ZN(n1580) );
  OAI211_X1 U2987 ( .C1(n5656), .C2(n5308), .A(n5831), .B(n5832), .ZN(n1579)
         );
  OAI222_X1 U2988 ( .A1(n5654), .A2(n5180), .B1(n5655), .B2(n5148), .C1(n5657), 
        .C2(n5276), .ZN(n1578) );
  OAI221_X1 U2989 ( .B1(n6925), .B2(n5084), .C1(n6353), .C2(n5116), .A(n1581), 
        .ZN(n1577) );
  AOI22_X1 U2990 ( .A1(n1582), .A2(n1453), .B1(n1583), .B2(n1455), .ZN(n1581)
         );
  AOI211_X1 U2991 ( .C1(n1584), .C2(n1457), .A(n1585), .B(n1586), .ZN(n1575)
         );
  OAI22_X1 U2992 ( .A1(n5637), .A2(n4732), .B1(n5647), .B2(n4636), .ZN(n1586)
         );
  OAI222_X1 U2993 ( .A1(n5642), .A2(n4572), .B1(n5648), .B2(n4540), .C1(n6936), 
        .C2(n4604), .ZN(n1585) );
  AOI221_X1 U2994 ( .B1(n6348), .B2(n1587), .C1(n1462), .C2(n1588), .A(n1589), 
        .ZN(n1574) );
  OAI22_X1 U2995 ( .A1(n4380), .A2(n1465), .B1(n5212), .B2(n1466), .ZN(n1589)
         );
  AOI222_X1 U2997 ( .A1(n1590), .A2(n1468), .B1(n1469), .B2(n1591), .C1(n1592), 
        .C2(n1472), .ZN(n1573) );
  AND4_X1 U2998 ( .A1(n1593), .A2(n1594), .A3(n1595), .A4(n1596), .ZN(n5407)
         );
  NOR4_X1 U2999 ( .A1(n1597), .A2(n1598), .A3(n1599), .A4(n1600), .ZN(n1596)
         );
  NAND3_X1 U3000 ( .A1(n5829), .A2(n5828), .A3(n5830), .ZN(n1600) );
  OAI211_X1 U3001 ( .C1(n5656), .C2(n5307), .A(n5826), .B(n5827), .ZN(n1599)
         );
  OAI222_X1 U3002 ( .A1(n5654), .A2(n5179), .B1(n5655), .B2(n5147), .C1(n5657), 
        .C2(n5275), .ZN(n1598) );
  OAI221_X1 U3003 ( .B1(n6925), .B2(n5083), .C1(n6353), .C2(n5115), .A(n1601), 
        .ZN(n1597) );
  AOI22_X1 U3004 ( .A1(n1602), .A2(n1453), .B1(n1603), .B2(n1455), .ZN(n1601)
         );
  AOI211_X1 U3005 ( .C1(n1604), .C2(n1457), .A(n1605), .B(n1606), .ZN(n1595)
         );
  OAI22_X1 U3006 ( .A1(n5637), .A2(n4731), .B1(n5647), .B2(n4635), .ZN(n1606)
         );
  OAI222_X1 U3007 ( .A1(n5642), .A2(n4571), .B1(n5648), .B2(n4539), .C1(n6936), 
        .C2(n4603), .ZN(n1605) );
  AOI221_X1 U3008 ( .B1(n6349), .B2(n1607), .C1(n1462), .C2(n1608), .A(n1609), 
        .ZN(n1594) );
  OAI22_X1 U3009 ( .A1(n4379), .A2(n1465), .B1(n5211), .B2(n1466), .ZN(n1609)
         );
  AOI222_X1 U3011 ( .A1(n1610), .A2(n1468), .B1(n1469), .B2(n1611), .C1(n1612), 
        .C2(n1472), .ZN(n1593) );
  AND4_X1 U3012 ( .A1(n1613), .A2(n1614), .A3(n1615), .A4(n1616), .ZN(n5404)
         );
  NOR4_X1 U3013 ( .A1(n1617), .A2(n1618), .A3(n1619), .A4(n1620), .ZN(n1616)
         );
  NAND3_X1 U3014 ( .A1(n5820), .A2(n5819), .A3(n5821), .ZN(n1620) );
  OAI211_X1 U3015 ( .C1(n5656), .C2(n5306), .A(n5817), .B(n5818), .ZN(n1619)
         );
  OAI222_X1 U3016 ( .A1(n5654), .A2(n5178), .B1(n5655), .B2(n5146), .C1(n5657), 
        .C2(n5274), .ZN(n1618) );
  OAI221_X1 U3017 ( .B1(n6925), .B2(n5082), .C1(n6352), .C2(n5114), .A(n1621), 
        .ZN(n1617) );
  AOI22_X1 U3018 ( .A1(n1622), .A2(n1453), .B1(n1623), .B2(n1455), .ZN(n1621)
         );
  AOI211_X1 U3019 ( .C1(n1624), .C2(n1457), .A(n1625), .B(n1626), .ZN(n1615)
         );
  OAI22_X1 U3020 ( .A1(n5637), .A2(n4730), .B1(n5647), .B2(n4634), .ZN(n1626)
         );
  OAI222_X1 U3021 ( .A1(n5642), .A2(n4570), .B1(n5648), .B2(n4538), .C1(n6936), 
        .C2(n4602), .ZN(n1625) );
  AOI221_X1 U3022 ( .B1(n6348), .B2(n1627), .C1(n1462), .C2(n1628), .A(n1629), 
        .ZN(n1614) );
  OAI22_X1 U3023 ( .A1(n4378), .A2(n1465), .B1(n5210), .B2(n1466), .ZN(n1629)
         );
  AOI222_X1 U3025 ( .A1(n1630), .A2(n1468), .B1(n1469), .B2(n1631), .C1(n1632), 
        .C2(n1472), .ZN(n1613) );
  AND4_X1 U3026 ( .A1(n1633), .A2(n1634), .A3(n1635), .A4(n1636), .ZN(n5401)
         );
  NOR4_X1 U3027 ( .A1(n1637), .A2(n1638), .A3(n1639), .A4(n1640), .ZN(n1636)
         );
  NAND3_X1 U3028 ( .A1(n5815), .A2(n5814), .A3(n5816), .ZN(n1640) );
  OAI211_X1 U3029 ( .C1(n5656), .C2(n5305), .A(n5812), .B(n5813), .ZN(n1639)
         );
  OAI222_X1 U3030 ( .A1(n5654), .A2(n5177), .B1(n5655), .B2(n5145), .C1(n5657), 
        .C2(n5273), .ZN(n1638) );
  OAI221_X1 U3031 ( .B1(n6925), .B2(n5081), .C1(n6352), .C2(n5113), .A(n1641), 
        .ZN(n1637) );
  AOI22_X1 U3032 ( .A1(n1642), .A2(n1453), .B1(n1643), .B2(n1455), .ZN(n1641)
         );
  AOI211_X1 U3033 ( .C1(n1644), .C2(n1457), .A(n1645), .B(n1646), .ZN(n1635)
         );
  OAI22_X1 U3034 ( .A1(n5637), .A2(n4729), .B1(n5647), .B2(n4633), .ZN(n1646)
         );
  OAI222_X1 U3035 ( .A1(n5642), .A2(n4569), .B1(n5648), .B2(n4537), .C1(n6936), 
        .C2(n4601), .ZN(n1645) );
  AOI221_X1 U3036 ( .B1(n6348), .B2(n1647), .C1(n1462), .C2(n1648), .A(n1649), 
        .ZN(n1634) );
  OAI22_X1 U3037 ( .A1(n4377), .A2(n1465), .B1(n5209), .B2(n1466), .ZN(n1649)
         );
  AOI222_X1 U3039 ( .A1(n1650), .A2(n1468), .B1(n1469), .B2(n1651), .C1(n1652), 
        .C2(n1472), .ZN(n1633) );
  AND4_X1 U3040 ( .A1(n1653), .A2(n1654), .A3(n1655), .A4(n1656), .ZN(n5398)
         );
  NOR4_X1 U3041 ( .A1(n1657), .A2(n1658), .A3(n1659), .A4(n1660), .ZN(n1656)
         );
  NAND3_X1 U3042 ( .A1(n5810), .A2(n5809), .A3(n5811), .ZN(n1660) );
  OAI211_X1 U3043 ( .C1(n5656), .C2(n5304), .A(n5807), .B(n5808), .ZN(n1659)
         );
  OAI222_X1 U3044 ( .A1(n5654), .A2(n5176), .B1(n5655), .B2(n5144), .C1(n5657), 
        .C2(n5272), .ZN(n1658) );
  OAI221_X1 U3045 ( .B1(n6925), .B2(n5080), .C1(n6352), .C2(n5112), .A(n1661), 
        .ZN(n1657) );
  AOI22_X1 U3046 ( .A1(n1662), .A2(n1453), .B1(n1663), .B2(n1455), .ZN(n1661)
         );
  AOI211_X1 U3047 ( .C1(n1664), .C2(n1457), .A(n1665), .B(n1666), .ZN(n1655)
         );
  OAI22_X1 U3048 ( .A1(n5637), .A2(n4728), .B1(n5647), .B2(n4632), .ZN(n1666)
         );
  OAI222_X1 U3049 ( .A1(n5642), .A2(n4568), .B1(n5648), .B2(n4536), .C1(n6936), 
        .C2(n4600), .ZN(n1665) );
  AOI221_X1 U3050 ( .B1(n6348), .B2(n1667), .C1(n1462), .C2(n1668), .A(n1669), 
        .ZN(n1654) );
  OAI22_X1 U3051 ( .A1(n4376), .A2(n1465), .B1(n5208), .B2(n1466), .ZN(n1669)
         );
  AOI222_X1 U3053 ( .A1(n1670), .A2(n1468), .B1(n1469), .B2(n1671), .C1(n1672), 
        .C2(n1472), .ZN(n1653) );
  AND4_X1 U3054 ( .A1(n1673), .A2(n1674), .A3(n1675), .A4(n1676), .ZN(n5395)
         );
  NOR4_X1 U3055 ( .A1(n1677), .A2(n1678), .A3(n1679), .A4(n1680), .ZN(n1676)
         );
  NAND3_X1 U3056 ( .A1(n5805), .A2(n5804), .A3(n5806), .ZN(n1680) );
  OAI211_X1 U3057 ( .C1(n5656), .C2(n5303), .A(n5802), .B(n5803), .ZN(n1679)
         );
  OAI222_X1 U3058 ( .A1(n5654), .A2(n5175), .B1(n5655), .B2(n5143), .C1(n5657), 
        .C2(n5271), .ZN(n1678) );
  OAI221_X1 U3059 ( .B1(n6925), .B2(n5079), .C1(n6352), .C2(n5111), .A(n1681), 
        .ZN(n1677) );
  AOI22_X1 U3060 ( .A1(n1682), .A2(n1453), .B1(n1683), .B2(n1455), .ZN(n1681)
         );
  AOI211_X1 U3061 ( .C1(n1684), .C2(n1457), .A(n1685), .B(n1686), .ZN(n1675)
         );
  OAI22_X1 U3062 ( .A1(n5637), .A2(n4727), .B1(n5647), .B2(n4631), .ZN(n1686)
         );
  OAI222_X1 U3063 ( .A1(n5642), .A2(n4567), .B1(n5648), .B2(n4535), .C1(n6936), 
        .C2(n4599), .ZN(n1685) );
  AOI221_X1 U3064 ( .B1(n6348), .B2(n1687), .C1(n1462), .C2(n1688), .A(n1689), 
        .ZN(n1674) );
  OAI22_X1 U3065 ( .A1(n4375), .A2(n1465), .B1(n5207), .B2(n1466), .ZN(n1689)
         );
  AOI222_X1 U3067 ( .A1(n1690), .A2(n1468), .B1(n1469), .B2(n1691), .C1(n1692), 
        .C2(n1472), .ZN(n1673) );
  AND4_X1 U3068 ( .A1(n1693), .A2(n1694), .A3(n1695), .A4(n1696), .ZN(n5392)
         );
  NOR4_X1 U3069 ( .A1(n1697), .A2(n1698), .A3(n1699), .A4(n1700), .ZN(n1696)
         );
  NAND3_X1 U3070 ( .A1(n5795), .A2(n5794), .A3(n5796), .ZN(n1700) );
  OAI211_X1 U3071 ( .C1(n5656), .C2(n5302), .A(n5792), .B(n5793), .ZN(n1699)
         );
  OAI222_X1 U3072 ( .A1(n5654), .A2(n5174), .B1(n5655), .B2(n5142), .C1(n5657), 
        .C2(n5270), .ZN(n1698) );
  OAI221_X1 U3073 ( .B1(n6925), .B2(n5078), .C1(n6353), .C2(n5110), .A(n1701), 
        .ZN(n1697) );
  AOI22_X1 U3074 ( .A1(n1702), .A2(n1453), .B1(n1703), .B2(n1455), .ZN(n1701)
         );
  AOI211_X1 U3075 ( .C1(n1704), .C2(n1457), .A(n1705), .B(n1706), .ZN(n1695)
         );
  OAI22_X1 U3076 ( .A1(n5637), .A2(n4726), .B1(n5647), .B2(n4630), .ZN(n1706)
         );
  OAI222_X1 U3077 ( .A1(n5642), .A2(n4566), .B1(n5648), .B2(n4534), .C1(n6936), 
        .C2(n4598), .ZN(n1705) );
  AOI221_X1 U3078 ( .B1(n6349), .B2(n1707), .C1(n1462), .C2(n1708), .A(n1709), 
        .ZN(n1694) );
  OAI22_X1 U3079 ( .A1(n4374), .A2(n1465), .B1(n5206), .B2(n1466), .ZN(n1709)
         );
  AOI222_X1 U3081 ( .A1(n1710), .A2(n1468), .B1(n1469), .B2(n1711), .C1(n1712), 
        .C2(n1472), .ZN(n1693) );
  AND4_X1 U3082 ( .A1(n1713), .A2(n1714), .A3(n1715), .A4(n1716), .ZN(n5389)
         );
  NOR4_X1 U3083 ( .A1(n1717), .A2(n1718), .A3(n1719), .A4(n1720), .ZN(n1716)
         );
  NAND3_X1 U3084 ( .A1(n5790), .A2(n5789), .A3(n5791), .ZN(n1720) );
  OAI211_X1 U3085 ( .C1(n5656), .C2(n5301), .A(n5787), .B(n5788), .ZN(n1719)
         );
  OAI222_X1 U3086 ( .A1(n5654), .A2(n5173), .B1(n5655), .B2(n5141), .C1(n5657), 
        .C2(n5269), .ZN(n1718) );
  OAI221_X1 U3087 ( .B1(n6925), .B2(n5077), .C1(n6352), .C2(n5109), .A(n1721), 
        .ZN(n1717) );
  AOI22_X1 U3088 ( .A1(n1722), .A2(n1453), .B1(n1723), .B2(n1455), .ZN(n1721)
         );
  AOI211_X1 U3089 ( .C1(n1724), .C2(n1457), .A(n1725), .B(n1726), .ZN(n1715)
         );
  OAI22_X1 U3090 ( .A1(n5637), .A2(n4725), .B1(n5647), .B2(n4629), .ZN(n1726)
         );
  OAI222_X1 U3091 ( .A1(n5642), .A2(n4565), .B1(n5648), .B2(n4533), .C1(n6936), 
        .C2(n4597), .ZN(n1725) );
  AOI221_X1 U3092 ( .B1(n6348), .B2(n1727), .C1(n1462), .C2(n1728), .A(n1729), 
        .ZN(n1714) );
  OAI22_X1 U3093 ( .A1(n4373), .A2(n1465), .B1(n5205), .B2(n1466), .ZN(n1729)
         );
  AOI222_X1 U3095 ( .A1(n1730), .A2(n1468), .B1(n1469), .B2(n1731), .C1(n1732), 
        .C2(n1472), .ZN(n1713) );
  AND4_X1 U3096 ( .A1(n1733), .A2(n1734), .A3(n1735), .A4(n1736), .ZN(n5386)
         );
  NOR4_X1 U3097 ( .A1(n1737), .A2(n1738), .A3(n1739), .A4(n1740), .ZN(n1736)
         );
  NAND3_X1 U3098 ( .A1(n5785), .A2(n5784), .A3(n5786), .ZN(n1740) );
  OAI211_X1 U3099 ( .C1(n5656), .C2(n5300), .A(n5782), .B(n5783), .ZN(n1739)
         );
  OAI222_X1 U3100 ( .A1(n5654), .A2(n5172), .B1(n5655), .B2(n5140), .C1(n5657), 
        .C2(n5268), .ZN(n1738) );
  OAI221_X1 U3101 ( .B1(n6925), .B2(n5076), .C1(n6353), .C2(n5108), .A(n1741), 
        .ZN(n1737) );
  AOI22_X1 U3102 ( .A1(n1742), .A2(n1453), .B1(n1743), .B2(n1455), .ZN(n1741)
         );
  AOI211_X1 U3103 ( .C1(n1744), .C2(n1457), .A(n1745), .B(n1746), .ZN(n1735)
         );
  OAI22_X1 U3104 ( .A1(n5637), .A2(n4724), .B1(n5647), .B2(n4628), .ZN(n1746)
         );
  OAI222_X1 U3105 ( .A1(n5642), .A2(n4564), .B1(n5648), .B2(n4532), .C1(n6936), 
        .C2(n4596), .ZN(n1745) );
  AOI221_X1 U3106 ( .B1(n6349), .B2(n1747), .C1(n1462), .C2(n1748), .A(n1749), 
        .ZN(n1734) );
  OAI22_X1 U3107 ( .A1(n4372), .A2(n1465), .B1(n5204), .B2(n1466), .ZN(n1749)
         );
  AOI222_X1 U3109 ( .A1(n1750), .A2(n1468), .B1(n1469), .B2(n1751), .C1(n1752), 
        .C2(n1472), .ZN(n1733) );
  AND4_X1 U3110 ( .A1(n1753), .A2(n1754), .A3(n1755), .A4(n1756), .ZN(n5383)
         );
  NOR4_X1 U3111 ( .A1(n1757), .A2(n1758), .A3(n1759), .A4(n1760), .ZN(n1756)
         );
  NAND3_X1 U3112 ( .A1(n5780), .A2(n5779), .A3(n5781), .ZN(n1760) );
  OAI211_X1 U3113 ( .C1(n5656), .C2(n5299), .A(n5777), .B(n5778), .ZN(n1759)
         );
  OAI222_X1 U3114 ( .A1(n5654), .A2(n5171), .B1(n5655), .B2(n5139), .C1(n5657), 
        .C2(n5267), .ZN(n1758) );
  OAI221_X1 U3115 ( .B1(n6925), .B2(n5075), .C1(n6353), .C2(n5107), .A(n1761), 
        .ZN(n1757) );
  AOI22_X1 U3116 ( .A1(n1762), .A2(n1453), .B1(n1763), .B2(n1455), .ZN(n1761)
         );
  AOI211_X1 U3117 ( .C1(n1764), .C2(n1457), .A(n1765), .B(n1766), .ZN(n1755)
         );
  OAI22_X1 U3118 ( .A1(n5637), .A2(n4723), .B1(n5647), .B2(n4627), .ZN(n1766)
         );
  OAI222_X1 U3119 ( .A1(n5642), .A2(n4563), .B1(n5648), .B2(n4531), .C1(n6936), 
        .C2(n4595), .ZN(n1765) );
  AOI221_X1 U3120 ( .B1(n6348), .B2(n1767), .C1(n1462), .C2(n1768), .A(n1769), 
        .ZN(n1754) );
  OAI22_X1 U3121 ( .A1(n4371), .A2(n1465), .B1(n5203), .B2(n1466), .ZN(n1769)
         );
  AOI222_X1 U3123 ( .A1(n1770), .A2(n1468), .B1(n1469), .B2(n1771), .C1(n1772), 
        .C2(n1472), .ZN(n1753) );
  AND4_X1 U3124 ( .A1(n1773), .A2(n1774), .A3(n1775), .A4(n1776), .ZN(n5380)
         );
  NOR4_X1 U3125 ( .A1(n1777), .A2(n1778), .A3(n1779), .A4(n1780), .ZN(n1776)
         );
  NAND3_X1 U3126 ( .A1(n5773), .A2(n5772), .A3(n5774), .ZN(n1780) );
  OAI211_X1 U3127 ( .C1(n5656), .C2(n5298), .A(n5770), .B(n5771), .ZN(n1779)
         );
  OAI222_X1 U3128 ( .A1(n5654), .A2(n5170), .B1(n5655), .B2(n5138), .C1(n5657), 
        .C2(n5266), .ZN(n1778) );
  OAI221_X1 U3129 ( .B1(n6925), .B2(n5074), .C1(n6353), .C2(n5106), .A(n1781), 
        .ZN(n1777) );
  AOI22_X1 U3130 ( .A1(n1782), .A2(n1453), .B1(n1783), .B2(n1455), .ZN(n1781)
         );
  AOI211_X1 U3131 ( .C1(n1784), .C2(n1457), .A(n1785), .B(n1786), .ZN(n1775)
         );
  OAI22_X1 U3132 ( .A1(n5637), .A2(n4722), .B1(n5647), .B2(n4626), .ZN(n1786)
         );
  OAI222_X1 U3133 ( .A1(n5642), .A2(n4562), .B1(n5648), .B2(n4530), .C1(n6936), 
        .C2(n4594), .ZN(n1785) );
  AOI221_X1 U3134 ( .B1(n6349), .B2(n1787), .C1(n1462), .C2(n1788), .A(n1789), 
        .ZN(n1774) );
  OAI22_X1 U3135 ( .A1(n4370), .A2(n1465), .B1(n5202), .B2(n1466), .ZN(n1789)
         );
  AOI222_X1 U3137 ( .A1(n1790), .A2(n1468), .B1(n1469), .B2(n1791), .C1(n1792), 
        .C2(n1472), .ZN(n1773) );
  AND4_X1 U3138 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(n5377)
         );
  NOR4_X1 U3139 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796)
         );
  NAND3_X1 U3140 ( .A1(n5766), .A2(n5765), .A3(n5767), .ZN(n1800) );
  OAI211_X1 U3141 ( .C1(n5656), .C2(n5297), .A(n5763), .B(n5764), .ZN(n1799)
         );
  OAI222_X1 U3142 ( .A1(n5654), .A2(n5169), .B1(n5655), .B2(n5137), .C1(n5657), 
        .C2(n5265), .ZN(n1798) );
  OAI221_X1 U3143 ( .B1(n6925), .B2(n5073), .C1(n6353), .C2(n5105), .A(n1801), 
        .ZN(n1797) );
  AOI22_X1 U3144 ( .A1(n1802), .A2(n1453), .B1(n1803), .B2(n1455), .ZN(n1801)
         );
  AOI211_X1 U3145 ( .C1(n1804), .C2(n1457), .A(n1805), .B(n1806), .ZN(n1795)
         );
  OAI22_X1 U3146 ( .A1(n5637), .A2(n4721), .B1(n5647), .B2(n4625), .ZN(n1806)
         );
  OAI222_X1 U3147 ( .A1(n5642), .A2(n4561), .B1(n5648), .B2(n4529), .C1(n6936), 
        .C2(n4593), .ZN(n1805) );
  AOI221_X1 U3148 ( .B1(n6348), .B2(n1807), .C1(n1462), .C2(n1808), .A(n1809), 
        .ZN(n1794) );
  OAI22_X1 U3149 ( .A1(n4369), .A2(n1465), .B1(n5201), .B2(n1466), .ZN(n1809)
         );
  AOI222_X1 U3151 ( .A1(n1810), .A2(n1468), .B1(n1469), .B2(n1811), .C1(n1812), 
        .C2(n1472), .ZN(n1793) );
  AND4_X1 U3152 ( .A1(n1813), .A2(n1814), .A3(n1815), .A4(n1816), .ZN(n5374)
         );
  NOR4_X1 U3153 ( .A1(n1817), .A2(n1818), .A3(n1819), .A4(n1820), .ZN(n1816)
         );
  NAND3_X1 U3154 ( .A1(n5758), .A2(n5757), .A3(n5759), .ZN(n1820) );
  OAI211_X1 U3155 ( .C1(n5656), .C2(n5296), .A(n5755), .B(n5756), .ZN(n1819)
         );
  OAI222_X1 U3156 ( .A1(n5654), .A2(n5168), .B1(n5655), .B2(n5136), .C1(n5657), 
        .C2(n5264), .ZN(n1818) );
  OAI221_X1 U3157 ( .B1(n6925), .B2(n5072), .C1(n6352), .C2(n5104), .A(n1821), 
        .ZN(n1817) );
  AOI22_X1 U3158 ( .A1(n1822), .A2(n1453), .B1(n1823), .B2(n1455), .ZN(n1821)
         );
  AOI211_X1 U3159 ( .C1(n1824), .C2(n1457), .A(n1825), .B(n1826), .ZN(n1815)
         );
  OAI22_X1 U3160 ( .A1(n5637), .A2(n4720), .B1(n5647), .B2(n4624), .ZN(n1826)
         );
  OAI222_X1 U3161 ( .A1(n5642), .A2(n4560), .B1(n5648), .B2(n4528), .C1(n6936), 
        .C2(n4592), .ZN(n1825) );
  AOI221_X1 U3162 ( .B1(n6349), .B2(n1827), .C1(n1462), .C2(n1828), .A(n1829), 
        .ZN(n1814) );
  OAI22_X1 U3163 ( .A1(n4368), .A2(n1465), .B1(n5200), .B2(n1466), .ZN(n1829)
         );
  AOI222_X1 U3165 ( .A1(n1830), .A2(n1468), .B1(n1469), .B2(n1831), .C1(n1832), 
        .C2(n1472), .ZN(n1813) );
  AND4_X1 U3166 ( .A1(n1833), .A2(n1834), .A3(n1835), .A4(n1836), .ZN(n5371)
         );
  NOR4_X1 U3167 ( .A1(n1837), .A2(n1838), .A3(n1839), .A4(n1840), .ZN(n1836)
         );
  NAND3_X1 U3168 ( .A1(n5749), .A2(n5748), .A3(n5750), .ZN(n1840) );
  OAI211_X1 U3169 ( .C1(n5656), .C2(n5295), .A(n5746), .B(n5747), .ZN(n1839)
         );
  OAI222_X1 U3170 ( .A1(n5654), .A2(n5167), .B1(n5655), .B2(n5135), .C1(n5657), 
        .C2(n5263), .ZN(n1838) );
  OAI221_X1 U3171 ( .B1(n6925), .B2(n5071), .C1(n6353), .C2(n5103), .A(n1841), 
        .ZN(n1837) );
  AOI22_X1 U3172 ( .A1(n1842), .A2(n1453), .B1(n1843), .B2(n1455), .ZN(n1841)
         );
  AOI211_X1 U3173 ( .C1(n1844), .C2(n1457), .A(n1845), .B(n1846), .ZN(n1835)
         );
  OAI22_X1 U3174 ( .A1(n5637), .A2(n4719), .B1(n5647), .B2(n4623), .ZN(n1846)
         );
  OAI222_X1 U3175 ( .A1(n5642), .A2(n4559), .B1(n5648), .B2(n4527), .C1(n6936), 
        .C2(n4591), .ZN(n1845) );
  AOI221_X1 U3176 ( .B1(n6349), .B2(n1847), .C1(n1462), .C2(n1848), .A(n1849), 
        .ZN(n1834) );
  OAI22_X1 U3177 ( .A1(n4367), .A2(n1465), .B1(n5199), .B2(n1466), .ZN(n1849)
         );
  AOI222_X1 U3179 ( .A1(n1850), .A2(n1468), .B1(n1469), .B2(n1851), .C1(n1852), 
        .C2(n1472), .ZN(n1833) );
  AND4_X1 U3180 ( .A1(n1853), .A2(n1854), .A3(n1855), .A4(n1856), .ZN(n5368)
         );
  NOR4_X1 U3181 ( .A1(n1857), .A2(n1858), .A3(n1859), .A4(n1860), .ZN(n1856)
         );
  NAND3_X1 U3182 ( .A1(n5744), .A2(n5743), .A3(n5745), .ZN(n1860) );
  OAI211_X1 U3183 ( .C1(n5656), .C2(n5294), .A(n5741), .B(n5742), .ZN(n1859)
         );
  OAI222_X1 U3184 ( .A1(n5654), .A2(n5166), .B1(n5655), .B2(n5134), .C1(n5657), 
        .C2(n5262), .ZN(n1858) );
  OAI221_X1 U3185 ( .B1(n6925), .B2(n5070), .C1(n6353), .C2(n5102), .A(n1861), 
        .ZN(n1857) );
  AOI22_X1 U3186 ( .A1(n1862), .A2(n1453), .B1(n1863), .B2(n1455), .ZN(n1861)
         );
  AOI211_X1 U3187 ( .C1(n1864), .C2(n1457), .A(n1865), .B(n1866), .ZN(n1855)
         );
  OAI22_X1 U3188 ( .A1(n5637), .A2(n4718), .B1(n5647), .B2(n4622), .ZN(n1866)
         );
  OAI222_X1 U3189 ( .A1(n5642), .A2(n4558), .B1(n5648), .B2(n4526), .C1(n6936), 
        .C2(n4590), .ZN(n1865) );
  AOI221_X1 U3190 ( .B1(n6349), .B2(n1867), .C1(n1462), .C2(n1868), .A(n1869), 
        .ZN(n1854) );
  OAI22_X1 U3191 ( .A1(n4366), .A2(n1465), .B1(n5198), .B2(n1466), .ZN(n1869)
         );
  AOI222_X1 U3193 ( .A1(n1870), .A2(n1468), .B1(n1469), .B2(n1871), .C1(n1872), 
        .C2(n1472), .ZN(n1853) );
  NOR4_X1 U3195 ( .A1(n1877), .A2(n1878), .A3(n1879), .A4(n1880), .ZN(n1876)
         );
  NAND3_X1 U3196 ( .A1(n5739), .A2(n5738), .A3(n5740), .ZN(n1880) );
  OAI211_X1 U3197 ( .C1(n5656), .C2(n5293), .A(n5736), .B(n5737), .ZN(n1879)
         );
  OAI222_X1 U3198 ( .A1(n5654), .A2(n5165), .B1(n5655), .B2(n5133), .C1(n5657), 
        .C2(n5261), .ZN(n1878) );
  OAI221_X1 U3199 ( .B1(n6925), .B2(n5069), .C1(n6352), .C2(n5101), .A(n1881), 
        .ZN(n1877) );
  AOI22_X1 U3200 ( .A1(n1882), .A2(n1453), .B1(n1883), .B2(n1455), .ZN(n1881)
         );
  AOI211_X1 U3201 ( .C1(n1884), .C2(n1457), .A(n1885), .B(n1886), .ZN(n1875)
         );
  OAI22_X1 U3202 ( .A1(n5637), .A2(n4717), .B1(n5647), .B2(n4621), .ZN(n1886)
         );
  OAI222_X1 U3203 ( .A1(n5642), .A2(n4557), .B1(n5648), .B2(n4525), .C1(n6936), 
        .C2(n4589), .ZN(n1885) );
  AOI221_X1 U3204 ( .B1(n6348), .B2(n1887), .C1(n1462), .C2(n1888), .A(n1889), 
        .ZN(n1874) );
  OAI22_X1 U3205 ( .A1(n4365), .A2(n1465), .B1(n5197), .B2(n1466), .ZN(n1889)
         );
  AOI222_X1 U3207 ( .A1(n1890), .A2(n1468), .B1(n1469), .B2(n1891), .C1(n1892), 
        .C2(n1472), .ZN(n1873) );
  AND4_X1 U3208 ( .A1(n1893), .A2(n1894), .A3(n1895), .A4(n1896), .ZN(n5362)
         );
  NOR4_X1 U3209 ( .A1(n1897), .A2(n1898), .A3(n1899), .A4(n1900), .ZN(n1896)
         );
  NAND3_X1 U3210 ( .A1(n5734), .A2(n5733), .A3(n5735), .ZN(n1900) );
  OAI211_X1 U3211 ( .C1(n5656), .C2(n5292), .A(n5731), .B(n5732), .ZN(n1899)
         );
  OAI222_X1 U3212 ( .A1(n5654), .A2(n5164), .B1(n5655), .B2(n5132), .C1(n5657), 
        .C2(n5260), .ZN(n1898) );
  OAI221_X1 U3213 ( .B1(n6925), .B2(n5068), .C1(n6353), .C2(n5100), .A(n1901), 
        .ZN(n1897) );
  AOI22_X1 U3214 ( .A1(n1902), .A2(n1453), .B1(n1903), .B2(n1455), .ZN(n1901)
         );
  AOI211_X1 U3215 ( .C1(n1904), .C2(n1457), .A(n1905), .B(n1906), .ZN(n1895)
         );
  OAI22_X1 U3216 ( .A1(n5637), .A2(n4716), .B1(n5647), .B2(n4620), .ZN(n1906)
         );
  OAI222_X1 U3217 ( .A1(n5642), .A2(n4556), .B1(n5648), .B2(n4524), .C1(n6936), 
        .C2(n4588), .ZN(n1905) );
  AOI221_X1 U3218 ( .B1(n6349), .B2(n1907), .C1(n1462), .C2(n1908), .A(n1909), 
        .ZN(n1894) );
  OAI22_X1 U3219 ( .A1(n4364), .A2(n1465), .B1(n5196), .B2(n1466), .ZN(n1909)
         );
  AOI222_X1 U3221 ( .A1(n1910), .A2(n1468), .B1(n1469), .B2(n1911), .C1(n1912), 
        .C2(n1472), .ZN(n1893) );
  NOR4_X1 U3223 ( .A1(n1917), .A2(n1918), .A3(n1919), .A4(n1920), .ZN(n1916)
         );
  NAND3_X1 U3224 ( .A1(n5724), .A2(n5723), .A3(n5725), .ZN(n1920) );
  OAI211_X1 U3225 ( .C1(n5656), .C2(n5291), .A(n5721), .B(n5722), .ZN(n1919)
         );
  OAI222_X1 U3226 ( .A1(n5654), .A2(n5163), .B1(n5655), .B2(n5131), .C1(n5657), 
        .C2(n5259), .ZN(n1918) );
  OAI221_X1 U3227 ( .B1(n6924), .B2(n5067), .C1(n6353), .C2(n5099), .A(n1921), 
        .ZN(n1917) );
  AOI22_X1 U3228 ( .A1(n1922), .A2(n1453), .B1(n1923), .B2(n1455), .ZN(n1921)
         );
  AOI211_X1 U3229 ( .C1(n1924), .C2(n1457), .A(n1925), .B(n1926), .ZN(n1915)
         );
  OAI22_X1 U3230 ( .A1(n5637), .A2(n4715), .B1(n5647), .B2(n4619), .ZN(n1926)
         );
  OAI222_X1 U3231 ( .A1(n5642), .A2(n4555), .B1(n5648), .B2(n4523), .C1(n6935), 
        .C2(n4587), .ZN(n1925) );
  AOI221_X1 U3232 ( .B1(n6349), .B2(n1927), .C1(n1462), .C2(n1928), .A(n1929), 
        .ZN(n1914) );
  OAI22_X1 U3233 ( .A1(n4363), .A2(n1465), .B1(n5195), .B2(n1466), .ZN(n1929)
         );
  AOI222_X1 U3235 ( .A1(n1930), .A2(n1468), .B1(n1469), .B2(n1931), .C1(n1932), 
        .C2(n1472), .ZN(n1913) );
  NOR4_X1 U3237 ( .A1(n1937), .A2(n1938), .A3(n1939), .A4(n1940), .ZN(n1936)
         );
  NAND3_X1 U3238 ( .A1(n5718), .A2(n5717), .A3(n5719), .ZN(n1940) );
  OAI211_X1 U3239 ( .C1(n5656), .C2(n5290), .A(n5715), .B(n5716), .ZN(n1939)
         );
  OAI222_X1 U3240 ( .A1(n5654), .A2(n5162), .B1(n5655), .B2(n5130), .C1(n5657), 
        .C2(n5258), .ZN(n1938) );
  OAI221_X1 U3241 ( .B1(n6925), .B2(n5066), .C1(n6352), .C2(n5098), .A(n1941), 
        .ZN(n1937) );
  AOI22_X1 U3242 ( .A1(n1942), .A2(n1453), .B1(n1943), .B2(n1455), .ZN(n1941)
         );
  AOI211_X1 U3243 ( .C1(n1944), .C2(n1457), .A(n1945), .B(n1946), .ZN(n1935)
         );
  OAI22_X1 U3244 ( .A1(n5637), .A2(n4714), .B1(n5647), .B2(n4618), .ZN(n1946)
         );
  OAI222_X1 U3245 ( .A1(n5642), .A2(n4554), .B1(n5648), .B2(n4522), .C1(n6936), 
        .C2(n4586), .ZN(n1945) );
  AOI221_X1 U3246 ( .B1(n6348), .B2(n1947), .C1(n1462), .C2(n1948), .A(n1949), 
        .ZN(n1934) );
  OAI22_X1 U3247 ( .A1(n4362), .A2(n1465), .B1(n5194), .B2(n1466), .ZN(n1949)
         );
  AOI222_X1 U3249 ( .A1(n1950), .A2(n1468), .B1(n1469), .B2(n1951), .C1(n1952), 
        .C2(n1472), .ZN(n1933) );
  AND4_X1 U3250 ( .A1(n1953), .A2(n1954), .A3(n1955), .A4(n1956), .ZN(n5353)
         );
  NOR4_X1 U3251 ( .A1(n1957), .A2(n1958), .A3(n1959), .A4(n1960), .ZN(n1956)
         );
  NAND3_X1 U3252 ( .A1(n5713), .A2(n5712), .A3(n5714), .ZN(n1960) );
  OAI211_X1 U3253 ( .C1(n5656), .C2(n5289), .A(n5710), .B(n5711), .ZN(n1959)
         );
  OAI222_X1 U3254 ( .A1(n5654), .A2(n5161), .B1(n5655), .B2(n5129), .C1(n5657), 
        .C2(n5257), .ZN(n1958) );
  OAI221_X1 U3255 ( .B1(n6925), .B2(n5065), .C1(n6352), .C2(n5097), .A(n1961), 
        .ZN(n1957) );
  AOI22_X1 U3256 ( .A1(n1962), .A2(n1453), .B1(n1963), .B2(n1455), .ZN(n1961)
         );
  AOI211_X1 U3257 ( .C1(n1964), .C2(n1457), .A(n1965), .B(n1966), .ZN(n1955)
         );
  OAI22_X1 U3258 ( .A1(n5637), .A2(n4713), .B1(n5647), .B2(n4617), .ZN(n1966)
         );
  OAI222_X1 U3259 ( .A1(n5642), .A2(n4553), .B1(n5648), .B2(n4521), .C1(n6936), 
        .C2(n4585), .ZN(n1965) );
  AOI221_X1 U3260 ( .B1(n6348), .B2(n1967), .C1(n1462), .C2(n1968), .A(n1969), 
        .ZN(n1954) );
  OAI22_X1 U3261 ( .A1(n4361), .A2(n1465), .B1(n5193), .B2(n1466), .ZN(n1969)
         );
  AOI222_X1 U3263 ( .A1(n1970), .A2(n1468), .B1(n1469), .B2(n1971), .C1(n1972), 
        .C2(n1472), .ZN(n1953) );
  AND4_X1 U3264 ( .A1(n1973), .A2(n1974), .A3(n1975), .A4(n1976), .ZN(n5350)
         );
  NOR4_X1 U3265 ( .A1(n1977), .A2(n1978), .A3(n1979), .A4(n1980), .ZN(n1976)
         );
  NAND3_X1 U3266 ( .A1(n5703), .A2(n5702), .A3(n5704), .ZN(n1980) );
  OAI211_X1 U3267 ( .C1(n5656), .C2(n5288), .A(n5700), .B(n5701), .ZN(n1979)
         );
  OAI222_X1 U3268 ( .A1(n5654), .A2(n5160), .B1(n5655), .B2(n5128), .C1(n5657), 
        .C2(n5256), .ZN(n1978) );
  OAI221_X1 U3269 ( .B1(n6925), .B2(n5064), .C1(n6352), .C2(n5096), .A(n1981), 
        .ZN(n1977) );
  AOI22_X1 U3270 ( .A1(n1982), .A2(n1453), .B1(n1983), .B2(n1455), .ZN(n1981)
         );
  AOI211_X1 U3271 ( .C1(n1984), .C2(n1457), .A(n1985), .B(n1986), .ZN(n1975)
         );
  OAI22_X1 U3272 ( .A1(n5637), .A2(n4712), .B1(n5647), .B2(n4616), .ZN(n1986)
         );
  OAI222_X1 U3273 ( .A1(n5642), .A2(n4552), .B1(n5648), .B2(n4520), .C1(n6936), 
        .C2(n4584), .ZN(n1985) );
  AOI221_X1 U3274 ( .B1(n6348), .B2(n1987), .C1(n1462), .C2(n1988), .A(n1989), 
        .ZN(n1974) );
  OAI22_X1 U3275 ( .A1(n4360), .A2(n1465), .B1(n5192), .B2(n1466), .ZN(n1989)
         );
  AOI222_X1 U3277 ( .A1(n1990), .A2(n1468), .B1(n1469), .B2(n1991), .C1(n1992), 
        .C2(n1472), .ZN(n1973) );
  AND4_X1 U3278 ( .A1(n1993), .A2(n1994), .A3(n1995), .A4(n1996), .ZN(n5347)
         );
  NOR4_X1 U3279 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(n1996)
         );
  NAND3_X1 U3280 ( .A1(n5693), .A2(n5692), .A3(n5694), .ZN(n2000) );
  OAI211_X1 U3281 ( .C1(n5656), .C2(n5287), .A(n5690), .B(n5691), .ZN(n1999)
         );
  OAI222_X1 U3282 ( .A1(n5654), .A2(n5159), .B1(n5655), .B2(n5127), .C1(n5657), 
        .C2(n5255), .ZN(n1998) );
  OAI221_X1 U3283 ( .B1(n6925), .B2(n5063), .C1(n6352), .C2(n5095), .A(n2001), 
        .ZN(n1997) );
  AOI22_X1 U3284 ( .A1(n2002), .A2(n1453), .B1(n2003), .B2(n1455), .ZN(n2001)
         );
  AOI211_X1 U3285 ( .C1(n2004), .C2(n1457), .A(n2005), .B(n2006), .ZN(n1995)
         );
  OAI22_X1 U3286 ( .A1(n5637), .A2(n4711), .B1(n5647), .B2(n4615), .ZN(n2006)
         );
  OAI222_X1 U3287 ( .A1(n5642), .A2(n4551), .B1(n5648), .B2(n4519), .C1(n6936), 
        .C2(n4583), .ZN(n2005) );
  AOI221_X1 U3288 ( .B1(n6348), .B2(n2007), .C1(n1462), .C2(n2008), .A(n2009), 
        .ZN(n1994) );
  OAI22_X1 U3289 ( .A1(n4359), .A2(n1465), .B1(n5191), .B2(n1466), .ZN(n2009)
         );
  AOI222_X1 U3291 ( .A1(n2010), .A2(n1468), .B1(n1469), .B2(n2011), .C1(n2012), 
        .C2(n1472), .ZN(n1993) );
  AND4_X1 U3292 ( .A1(n2013), .A2(n2014), .A3(n2015), .A4(n2016), .ZN(n5344)
         );
  NOR4_X1 U3293 ( .A1(n2017), .A2(n2018), .A3(n2019), .A4(n2020), .ZN(n2016)
         );
  NAND3_X1 U3294 ( .A1(n5683), .A2(n5682), .A3(n5684), .ZN(n2020) );
  OAI211_X1 U3295 ( .C1(n5656), .C2(n5286), .A(n5680), .B(n5681), .ZN(n2019)
         );
  OAI222_X1 U3296 ( .A1(n5654), .A2(n5158), .B1(n5655), .B2(n5126), .C1(n5657), 
        .C2(n5254), .ZN(n2018) );
  OAI221_X1 U3297 ( .B1(n6925), .B2(n5062), .C1(n6352), .C2(n5094), .A(n2021), 
        .ZN(n2017) );
  AOI22_X1 U3298 ( .A1(n2022), .A2(n1453), .B1(n2023), .B2(n1455), .ZN(n2021)
         );
  AOI211_X1 U3299 ( .C1(n2024), .C2(n1457), .A(n2025), .B(n2026), .ZN(n2015)
         );
  OAI22_X1 U3300 ( .A1(n5637), .A2(n4710), .B1(n5647), .B2(n4614), .ZN(n2026)
         );
  OAI222_X1 U3301 ( .A1(n5642), .A2(n4550), .B1(n5648), .B2(n4518), .C1(n6936), 
        .C2(n4582), .ZN(n2025) );
  AOI221_X1 U3302 ( .B1(n6349), .B2(n2027), .C1(n1462), .C2(n2028), .A(n2029), 
        .ZN(n2014) );
  OAI22_X1 U3303 ( .A1(n4358), .A2(n1465), .B1(n5190), .B2(n1466), .ZN(n2029)
         );
  AOI222_X1 U3305 ( .A1(n2030), .A2(n1468), .B1(n1469), .B2(n2031), .C1(n2032), 
        .C2(n1472), .ZN(n2013) );
  AND4_X1 U3306 ( .A1(n2033), .A2(n2034), .A3(n2035), .A4(n2036), .ZN(n5341)
         );
  NOR4_X1 U3307 ( .A1(n2037), .A2(n2038), .A3(n2039), .A4(n2040), .ZN(n2036)
         );
  NAND3_X1 U3308 ( .A1(n5673), .A2(n5672), .A3(n5674), .ZN(n2040) );
  OAI211_X1 U3309 ( .C1(n5656), .C2(n5285), .A(n5670), .B(n5671), .ZN(n2039)
         );
  OAI222_X1 U3310 ( .A1(n5654), .A2(n5157), .B1(n5655), .B2(n5125), .C1(n5657), 
        .C2(n5253), .ZN(n2038) );
  OAI221_X1 U3311 ( .B1(n6925), .B2(n5061), .C1(n6353), .C2(n5093), .A(n2041), 
        .ZN(n2037) );
  AOI22_X1 U3312 ( .A1(n2042), .A2(n1453), .B1(n2043), .B2(n1455), .ZN(n2041)
         );
  AOI211_X1 U3313 ( .C1(n2044), .C2(n1457), .A(n2045), .B(n2046), .ZN(n2035)
         );
  OAI22_X1 U3314 ( .A1(n5637), .A2(n4709), .B1(n5647), .B2(n4613), .ZN(n2046)
         );
  OAI222_X1 U3315 ( .A1(n5642), .A2(n4549), .B1(n5648), .B2(n4517), .C1(n6936), 
        .C2(n4581), .ZN(n2045) );
  AOI221_X1 U3316 ( .B1(n6349), .B2(n2047), .C1(n1462), .C2(n2048), .A(n2049), 
        .ZN(n2034) );
  OAI22_X1 U3317 ( .A1(n4357), .A2(n1465), .B1(n5189), .B2(n1466), .ZN(n2049)
         );
  AOI222_X1 U3319 ( .A1(n2050), .A2(n1468), .B1(n1469), .B2(n2051), .C1(n2052), 
        .C2(n1472), .ZN(n2033) );
  AND4_X1 U3320 ( .A1(n2053), .A2(n2054), .A3(n2055), .A4(n2056), .ZN(n5338)
         );
  NOR4_X1 U3321 ( .A1(n2057), .A2(n2058), .A3(n2059), .A4(n2060), .ZN(n2056)
         );
  NAND3_X1 U3322 ( .A1(n5661), .A2(n5660), .A3(n5662), .ZN(n2060) );
  OAI211_X1 U3323 ( .C1(n5656), .C2(n5284), .A(n5658), .B(n5659), .ZN(n2059)
         );
  OAI222_X1 U3324 ( .A1(n5654), .A2(n5156), .B1(n5655), .B2(n5124), .C1(n5657), 
        .C2(n5252), .ZN(n2058) );
  OAI221_X1 U3325 ( .B1(n6925), .B2(n5060), .C1(n6353), .C2(n5092), .A(n2061), 
        .ZN(n2057) );
  AOI22_X1 U3326 ( .A1(n2062), .A2(n1453), .B1(n2063), .B2(n1455), .ZN(n2061)
         );
  AOI211_X1 U3327 ( .C1(n2064), .C2(n1457), .A(n2065), .B(n2066), .ZN(n2055)
         );
  OAI22_X1 U3328 ( .A1(n5637), .A2(n4708), .B1(n5647), .B2(n4612), .ZN(n2066)
         );
  OAI222_X1 U3329 ( .A1(n5642), .A2(n4548), .B1(n5648), .B2(n4516), .C1(n6936), 
        .C2(n4580), .ZN(n2065) );
  AOI221_X1 U3330 ( .B1(n6349), .B2(n2067), .C1(n1462), .C2(n2068), .A(n2069), 
        .ZN(n2054) );
  OAI22_X1 U3331 ( .A1(n4356), .A2(n1465), .B1(n5188), .B2(n1466), .ZN(n2069)
         );
  AOI222_X1 U3333 ( .A1(n2070), .A2(n1468), .B1(n1469), .B2(n2071), .C1(n2072), 
        .C2(n1472), .ZN(n2053) );
  AND4_X1 U3334 ( .A1(n2073), .A2(n2074), .A3(n2075), .A4(n2076), .ZN(n5333)
         );
  NOR4_X1 U3335 ( .A1(n2077), .A2(n2078), .A3(n2079), .A4(n2080), .ZN(n2076)
         );
  NAND3_X1 U3336 ( .A1(n5644), .A2(n5639), .A3(n5651), .ZN(n2080) );
  OAI211_X1 U3337 ( .C1(n5656), .C2(n5283), .A(n5629), .B(n5634), .ZN(n2079)
         );
  OAI222_X1 U3338 ( .A1(n5654), .A2(n5155), .B1(n5655), .B2(n5123), .C1(n5657), 
        .C2(n5251), .ZN(n2078) );
  OAI221_X1 U3339 ( .B1(n6925), .B2(n5059), .C1(n6352), .C2(n5091), .A(n2081), 
        .ZN(n2077) );
  AOI22_X1 U3340 ( .A1(n2082), .A2(n1453), .B1(n2083), .B2(n1455), .ZN(n2081)
         );
  AOI211_X1 U3343 ( .C1(n2084), .C2(n1457), .A(n2085), .B(n2086), .ZN(n2075)
         );
  OAI22_X1 U3344 ( .A1(n5637), .A2(n4707), .B1(n5647), .B2(n4611), .ZN(n2086)
         );
  OAI222_X1 U3345 ( .A1(n5642), .A2(n4547), .B1(n5648), .B2(n4515), .C1(n6936), 
        .C2(n4579), .ZN(n2085) );
  AOI221_X1 U3347 ( .B1(n6348), .B2(n2087), .C1(n1462), .C2(n2088), .A(n2089), 
        .ZN(n2074) );
  OAI22_X1 U3348 ( .A1(n4355), .A2(n1465), .B1(n5187), .B2(n1466), .ZN(n2089)
         );
  INV_X1 U3352 ( .A(n5892), .ZN(n2090) );
  AOI222_X1 U3355 ( .A1(n2091), .A2(n1468), .B1(n1469), .B2(n2092), .C1(n2093), 
        .C2(n1472), .ZN(n2073) );
  AND4_X1 U3360 ( .A1(n2094), .A2(n2095), .A3(n2096), .A4(n2097), .ZN(n5324)
         );
  NOR4_X1 U3361 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(n2097)
         );
  NAND3_X1 U3362 ( .A1(n5520), .A2(n5519), .A3(n5521), .ZN(n2101) );
  OAI211_X1 U3363 ( .C1(n5462), .C2(n5314), .A(n5517), .B(n5518), .ZN(n2100)
         );
  OAI222_X1 U3364 ( .A1(n5460), .A2(n5186), .B1(n5461), .B2(n5154), .C1(n5463), 
        .C2(n5282), .ZN(n2099) );
  OAI221_X1 U3365 ( .B1(n5433), .B2(n5090), .C1(n5434), .C2(n5122), .A(n2102), 
        .ZN(n2098) );
  AOI22_X1 U3366 ( .A1(n1452), .A2(n2103), .B1(n1454), .B2(n2104), .ZN(n2102)
         );
  AOI211_X1 U3369 ( .C1(n1456), .C2(n2105), .A(n2106), .B(n2107), .ZN(n2096)
         );
  OAI22_X1 U3370 ( .A1(n5443), .A2(n4738), .B1(n5453), .B2(n4642), .ZN(n2107)
         );
  OAI222_X1 U3371 ( .A1(n5448), .A2(n4578), .B1(n5454), .B2(n4546), .C1(n5449), 
        .C2(n4610), .ZN(n2106) );
  AOI221_X1 U3373 ( .B1(n2108), .B2(n1463), .C1(n2109), .C2(n2110), .A(n2111), 
        .ZN(n2095) );
  OAI22_X1 U3374 ( .A1(n4386), .A2(n6901), .B1(n4994), .B2(n2113), .ZN(n2111)
         );
  AOI222_X1 U3377 ( .A1(n1467), .A2(n2114), .B1(n2115), .B2(n1470), .C1(n1471), 
        .C2(n2116), .ZN(n2094) );
  AND4_X1 U3381 ( .A1(n2117), .A2(n2118), .A3(n2119), .A4(n2120), .ZN(n5323)
         );
  NOR4_X1 U3382 ( .A1(n2121), .A2(n2122), .A3(n2123), .A4(n2124), .ZN(n2120)
         );
  NAND3_X1 U3383 ( .A1(n5512), .A2(n5511), .A3(n5513), .ZN(n2124) );
  OAI211_X1 U3384 ( .C1(n5462), .C2(n5298), .A(n5509), .B(n5510), .ZN(n2123)
         );
  OAI222_X1 U3385 ( .A1(n5460), .A2(n5170), .B1(n5461), .B2(n5138), .C1(n5463), 
        .C2(n5266), .ZN(n2122) );
  OAI221_X1 U3386 ( .B1(n5433), .B2(n5074), .C1(n5434), .C2(n5106), .A(n2125), 
        .ZN(n2121) );
  AOI22_X1 U3387 ( .A1(n1782), .A2(n2103), .B1(n1783), .B2(n2104), .ZN(n2125)
         );
  AOI211_X1 U3390 ( .C1(n1784), .C2(n2105), .A(n2126), .B(n2127), .ZN(n2119)
         );
  OAI22_X1 U3391 ( .A1(n5443), .A2(n4722), .B1(n5453), .B2(n4626), .ZN(n2127)
         );
  OAI222_X1 U3392 ( .A1(n5448), .A2(n4562), .B1(n5454), .B2(n4530), .C1(n5449), 
        .C2(n4594), .ZN(n2126) );
  AOI221_X1 U3394 ( .B1(n2108), .B2(n1788), .C1(n2109), .C2(n2128), .A(n2129), 
        .ZN(n2118) );
  OAI22_X1 U3395 ( .A1(n4370), .A2(n6901), .B1(n4978), .B2(n2113), .ZN(n2129)
         );
  AOI222_X1 U3398 ( .A1(n1790), .A2(n2114), .B1(n2115), .B2(n1791), .C1(n1792), 
        .C2(n2116), .ZN(n2117) );
  NOR4_X1 U3403 ( .A1(n2134), .A2(n2135), .A3(n2136), .A4(n2137), .ZN(n2133)
         );
  NAND3_X1 U3404 ( .A1(n5504), .A2(n5503), .A3(n5505), .ZN(n2137) );
  OAI211_X1 U3405 ( .C1(n5462), .C2(n5297), .A(n5501), .B(n5502), .ZN(n2136)
         );
  OAI222_X1 U3406 ( .A1(n5460), .A2(n5169), .B1(n5461), .B2(n5137), .C1(n5463), 
        .C2(n5265), .ZN(n2135) );
  OAI221_X1 U3407 ( .B1(n5433), .B2(n5073), .C1(n5434), .C2(n5105), .A(n2138), 
        .ZN(n2134) );
  AOI22_X1 U3408 ( .A1(n1802), .A2(n2103), .B1(n1803), .B2(n2104), .ZN(n2138)
         );
  AOI211_X1 U3411 ( .C1(n1804), .C2(n2105), .A(n2139), .B(n2140), .ZN(n2132)
         );
  OAI22_X1 U3412 ( .A1(n5443), .A2(n4721), .B1(n5453), .B2(n4625), .ZN(n2140)
         );
  OAI222_X1 U3413 ( .A1(n5448), .A2(n4561), .B1(n5454), .B2(n4529), .C1(n5449), 
        .C2(n4593), .ZN(n2139) );
  AOI221_X1 U3415 ( .B1(n2108), .B2(n1808), .C1(n2109), .C2(n2141), .A(n2142), 
        .ZN(n2131) );
  OAI22_X1 U3416 ( .A1(n4369), .A2(n6900), .B1(n4977), .B2(n2113), .ZN(n2142)
         );
  AOI222_X1 U3419 ( .A1(n1810), .A2(n2114), .B1(n2115), .B2(n1811), .C1(n1812), 
        .C2(n2116), .ZN(n2130) );
  AND4_X1 U3423 ( .A1(n2143), .A2(n2144), .A3(n2145), .A4(n2146), .ZN(n5321)
         );
  NOR4_X1 U3424 ( .A1(n2147), .A2(n2148), .A3(n2149), .A4(n2150), .ZN(n2146)
         );
  NAND3_X1 U3425 ( .A1(n5496), .A2(n5495), .A3(n5497), .ZN(n2150) );
  OAI211_X1 U3426 ( .C1(n5462), .C2(n5296), .A(n5493), .B(n5494), .ZN(n2149)
         );
  OAI222_X1 U3427 ( .A1(n5460), .A2(n5168), .B1(n5461), .B2(n5136), .C1(n5463), 
        .C2(n5264), .ZN(n2148) );
  OAI221_X1 U3428 ( .B1(n5433), .B2(n5072), .C1(n5434), .C2(n5104), .A(n2151), 
        .ZN(n2147) );
  AOI22_X1 U3429 ( .A1(n1822), .A2(n2103), .B1(n1823), .B2(n2104), .ZN(n2151)
         );
  AOI211_X1 U3432 ( .C1(n1824), .C2(n2105), .A(n2152), .B(n2153), .ZN(n2145)
         );
  OAI22_X1 U3433 ( .A1(n5443), .A2(n4720), .B1(n5453), .B2(n4624), .ZN(n2153)
         );
  OAI222_X1 U3434 ( .A1(n5448), .A2(n4560), .B1(n5454), .B2(n4528), .C1(n5449), 
        .C2(n4592), .ZN(n2152) );
  AOI221_X1 U3436 ( .B1(n2108), .B2(n1828), .C1(n2109), .C2(n2154), .A(n2155), 
        .ZN(n2144) );
  OAI22_X1 U3437 ( .A1(n4368), .A2(n6901), .B1(n4976), .B2(n2113), .ZN(n2155)
         );
  AOI222_X1 U3440 ( .A1(n1830), .A2(n2114), .B1(n2115), .B2(n1831), .C1(n1832), 
        .C2(n2116), .ZN(n2143) );
  NOR4_X1 U3445 ( .A1(n2160), .A2(n2161), .A3(n2162), .A4(n2163), .ZN(n2159)
         );
  NAND3_X1 U3446 ( .A1(n5488), .A2(n5487), .A3(n5489), .ZN(n2163) );
  OAI211_X1 U3447 ( .C1(n5462), .C2(n5295), .A(n5485), .B(n5486), .ZN(n2162)
         );
  OAI222_X1 U3448 ( .A1(n5460), .A2(n5167), .B1(n5461), .B2(n5135), .C1(n5463), 
        .C2(n5263), .ZN(n2161) );
  OAI221_X1 U3449 ( .B1(n5433), .B2(n5071), .C1(n5434), .C2(n5103), .A(n2164), 
        .ZN(n2160) );
  AOI22_X1 U3450 ( .A1(n1842), .A2(n2103), .B1(n1843), .B2(n2104), .ZN(n2164)
         );
  AOI211_X1 U3453 ( .C1(n1844), .C2(n2105), .A(n2165), .B(n2166), .ZN(n2158)
         );
  OAI22_X1 U3454 ( .A1(n5443), .A2(n4719), .B1(n5453), .B2(n4623), .ZN(n2166)
         );
  OAI222_X1 U3455 ( .A1(n5448), .A2(n4559), .B1(n5454), .B2(n4527), .C1(n5449), 
        .C2(n4591), .ZN(n2165) );
  AOI221_X1 U3457 ( .B1(n2108), .B2(n1848), .C1(n2109), .C2(n2167), .A(n2168), 
        .ZN(n2157) );
  OAI22_X1 U3458 ( .A1(n4367), .A2(n6902), .B1(n4975), .B2(n2113), .ZN(n2168)
         );
  AOI222_X1 U3461 ( .A1(n1850), .A2(n2114), .B1(n2115), .B2(n1851), .C1(n1852), 
        .C2(n2116), .ZN(n2156) );
  AND4_X1 U3465 ( .A1(n2169), .A2(n2170), .A3(n2171), .A4(n2172), .ZN(n5319)
         );
  NOR4_X1 U3466 ( .A1(n2173), .A2(n2174), .A3(n2175), .A4(n2176), .ZN(n2172)
         );
  NAND3_X1 U3467 ( .A1(n5480), .A2(n5479), .A3(n5481), .ZN(n2176) );
  OAI211_X1 U3468 ( .C1(n5462), .C2(n5294), .A(n5477), .B(n5478), .ZN(n2175)
         );
  OAI222_X1 U3469 ( .A1(n5460), .A2(n5166), .B1(n5461), .B2(n5134), .C1(n5463), 
        .C2(n5262), .ZN(n2174) );
  OAI221_X1 U3470 ( .B1(n5433), .B2(n5070), .C1(n5434), .C2(n5102), .A(n2177), 
        .ZN(n2173) );
  AOI22_X1 U3471 ( .A1(n1862), .A2(n2103), .B1(n1863), .B2(n2104), .ZN(n2177)
         );
  AOI211_X1 U3474 ( .C1(n1864), .C2(n2105), .A(n2178), .B(n2179), .ZN(n2171)
         );
  OAI22_X1 U3475 ( .A1(n5443), .A2(n4718), .B1(n5453), .B2(n4622), .ZN(n2179)
         );
  OAI222_X1 U3476 ( .A1(n5448), .A2(n4558), .B1(n5454), .B2(n4526), .C1(n5449), 
        .C2(n4590), .ZN(n2178) );
  AOI221_X1 U3478 ( .B1(n2108), .B2(n1868), .C1(n2109), .C2(n2180), .A(n2181), 
        .ZN(n2170) );
  OAI22_X1 U3479 ( .A1(n4366), .A2(n6900), .B1(n4974), .B2(n2113), .ZN(n2181)
         );
  AOI222_X1 U3482 ( .A1(n1870), .A2(n2114), .B1(n2115), .B2(n1871), .C1(n1872), 
        .C2(n2116), .ZN(n2169) );
  NOR4_X1 U3487 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2185)
         );
  NAND3_X1 U3488 ( .A1(n5472), .A2(n5471), .A3(n5473), .ZN(n2189) );
  OAI211_X1 U3489 ( .C1(n5462), .C2(n5293), .A(n5469), .B(n5470), .ZN(n2188)
         );
  OAI222_X1 U3490 ( .A1(n5460), .A2(n5165), .B1(n5461), .B2(n5133), .C1(n5463), 
        .C2(n5261), .ZN(n2187) );
  OAI221_X1 U3491 ( .B1(n5433), .B2(n5069), .C1(n5434), .C2(n5101), .A(n2190), 
        .ZN(n2186) );
  AOI22_X1 U3492 ( .A1(n1882), .A2(n2103), .B1(n1883), .B2(n2104), .ZN(n2190)
         );
  AOI211_X1 U3495 ( .C1(n1884), .C2(n2105), .A(n2191), .B(n2192), .ZN(n2184)
         );
  OAI22_X1 U3496 ( .A1(n5443), .A2(n4717), .B1(n5453), .B2(n4621), .ZN(n2192)
         );
  OAI222_X1 U3497 ( .A1(n5448), .A2(n4557), .B1(n5454), .B2(n4525), .C1(n5449), 
        .C2(n4589), .ZN(n2191) );
  AOI221_X1 U3499 ( .B1(n2108), .B2(n1888), .C1(n2109), .C2(n2193), .A(n2194), 
        .ZN(n2183) );
  OAI22_X1 U3500 ( .A1(n4365), .A2(n6901), .B1(n4973), .B2(n2113), .ZN(n2194)
         );
  AOI222_X1 U3503 ( .A1(n1890), .A2(n2114), .B1(n2115), .B2(n1891), .C1(n1892), 
        .C2(n2116), .ZN(n2182) );
  AND4_X1 U3507 ( .A1(n2195), .A2(n2196), .A3(n2197), .A4(n2198), .ZN(n5317)
         );
  NOR4_X1 U3508 ( .A1(n2199), .A2(n2200), .A3(n2201), .A4(n2202), .ZN(n2198)
         );
  NAND3_X1 U3509 ( .A1(n5450), .A2(n5445), .A3(n5457), .ZN(n2202) );
  OAI211_X1 U3510 ( .C1(n5462), .C2(n5291), .A(n5435), .B(n5440), .ZN(n2201)
         );
  OAI222_X1 U3511 ( .A1(n5460), .A2(n5163), .B1(n5461), .B2(n5131), .C1(n5463), 
        .C2(n5259), .ZN(n2200) );
  OAI221_X1 U3512 ( .B1(n5433), .B2(n5067), .C1(n5434), .C2(n5099), .A(n2203), 
        .ZN(n2199) );
  AOI22_X1 U3513 ( .A1(n1922), .A2(n2103), .B1(n1923), .B2(n2104), .ZN(n2203)
         );
  AOI211_X1 U3516 ( .C1(n1924), .C2(n2105), .A(n2204), .B(n2205), .ZN(n2197)
         );
  OAI22_X1 U3517 ( .A1(n5443), .A2(n4715), .B1(n5453), .B2(n4619), .ZN(n2205)
         );
  OAI222_X1 U3518 ( .A1(n5448), .A2(n4555), .B1(n5454), .B2(n4523), .C1(n5449), 
        .C2(n4587), .ZN(n2204) );
  AOI221_X1 U3520 ( .B1(n2108), .B2(n1928), .C1(n2109), .C2(n2206), .A(n2207), 
        .ZN(n2196) );
  OAI22_X1 U3521 ( .A1(n4363), .A2(n6900), .B1(n4971), .B2(n2113), .ZN(n2207)
         );
  AOI222_X1 U3524 ( .A1(n1930), .A2(n2114), .B1(n2115), .B2(n1931), .C1(n1932), 
        .C2(n2116), .ZN(n2195) );
  NAND3_X1 U3530 ( .A1(n6272), .A2(n6268), .A3(n6277), .ZN(n2215) );
  OAI211_X1 U3531 ( .C1(n5462), .C2(n5290), .A(n6257), .B(n6264), .ZN(n2214)
         );
  OAI222_X1 U3532 ( .A1(n5460), .A2(n5162), .B1(n5461), .B2(n5130), .C1(n5463), 
        .C2(n5258), .ZN(n2213) );
  OAI221_X1 U3533 ( .B1(n5433), .B2(n5066), .C1(n5434), .C2(n5098), .A(n2216), 
        .ZN(n2212) );
  AOI22_X1 U3534 ( .A1(n1942), .A2(n2103), .B1(n1943), .B2(n2104), .ZN(n2216)
         );
  AOI211_X1 U3537 ( .C1(n1944), .C2(n2105), .A(n2217), .B(n2218), .ZN(n2210)
         );
  OAI22_X1 U3538 ( .A1(n5443), .A2(n4714), .B1(n5453), .B2(n4618), .ZN(n2218)
         );
  OAI222_X1 U3539 ( .A1(n5448), .A2(n4554), .B1(n5454), .B2(n4522), .C1(n5449), 
        .C2(n4586), .ZN(n2217) );
  AOI221_X1 U3541 ( .B1(n2108), .B2(n1948), .C1(n2109), .C2(n2219), .A(n2220), 
        .ZN(n2209) );
  OAI22_X1 U3542 ( .A1(n4362), .A2(n6902), .B1(n4970), .B2(n2113), .ZN(n2220)
         );
  AOI222_X1 U3545 ( .A1(n1950), .A2(n2114), .B1(n2115), .B2(n1951), .C1(n1952), 
        .C2(n2116), .ZN(n2208) );
  NAND2_X1 U3549 ( .A1(n1012), .A2(n1095), .ZN(dmem_read) );
  NAND2_X1 U3551 ( .A1(n1012), .A2(n1090), .ZN(dmem_ishalf) );
  NAND2_X1 U3553 ( .A1(n1083), .A2(n1012), .ZN(dmem_isbyte) );
  INV_X1 U3554 ( .A(\UUT/x_we ), .ZN(n1012) );
  NOR2_X1 U3556 ( .A1(\UUT/regfile/N267 ), .A2(n2221), .ZN(\UUT/regfile/N269 )
         );
  INV_X1 U3557 ( .A(n5877), .ZN(n2221) );
  OAI211_X1 U3558 ( .C1(\UUT/Mpath/the_alu/N81 ), .C2(n7215), .A(n2222), .B(
        n2223), .ZN(\UUT/daddr_out [1]) );
  AOI22_X1 U3559 ( .A1(\UUT/Mpath/the_alu/diff[1] ), .A2(n1223), .B1(
        \UUT/Mpath/the_alu/sum[1] ), .B2(n7213), .ZN(n2223) );
  AOI22_X1 U3560 ( .A1(\UUT/Mpath/the_alu/N82 ), .A2(n2224), .B1(n2225), .B2(
        n2226), .ZN(n2222) );
  INV_X1 U3561 ( .A(\UUT/Mpath/the_alu/N82 ), .ZN(n2226) );
  OAI221_X1 U3562 ( .B1(n2227), .B2(n1301), .C1(\UUT/Mpath/the_alu/N81 ), .C2(
        n1303), .A(n1304), .ZN(n2225) );
  NAND2_X1 U3563 ( .A1(n6323), .A2(\UUT/Mpath/the_alu/N492 ), .ZN(n1303) );
  OAI22_X1 U3564 ( .A1(\UUT/Mpath/the_alu/N81 ), .A2(n1301), .B1(n1305), .B2(
        n2227), .ZN(n2224) );
  INV_X1 U3565 ( .A(\UUT/Mpath/the_alu/N81 ), .ZN(n2227) );
  INV_X1 U3568 ( .A(\UUT/Mpath/the_alu/N486 ), .ZN(n2229) );
  INV_X1 U3572 ( .A(n6324), .ZN(n2230) );
  INV_X1 U3574 ( .A(n2228), .ZN(n2231) );
  NAND2_X1 U3576 ( .A1(n2232), .A2(n2233), .ZN(\UUT/daddr_out [0]) );
  AOI21_X1 U3577 ( .B1(\UUT/Mpath/the_alu/diff[0] ), .B2(n1223), .A(n2234), 
        .ZN(n2233) );
  NOR3_X1 U3578 ( .A1(n2235), .A2(n2236), .A3(n7213), .ZN(n2234) );
  AOI22_X1 U3579 ( .A1(n2237), .A2(\UUT/Mpath/the_alu/N93 ), .B1(
        \UUT/Mpath/the_alu/N91 ), .B2(n2238), .ZN(n2236) );
  AND2_X1 U3580 ( .A1(\UUT/Mpath/the_alu/N498 ), .A2(\UUT/Mpath/the_alu/N503 ), 
        .ZN(n2237) );
  INV_X1 U3582 ( .A(n2235), .ZN(n2239) );
  AOI22_X1 U3583 ( .A1(\UUT/Mpath/the_alu/sum[0] ), .A2(n7213), .B1(n6326), 
        .B2(n6323), .ZN(n2232) );
  INV_X1 U3585 ( .A(\UUT/Mpath/the_alu/N503 ), .ZN(n2238) );
  INV_X1 U3588 ( .A(\UUT/Mpath/the_alu/N468 ), .ZN(n2240) );
  INV_X1 U3589 ( .A(n1061), .ZN(\UUT/d_mul_command [5]) );
  NAND2_X1 U3590 ( .A1(n2241), .A2(\UUT/Mcontrol/d_sampled_finstr [5]), .ZN(
        n1061) );
  INV_X1 U3591 ( .A(n1053), .ZN(\UUT/d_mul_command [4]) );
  NAND2_X1 U3592 ( .A1(n2241), .A2(n7202), .ZN(n1053) );
  NAND2_X1 U3593 ( .A1(n2241), .A2(n5327), .ZN(\UUT/d_mul_command [3]) );
  NAND2_X1 U3594 ( .A1(n2241), .A2(n7210), .ZN(\UUT/d_mul_command [2]) );
  NAND2_X1 U3595 ( .A1(n2241), .A2(n5329), .ZN(\UUT/d_mul_command [1]) );
  NAND2_X1 U3596 ( .A1(n2241), .A2(n5330), .ZN(\UUT/d_mul_command [0]) );
  AND2_X1 U3597 ( .A1(n1039), .A2(\UUT/Mcontrol/Operation_decoding32/N2043 ), 
        .ZN(n2241) );
  INV_X1 U3598 ( .A(\UUT/Mcontrol/st_logic/N42 ), .ZN(\UUT/byp_controlB[0] )
         );
  INV_X1 U3599 ( .A(n84), .ZN(\UUT/break_code[23] ) );
  AOI221_X1 U3600 ( .B1(n5970), .B2(n2242), .C1(\UUT/Mcontrol/d_instr [7]), 
        .C2(n2243), .A(n2244), .ZN(n84) );
  INV_X1 U3601 ( .A(n294), .ZN(\UUT/break_code[22] ) );
  AOI221_X1 U3602 ( .B1(n5981), .B2(n2242), .C1(n2243), .C2(
        \UUT/Mcontrol/d_instr [6]), .A(n2244), .ZN(n294) );
  INV_X1 U3603 ( .A(n325), .ZN(\UUT/break_code[21] ) );
  INV_X1 U3605 ( .A(n348), .ZN(\UUT/break_code[20] ) );
  OAI21_X1 U3607 ( .B1(n947), .B2(n202), .A(n2245), .ZN(n2244) );
  NAND3_X1 U3608 ( .A1(\UUT/Mcontrol/d_sampled_finstr [15]), .A2(n6982), .A3(
        n451), .ZN(n202) );
  NOR2_X1 U3609 ( .A1(n946), .A2(n947), .ZN(n2242) );
  NAND2_X1 U3610 ( .A1(n6968), .A2(n451), .ZN(n946) );
  INV_X1 U3611 ( .A(n2246), .ZN(n6002) );
  NAND4_X1 U3612 ( .A1(n1097), .A2(\UUT/Mcontrol/Operation_decoding32/N1987 ), 
        .A3(n7101), .A4(n6875), .ZN(n2246) );
  OAI21_X1 U3615 ( .B1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .B2(n2247), 
        .A(n2248), .ZN(n1097) );
  NAND3_X1 U3616 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2005 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N2017 ), .ZN(n2248) );
  INV_X1 U3617 ( .A(\UUT/Mcontrol/Operation_decoding32/N1999 ), .ZN(n2247) );
  NAND2_X1 U3618 ( .A1(n2249), .A2(n2250), .ZN(\UUT/break_code[1] ) );
  NAND3_X1 U3619 ( .A1(n5960), .A2(n7098), .A3(\UUT/Mcontrol/d_instr [7]), 
        .ZN(n2250) );
  NAND2_X1 U3620 ( .A1(\UUT/Mcontrol/d_instr [1]), .A2(n2251), .ZN(n2249) );
  INV_X1 U3621 ( .A(n2252), .ZN(n2251) );
  INV_X1 U3624 ( .A(n6015), .ZN(n2254) );
  INV_X1 U3627 ( .A(n6027), .ZN(n2257) );
  OAI221_X1 U3628 ( .B1(n2253), .B2(n2258), .C1(n5329), .C2(n2255), .A(n2256), 
        .ZN(\UUT/break_code[17] ) );
  INV_X1 U3629 ( .A(\UUT/Mcontrol/d_sampled_finstr [1]), .ZN(n5329) );
  INV_X1 U3630 ( .A(n6048), .ZN(n2258) );
  OAI221_X1 U3631 ( .B1(n2253), .B2(n2259), .C1(n5330), .C2(n2255), .A(n2256), 
        .ZN(\UUT/break_code[16] ) );
  AOI21_X1 U3632 ( .B1(n5920), .B2(n6016), .A(n456), .ZN(n2256) );
  INV_X1 U3633 ( .A(n2245), .ZN(n456) );
  NAND2_X1 U3634 ( .A1(n482), .A2(n1119), .ZN(n2245) );
  INV_X1 U3635 ( .A(n1048), .ZN(n1119) );
  INV_X1 U3636 ( .A(n2243), .ZN(n2255) );
  NOR2_X1 U3637 ( .A1(n451), .A2(n947), .ZN(n2243) );
  INV_X1 U3638 ( .A(n7096), .ZN(n451) );
  INV_X1 U3639 ( .A(\UUT/Mcontrol/d_sampled_finstr [0]), .ZN(n5330) );
  INV_X1 U3640 ( .A(n6060), .ZN(n2259) );
  NAND2_X1 U3641 ( .A1(n5920), .A2(n6849), .ZN(n2253) );
  INV_X1 U3645 ( .A(n6871), .ZN(n1038) );
  INV_X1 U3647 ( .A(n475), .ZN(\UUT/break_code[15] ) );
  AOI22_X1 U3648 ( .A1(n6071), .A2(n482), .B1(n479), .B2(n480), .ZN(n475) );
  INV_X1 U3649 ( .A(n6074), .ZN(n479) );
  NOR2_X1 U3650 ( .A1(n1058), .A2(n5720), .ZN(n482) );
  OAI21_X1 U3652 ( .B1(n5902), .B2(n2260), .A(n2261), .ZN(\UUT/break_code[14] ) );
  NAND2_X1 U3653 ( .A1(n6085), .A2(n2262), .ZN(n2261) );
  OAI21_X1 U3655 ( .B1(n5903), .B2(n2260), .A(n2263), .ZN(\UUT/break_code[13] ) );
  NAND2_X1 U3656 ( .A1(n6095), .A2(n2262), .ZN(n2263) );
  NAND3_X1 U3659 ( .A1(n5960), .A2(n7098), .A3(\UUT/Mcontrol/d_instr [6]), 
        .ZN(n2264) );
  NOR2_X1 U3661 ( .A1(n7062), .A2(n1058), .ZN(n1056) );
  INV_X1 U3663 ( .A(n5966), .ZN(n5382) );
  NOR4_X1 U3665 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n2269)
         );
  NAND3_X1 U3666 ( .A1(n5964), .A2(n5963), .A3(n5965), .ZN(n2273) );
  OAI211_X1 U3667 ( .C1(n5462), .C2(n5299), .A(n5961), .B(n5962), .ZN(n2272)
         );
  OAI222_X1 U3668 ( .A1(n5460), .A2(n5171), .B1(n5461), .B2(n5139), .C1(n5463), 
        .C2(n5267), .ZN(n2271) );
  OAI221_X1 U3669 ( .B1(n5433), .B2(n5075), .C1(n5434), .C2(n5107), .A(n2274), 
        .ZN(n2270) );
  AOI22_X1 U3670 ( .A1(n1762), .A2(n2103), .B1(n1763), .B2(n2104), .ZN(n2274)
         );
  AOI211_X1 U3673 ( .C1(n1764), .C2(n2105), .A(n2275), .B(n2276), .ZN(n2268)
         );
  OAI22_X1 U3674 ( .A1(n5443), .A2(n4723), .B1(n5453), .B2(n4627), .ZN(n2276)
         );
  OAI222_X1 U3675 ( .A1(n5448), .A2(n4563), .B1(n5454), .B2(n4531), .C1(n5449), 
        .C2(n4595), .ZN(n2275) );
  AOI221_X1 U3677 ( .B1(n2108), .B2(n1768), .C1(n2109), .C2(n2277), .A(n2278), 
        .ZN(n2267) );
  OAI22_X1 U3678 ( .A1(n4371), .A2(n6901), .B1(n4979), .B2(n2113), .ZN(n2278)
         );
  AOI222_X1 U3681 ( .A1(n1770), .A2(n2114), .B1(n2115), .B2(n1771), .C1(n1772), 
        .C2(n2116), .ZN(n2266) );
  INV_X1 U3686 ( .A(n5977), .ZN(n5385) );
  NOR4_X1 U3688 ( .A1(n2283), .A2(n2284), .A3(n2285), .A4(n2286), .ZN(n2282)
         );
  NAND3_X1 U3689 ( .A1(n5975), .A2(n5974), .A3(n5976), .ZN(n2286) );
  OAI211_X1 U3690 ( .C1(n5462), .C2(n5300), .A(n5972), .B(n5973), .ZN(n2285)
         );
  OAI222_X1 U3691 ( .A1(n5460), .A2(n5172), .B1(n5461), .B2(n5140), .C1(n5463), 
        .C2(n5268), .ZN(n2284) );
  OAI221_X1 U3692 ( .B1(n5433), .B2(n5076), .C1(n5434), .C2(n5108), .A(n2287), 
        .ZN(n2283) );
  AOI22_X1 U3693 ( .A1(n1742), .A2(n2103), .B1(n1743), .B2(n2104), .ZN(n2287)
         );
  AOI211_X1 U3696 ( .C1(n1744), .C2(n2105), .A(n2288), .B(n2289), .ZN(n2281)
         );
  OAI22_X1 U3697 ( .A1(n5443), .A2(n4724), .B1(n5453), .B2(n4628), .ZN(n2289)
         );
  OAI222_X1 U3698 ( .A1(n5448), .A2(n4564), .B1(n5454), .B2(n4532), .C1(n5449), 
        .C2(n4596), .ZN(n2288) );
  AOI221_X1 U3700 ( .B1(n2108), .B2(n1748), .C1(n2109), .C2(n2290), .A(n2291), 
        .ZN(n2280) );
  OAI22_X1 U3701 ( .A1(n4372), .A2(n6902), .B1(n4980), .B2(n2113), .ZN(n2291)
         );
  AOI222_X1 U3704 ( .A1(n1750), .A2(n2114), .B1(n2115), .B2(n1751), .C1(n1752), 
        .C2(n2116), .ZN(n2279) );
  NOR4_X1 U3711 ( .A1(n2296), .A2(n2297), .A3(n2298), .A4(n2299), .ZN(n2295)
         );
  NAND3_X1 U3712 ( .A1(n5985), .A2(n5984), .A3(n5986), .ZN(n2299) );
  OAI211_X1 U3713 ( .C1(n5462), .C2(n5301), .A(n5982), .B(n5983), .ZN(n2298)
         );
  OAI222_X1 U3714 ( .A1(n5460), .A2(n5173), .B1(n5461), .B2(n5141), .C1(n5463), 
        .C2(n5269), .ZN(n2297) );
  OAI221_X1 U3715 ( .B1(n5433), .B2(n5077), .C1(n5434), .C2(n5109), .A(n2300), 
        .ZN(n2296) );
  AOI22_X1 U3716 ( .A1(n1722), .A2(n2103), .B1(n1723), .B2(n2104), .ZN(n2300)
         );
  AOI211_X1 U3719 ( .C1(n1724), .C2(n2105), .A(n2301), .B(n2302), .ZN(n2294)
         );
  OAI22_X1 U3720 ( .A1(n5443), .A2(n4725), .B1(n5453), .B2(n4629), .ZN(n2302)
         );
  OAI222_X1 U3721 ( .A1(n5448), .A2(n4565), .B1(n5454), .B2(n4533), .C1(n5449), 
        .C2(n4597), .ZN(n2301) );
  AOI221_X1 U3723 ( .B1(n2108), .B2(n1728), .C1(n2109), .C2(n2303), .A(n2304), 
        .ZN(n2293) );
  OAI22_X1 U3724 ( .A1(n4373), .A2(n6902), .B1(n4981), .B2(n2113), .ZN(n2304)
         );
  AOI222_X1 U3727 ( .A1(n1730), .A2(n2114), .B1(n2115), .B2(n1731), .C1(n1732), 
        .C2(n2116), .ZN(n2292) );
  INV_X1 U3732 ( .A(n5997), .ZN(n5391) );
  AND4_X1 U3733 ( .A1(n2305), .A2(n2306), .A3(n2307), .A4(n2308), .ZN(n360) );
  NOR4_X1 U3734 ( .A1(n2309), .A2(n2310), .A3(n2311), .A4(n2312), .ZN(n2308)
         );
  NAND3_X1 U3735 ( .A1(n5995), .A2(n5994), .A3(n5996), .ZN(n2312) );
  OAI211_X1 U3736 ( .C1(n5462), .C2(n5302), .A(n5992), .B(n5993), .ZN(n2311)
         );
  OAI222_X1 U3737 ( .A1(n5460), .A2(n5174), .B1(n5461), .B2(n5142), .C1(n5463), 
        .C2(n5270), .ZN(n2310) );
  OAI221_X1 U3738 ( .B1(n5433), .B2(n5078), .C1(n5434), .C2(n5110), .A(n2313), 
        .ZN(n2309) );
  AOI22_X1 U3739 ( .A1(n1702), .A2(n2103), .B1(n1703), .B2(n2104), .ZN(n2313)
         );
  AOI211_X1 U3742 ( .C1(n1704), .C2(n2105), .A(n2314), .B(n2315), .ZN(n2307)
         );
  OAI22_X1 U3743 ( .A1(n5443), .A2(n4726), .B1(n5453), .B2(n4630), .ZN(n2315)
         );
  OAI222_X1 U3744 ( .A1(n5448), .A2(n4566), .B1(n5454), .B2(n4534), .C1(n5449), 
        .C2(n4598), .ZN(n2314) );
  AOI221_X1 U3746 ( .B1(n2108), .B2(n1708), .C1(n2109), .C2(n2316), .A(n2317), 
        .ZN(n2306) );
  OAI22_X1 U3747 ( .A1(n4374), .A2(n6902), .B1(n4982), .B2(n2113), .ZN(n2317)
         );
  AOI222_X1 U3750 ( .A1(n1710), .A2(n2114), .B1(n2115), .B2(n1711), .C1(n1712), 
        .C2(n2116), .ZN(n2305) );
  OAI222_X1 U3754 ( .A1(n5396), .A2(n5432), .B1(n5431), .B2(n854), .C1(n5394), 
        .C2(n5430), .ZN(\UUT/branch_rega [1]) );
  INV_X1 U3755 ( .A(n5955), .ZN(n5394) );
  AND4_X1 U3756 ( .A1(n2318), .A2(n2319), .A3(n2320), .A4(n2321), .ZN(n854) );
  NOR4_X1 U3757 ( .A1(n2322), .A2(n2323), .A3(n2324), .A4(n2325), .ZN(n2321)
         );
  NAND3_X1 U3758 ( .A1(n5953), .A2(n5952), .A3(n5954), .ZN(n2325) );
  OAI211_X1 U3759 ( .C1(n5462), .C2(n5303), .A(n5950), .B(n5951), .ZN(n2324)
         );
  OAI222_X1 U3760 ( .A1(n5460), .A2(n5175), .B1(n5461), .B2(n5143), .C1(n5463), 
        .C2(n5271), .ZN(n2323) );
  OAI221_X1 U3761 ( .B1(n5433), .B2(n5079), .C1(n5434), .C2(n5111), .A(n2326), 
        .ZN(n2322) );
  AOI22_X1 U3762 ( .A1(n1682), .A2(n2103), .B1(n1683), .B2(n2104), .ZN(n2326)
         );
  AOI211_X1 U3765 ( .C1(n1684), .C2(n2105), .A(n2327), .B(n2328), .ZN(n2320)
         );
  OAI22_X1 U3766 ( .A1(n5443), .A2(n4727), .B1(n5453), .B2(n4631), .ZN(n2328)
         );
  OAI222_X1 U3767 ( .A1(n5448), .A2(n4567), .B1(n5454), .B2(n4535), .C1(n5449), 
        .C2(n4599), .ZN(n2327) );
  AOI221_X1 U3769 ( .B1(n2108), .B2(n1688), .C1(n2109), .C2(n2329), .A(n2330), 
        .ZN(n2319) );
  OAI22_X1 U3770 ( .A1(n4375), .A2(n6901), .B1(n4983), .B2(n2113), .ZN(n2330)
         );
  AOI222_X1 U3773 ( .A1(n1690), .A2(n2114), .B1(n2115), .B2(n1691), .C1(n1692), 
        .C2(n2116), .ZN(n2318) );
  INV_X1 U3778 ( .A(n6010), .ZN(n5397) );
  AND4_X1 U3779 ( .A1(n2331), .A2(n2332), .A3(n2333), .A4(n2334), .ZN(n387) );
  NOR4_X1 U3780 ( .A1(n2335), .A2(n2336), .A3(n2337), .A4(n2338), .ZN(n2334)
         );
  NAND3_X1 U3781 ( .A1(n6008), .A2(n6007), .A3(n6009), .ZN(n2338) );
  OAI211_X1 U3782 ( .C1(n5462), .C2(n5304), .A(n6005), .B(n6006), .ZN(n2337)
         );
  OAI222_X1 U3783 ( .A1(n5460), .A2(n5176), .B1(n5461), .B2(n5144), .C1(n5463), 
        .C2(n5272), .ZN(n2336) );
  OAI221_X1 U3784 ( .B1(n5433), .B2(n5080), .C1(n5434), .C2(n5112), .A(n2339), 
        .ZN(n2335) );
  AOI22_X1 U3785 ( .A1(n1662), .A2(n2103), .B1(n1663), .B2(n2104), .ZN(n2339)
         );
  AOI211_X1 U3788 ( .C1(n1664), .C2(n2105), .A(n2340), .B(n2341), .ZN(n2333)
         );
  OAI22_X1 U3789 ( .A1(n5443), .A2(n4728), .B1(n5453), .B2(n4632), .ZN(n2341)
         );
  OAI222_X1 U3790 ( .A1(n5448), .A2(n4568), .B1(n5454), .B2(n4536), .C1(n5449), 
        .C2(n4600), .ZN(n2340) );
  AOI221_X1 U3792 ( .B1(n2108), .B2(n1668), .C1(n2109), .C2(n2342), .A(n2343), 
        .ZN(n2332) );
  OAI22_X1 U3793 ( .A1(n4376), .A2(n6902), .B1(n4984), .B2(n2113), .ZN(n2343)
         );
  AOI222_X1 U3796 ( .A1(n1670), .A2(n2114), .B1(n2115), .B2(n1671), .C1(n1672), 
        .C2(n2116), .ZN(n2331) );
  INV_X1 U3801 ( .A(n6023), .ZN(n5400) );
  NOR4_X1 U3803 ( .A1(n2348), .A2(n2349), .A3(n2350), .A4(n2351), .ZN(n2347)
         );
  NAND3_X1 U3804 ( .A1(n6021), .A2(n6020), .A3(n6022), .ZN(n2351) );
  OAI211_X1 U3805 ( .C1(n5462), .C2(n5305), .A(n6018), .B(n6019), .ZN(n2350)
         );
  OAI222_X1 U3806 ( .A1(n5460), .A2(n5177), .B1(n5461), .B2(n5145), .C1(n5463), 
        .C2(n5273), .ZN(n2349) );
  OAI221_X1 U3807 ( .B1(n5433), .B2(n5081), .C1(n5434), .C2(n5113), .A(n2352), 
        .ZN(n2348) );
  AOI22_X1 U3808 ( .A1(n1642), .A2(n2103), .B1(n1643), .B2(n2104), .ZN(n2352)
         );
  AOI211_X1 U3811 ( .C1(n1644), .C2(n2105), .A(n2353), .B(n2354), .ZN(n2346)
         );
  OAI22_X1 U3812 ( .A1(n5443), .A2(n4729), .B1(n5453), .B2(n4633), .ZN(n2354)
         );
  OAI222_X1 U3813 ( .A1(n5448), .A2(n4569), .B1(n5454), .B2(n4537), .C1(n5449), 
        .C2(n4601), .ZN(n2353) );
  AOI221_X1 U3815 ( .B1(n2108), .B2(n1648), .C1(n2109), .C2(n2355), .A(n2356), 
        .ZN(n2345) );
  OAI22_X1 U3816 ( .A1(n4377), .A2(n6901), .B1(n4985), .B2(n2113), .ZN(n2356)
         );
  AOI222_X1 U3819 ( .A1(n1650), .A2(n2114), .B1(n2115), .B2(n1651), .C1(n1652), 
        .C2(n2116), .ZN(n2344) );
  INV_X1 U3824 ( .A(n6044), .ZN(n5403) );
  AND4_X1 U3825 ( .A1(n2357), .A2(n2358), .A3(n2359), .A4(n2360), .ZN(n435) );
  NOR4_X1 U3826 ( .A1(n2361), .A2(n2362), .A3(n2363), .A4(n2364), .ZN(n2360)
         );
  NAND3_X1 U3827 ( .A1(n6042), .A2(n6041), .A3(n6043), .ZN(n2364) );
  OAI211_X1 U3828 ( .C1(n5462), .C2(n5306), .A(n6039), .B(n6040), .ZN(n2363)
         );
  OAI222_X1 U3829 ( .A1(n5460), .A2(n5178), .B1(n5461), .B2(n5146), .C1(n5463), 
        .C2(n5274), .ZN(n2362) );
  OAI221_X1 U3830 ( .B1(n5433), .B2(n5082), .C1(n5434), .C2(n5114), .A(n2365), 
        .ZN(n2361) );
  AOI22_X1 U3831 ( .A1(n1622), .A2(n2103), .B1(n1623), .B2(n2104), .ZN(n2365)
         );
  AOI211_X1 U3834 ( .C1(n1624), .C2(n2105), .A(n2366), .B(n2367), .ZN(n2359)
         );
  OAI22_X1 U3835 ( .A1(n5443), .A2(n4730), .B1(n5453), .B2(n4634), .ZN(n2367)
         );
  OAI222_X1 U3836 ( .A1(n5448), .A2(n4570), .B1(n5454), .B2(n4538), .C1(n5449), 
        .C2(n4602), .ZN(n2366) );
  AOI221_X1 U3838 ( .B1(n2108), .B2(n1628), .C1(n2109), .C2(n2368), .A(n2369), 
        .ZN(n2358) );
  OAI22_X1 U3839 ( .A1(n4378), .A2(n6902), .B1(n4986), .B2(n2113), .ZN(n2369)
         );
  AOI222_X1 U3842 ( .A1(n1630), .A2(n2114), .B1(n2115), .B2(n1631), .C1(n1632), 
        .C2(n2116), .ZN(n2357) );
  OAI222_X1 U3846 ( .A1(n5408), .A2(n5432), .B1(n5431), .B2(n464), .C1(n5406), 
        .C2(n5430), .ZN(\UUT/branch_rega [16]) );
  INV_X1 U3847 ( .A(n6056), .ZN(n5406) );
  AND4_X1 U3848 ( .A1(n2370), .A2(n2371), .A3(n2372), .A4(n2373), .ZN(n464) );
  NOR4_X1 U3849 ( .A1(n2374), .A2(n2375), .A3(n2376), .A4(n2377), .ZN(n2373)
         );
  NAND3_X1 U3850 ( .A1(n6054), .A2(n6053), .A3(n6055), .ZN(n2377) );
  OAI211_X1 U3851 ( .C1(n5462), .C2(n5307), .A(n6051), .B(n6052), .ZN(n2376)
         );
  OAI222_X1 U3852 ( .A1(n5460), .A2(n5179), .B1(n5461), .B2(n5147), .C1(n5463), 
        .C2(n5275), .ZN(n2375) );
  OAI221_X1 U3853 ( .B1(n5433), .B2(n5083), .C1(n5434), .C2(n5115), .A(n2378), 
        .ZN(n2374) );
  AOI22_X1 U3854 ( .A1(n1602), .A2(n2103), .B1(n1603), .B2(n2104), .ZN(n2378)
         );
  AOI211_X1 U3857 ( .C1(n1604), .C2(n2105), .A(n2379), .B(n2380), .ZN(n2372)
         );
  OAI22_X1 U3858 ( .A1(n5443), .A2(n4731), .B1(n5453), .B2(n4635), .ZN(n2380)
         );
  OAI222_X1 U3859 ( .A1(n5448), .A2(n4571), .B1(n5454), .B2(n4539), .C1(n5449), 
        .C2(n4603), .ZN(n2379) );
  AOI221_X1 U3861 ( .B1(n2108), .B2(n1608), .C1(n2109), .C2(n2381), .A(n2382), 
        .ZN(n2371) );
  OAI22_X1 U3862 ( .A1(n4379), .A2(n6901), .B1(n4987), .B2(n2113), .ZN(n2382)
         );
  AOI222_X1 U3865 ( .A1(n1610), .A2(n2114), .B1(n2115), .B2(n1611), .C1(n1612), 
        .C2(n2116), .ZN(n2370) );
  OAI222_X1 U3869 ( .A1(n5411), .A2(n5432), .B1(n5431), .B2(n492), .C1(n5409), 
        .C2(n5430), .ZN(\UUT/branch_rega [15]) );
  INV_X1 U3870 ( .A(n6067), .ZN(n5409) );
  AND4_X1 U3871 ( .A1(n2383), .A2(n2384), .A3(n2385), .A4(n2386), .ZN(n492) );
  NOR4_X1 U3872 ( .A1(n2387), .A2(n2388), .A3(n2389), .A4(n2390), .ZN(n2386)
         );
  NAND3_X1 U3873 ( .A1(n6065), .A2(n6064), .A3(n6066), .ZN(n2390) );
  OAI211_X1 U3874 ( .C1(n5462), .C2(n5308), .A(n6062), .B(n6063), .ZN(n2389)
         );
  OAI222_X1 U3875 ( .A1(n5460), .A2(n5180), .B1(n5461), .B2(n5148), .C1(n5463), 
        .C2(n5276), .ZN(n2388) );
  OAI221_X1 U3876 ( .B1(n5433), .B2(n5084), .C1(n5434), .C2(n5116), .A(n2391), 
        .ZN(n2387) );
  AOI22_X1 U3877 ( .A1(n1582), .A2(n2103), .B1(n1583), .B2(n2104), .ZN(n2391)
         );
  AOI211_X1 U3880 ( .C1(n1584), .C2(n2105), .A(n2392), .B(n2393), .ZN(n2385)
         );
  OAI22_X1 U3881 ( .A1(n5443), .A2(n4732), .B1(n5453), .B2(n4636), .ZN(n2393)
         );
  OAI222_X1 U3882 ( .A1(n5448), .A2(n4572), .B1(n5454), .B2(n4540), .C1(n5449), 
        .C2(n4604), .ZN(n2392) );
  AOI221_X1 U3884 ( .B1(n2108), .B2(n1588), .C1(n2109), .C2(n2394), .A(n2395), 
        .ZN(n2384) );
  OAI22_X1 U3885 ( .A1(n4380), .A2(n6902), .B1(n4988), .B2(n2113), .ZN(n2395)
         );
  AOI222_X1 U3888 ( .A1(n1590), .A2(n2114), .B1(n2115), .B2(n1591), .C1(n1592), 
        .C2(n2116), .ZN(n2383) );
  OAI222_X1 U3892 ( .A1(n5414), .A2(n5432), .B1(n5431), .B2(n519), .C1(n5412), 
        .C2(n5430), .ZN(\UUT/branch_rega [14]) );
  INV_X1 U3893 ( .A(n6081), .ZN(n5412) );
  AND4_X1 U3894 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(n519) );
  NOR4_X1 U3895 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2399)
         );
  NAND3_X1 U3896 ( .A1(n6079), .A2(n6078), .A3(n6080), .ZN(n2403) );
  OAI211_X1 U3897 ( .C1(n5462), .C2(n5309), .A(n6076), .B(n6077), .ZN(n2402)
         );
  OAI222_X1 U3898 ( .A1(n5460), .A2(n5181), .B1(n5461), .B2(n5149), .C1(n5463), 
        .C2(n5277), .ZN(n2401) );
  OAI221_X1 U3899 ( .B1(n5433), .B2(n5085), .C1(n5434), .C2(n5117), .A(n2404), 
        .ZN(n2400) );
  AOI22_X1 U3900 ( .A1(n1562), .A2(n2103), .B1(n1563), .B2(n2104), .ZN(n2404)
         );
  AOI211_X1 U3903 ( .C1(n1564), .C2(n2105), .A(n2405), .B(n2406), .ZN(n2398)
         );
  OAI22_X1 U3904 ( .A1(n5443), .A2(n4733), .B1(n5453), .B2(n4637), .ZN(n2406)
         );
  OAI222_X1 U3905 ( .A1(n5448), .A2(n4573), .B1(n5454), .B2(n4541), .C1(n5449), 
        .C2(n4605), .ZN(n2405) );
  AOI221_X1 U3907 ( .B1(n2108), .B2(n1568), .C1(n2109), .C2(n2407), .A(n2408), 
        .ZN(n2397) );
  OAI22_X1 U3908 ( .A1(n4381), .A2(n6901), .B1(n4989), .B2(n2113), .ZN(n2408)
         );
  AOI222_X1 U3911 ( .A1(n1570), .A2(n2114), .B1(n2115), .B2(n1571), .C1(n1572), 
        .C2(n2116), .ZN(n2396) );
  INV_X1 U3916 ( .A(n6091), .ZN(n5415) );
  AND4_X1 U3917 ( .A1(n2409), .A2(n2410), .A3(n2411), .A4(n2412), .ZN(n543) );
  NOR4_X1 U3918 ( .A1(n2413), .A2(n2414), .A3(n2415), .A4(n2416), .ZN(n2412)
         );
  NAND3_X1 U3919 ( .A1(n6089), .A2(n6088), .A3(n6090), .ZN(n2416) );
  OAI211_X1 U3920 ( .C1(n5462), .C2(n5310), .A(n6086), .B(n6087), .ZN(n2415)
         );
  OAI222_X1 U3921 ( .A1(n5460), .A2(n5182), .B1(n5461), .B2(n5150), .C1(n5463), 
        .C2(n5278), .ZN(n2414) );
  OAI221_X1 U3922 ( .B1(n5433), .B2(n5086), .C1(n5434), .C2(n5118), .A(n2417), 
        .ZN(n2413) );
  AOI22_X1 U3923 ( .A1(n1542), .A2(n2103), .B1(n1543), .B2(n2104), .ZN(n2417)
         );
  AOI211_X1 U3926 ( .C1(n1544), .C2(n2105), .A(n2418), .B(n2419), .ZN(n2411)
         );
  OAI22_X1 U3927 ( .A1(n5443), .A2(n4734), .B1(n5453), .B2(n4638), .ZN(n2419)
         );
  OAI222_X1 U3928 ( .A1(n5448), .A2(n4574), .B1(n5454), .B2(n4542), .C1(n5449), 
        .C2(n4606), .ZN(n2418) );
  AOI221_X1 U3930 ( .B1(n2108), .B2(n1548), .C1(n2109), .C2(n2420), .A(n2421), 
        .ZN(n2410) );
  OAI22_X1 U3931 ( .A1(n4382), .A2(n6902), .B1(n4990), .B2(n2113), .ZN(n2421)
         );
  AOI222_X1 U3934 ( .A1(n1550), .A2(n2114), .B1(n2115), .B2(n1551), .C1(n1552), 
        .C2(n2116), .ZN(n2409) );
  INV_X1 U3938 ( .A(\UUT/Mpath/the_alu/N491 ), .ZN(\UUT/Mpath/the_alu/N492 )
         );
  NAND2_X1 U3939 ( .A1(\UUT/Mcontrol/bp_logicB/memory_main ), .A2(n2422), .ZN(
        \UUT/Mcontrol/st_logic/N42 ) );
  INV_X1 U3940 ( .A(\UUT/Mcontrol/bp_logicB/exec_main ), .ZN(n2422) );
  OAI221_X1 U3941 ( .B1(n984), .B2(n978), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2423), .A(n2424), .ZN(
        \UUT/Mcontrol/Program_counter/N8 ) );
  AOI22_X1 U3942 ( .A1(n985), .A2(n7327), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [2]), .B2(n6932), .ZN(n2424) );
  INV_X1 U3945 ( .A(\UUT/branch_rega [2]), .ZN(n2423) );
  INV_X1 U3947 ( .A(n6209), .ZN(n5361) );
  AND4_X1 U3948 ( .A1(n2427), .A2(n2428), .A3(n2429), .A4(n2430), .ZN(n816) );
  NOR4_X1 U3949 ( .A1(n2431), .A2(n2432), .A3(n2433), .A4(n2434), .ZN(n2430)
         );
  NAND3_X1 U3950 ( .A1(n6207), .A2(n6206), .A3(n6208), .ZN(n2434) );
  OAI211_X1 U3951 ( .C1(n5462), .C2(n5292), .A(n6204), .B(n6205), .ZN(n2433)
         );
  OAI222_X1 U3952 ( .A1(n5460), .A2(n5164), .B1(n5461), .B2(n5132), .C1(n5463), 
        .C2(n5260), .ZN(n2432) );
  OAI221_X1 U3953 ( .B1(n5433), .B2(n5068), .C1(n5434), .C2(n5100), .A(n2435), 
        .ZN(n2431) );
  AOI22_X1 U3954 ( .A1(n1902), .A2(n2103), .B1(n1903), .B2(n2104), .ZN(n2435)
         );
  AOI211_X1 U3957 ( .C1(n1904), .C2(n2105), .A(n2436), .B(n2437), .ZN(n2429)
         );
  OAI22_X1 U3958 ( .A1(n5443), .A2(n4716), .B1(n5453), .B2(n4620), .ZN(n2437)
         );
  OAI222_X1 U3959 ( .A1(n5448), .A2(n4556), .B1(n5454), .B2(n4524), .C1(n5449), 
        .C2(n4588), .ZN(n2436) );
  AOI221_X1 U3961 ( .B1(n2108), .B2(n1908), .C1(n2109), .C2(n2438), .A(n2439), 
        .ZN(n2428) );
  OAI22_X1 U3962 ( .A1(n4364), .A2(n6902), .B1(n4972), .B2(n2113), .ZN(n2439)
         );
  AOI222_X1 U3965 ( .A1(n1910), .A2(n2114), .B1(n2115), .B2(n1911), .C1(n1912), 
        .C2(n2116), .ZN(n2427) );
  INV_X1 U3969 ( .A(\UUT/jar_in [2]), .ZN(n978) );
  OAI221_X1 U3970 ( .B1(n984), .B2(n968), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2440), .A(n2441), .ZN(
        \UUT/Mcontrol/Program_counter/N28 ) );
  AOI22_X1 U3971 ( .A1(n985), .A2(\UUT/break_code[12] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [12]), .B2(n983), .ZN(n2441) );
  OAI21_X1 U3972 ( .B1(n5905), .B2(n2260), .A(n2442), .ZN(\UUT/break_code[12] ) );
  NAND2_X1 U3973 ( .A1(n6224), .A2(n2262), .ZN(n2442) );
  INV_X1 U3975 ( .A(\UUT/branch_rega [12]), .ZN(n2440) );
  AND4_X1 U3978 ( .A1(n2443), .A2(n2444), .A3(n2445), .A4(n2446), .ZN(n568) );
  NOR4_X1 U3979 ( .A1(n2447), .A2(n2448), .A3(n2449), .A4(n2450), .ZN(n2446)
         );
  NAND3_X1 U3980 ( .A1(n6219), .A2(n6218), .A3(n6220), .ZN(n2450) );
  OAI211_X1 U3981 ( .C1(n5462), .C2(n5311), .A(n6216), .B(n6217), .ZN(n2449)
         );
  OAI222_X1 U3982 ( .A1(n5460), .A2(n5183), .B1(n5461), .B2(n5151), .C1(n5463), 
        .C2(n5279), .ZN(n2448) );
  OAI221_X1 U3983 ( .B1(n5433), .B2(n5087), .C1(n5434), .C2(n5119), .A(n2451), 
        .ZN(n2447) );
  AOI22_X1 U3984 ( .A1(n1522), .A2(n2103), .B1(n1523), .B2(n2104), .ZN(n2451)
         );
  AOI211_X1 U3987 ( .C1(n1524), .C2(n2105), .A(n2452), .B(n2453), .ZN(n2445)
         );
  OAI22_X1 U3988 ( .A1(n5443), .A2(n4735), .B1(n5453), .B2(n4639), .ZN(n2453)
         );
  OAI222_X1 U3989 ( .A1(n5448), .A2(n4575), .B1(n5454), .B2(n4543), .C1(n5449), 
        .C2(n4607), .ZN(n2452) );
  AOI221_X1 U3991 ( .B1(n2108), .B2(n1528), .C1(n2109), .C2(n2454), .A(n2455), 
        .ZN(n2444) );
  OAI22_X1 U3992 ( .A1(n4383), .A2(n6901), .B1(n4991), .B2(n2113), .ZN(n2455)
         );
  AOI222_X1 U3995 ( .A1(n1530), .A2(n2114), .B1(n2115), .B2(n1531), .C1(n1532), 
        .C2(n2116), .ZN(n2443) );
  INV_X1 U3999 ( .A(\UUT/jar_in [12]), .ZN(n968) );
  OAI221_X1 U4000 ( .B1(n984), .B2(n969), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2456), .A(n2457), .ZN(
        \UUT/Mcontrol/Program_counter/N26 ) );
  AOI22_X1 U4001 ( .A1(n985), .A2(\UUT/break_code[11] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [11]), .B2(n983), .ZN(n2457) );
  OAI21_X1 U4002 ( .B1(n5906), .B2(n2260), .A(n2458), .ZN(\UUT/break_code[11] ) );
  NAND2_X1 U4003 ( .A1(n6233), .A2(n2262), .ZN(n2458) );
  INV_X1 U4005 ( .A(\UUT/branch_rega [11]), .ZN(n2456) );
  OAI222_X1 U4006 ( .A1(n5423), .A2(n5432), .B1(n5431), .B2(n592), .C1(n5421), 
        .C2(n5430), .ZN(\UUT/branch_rega [11]) );
  INV_X1 U4007 ( .A(n6230), .ZN(n5421) );
  AND4_X1 U4008 ( .A1(n2459), .A2(n2460), .A3(n2461), .A4(n2462), .ZN(n592) );
  NOR4_X1 U4009 ( .A1(n2463), .A2(n2464), .A3(n2465), .A4(n2466), .ZN(n2462)
         );
  NAND3_X1 U4010 ( .A1(n6228), .A2(n6227), .A3(n6229), .ZN(n2466) );
  OAI211_X1 U4011 ( .C1(n5462), .C2(n5312), .A(n6225), .B(n6226), .ZN(n2465)
         );
  OAI222_X1 U4012 ( .A1(n5460), .A2(n5184), .B1(n5461), .B2(n5152), .C1(n5463), 
        .C2(n5280), .ZN(n2464) );
  OAI221_X1 U4013 ( .B1(n5433), .B2(n5088), .C1(n5434), .C2(n5120), .A(n2467), 
        .ZN(n2463) );
  AOI22_X1 U4014 ( .A1(n1502), .A2(n2103), .B1(n1503), .B2(n2104), .ZN(n2467)
         );
  AOI211_X1 U4017 ( .C1(n1504), .C2(n2105), .A(n2468), .B(n2469), .ZN(n2461)
         );
  OAI22_X1 U4018 ( .A1(n5443), .A2(n4736), .B1(n5453), .B2(n4640), .ZN(n2469)
         );
  OAI222_X1 U4019 ( .A1(n5448), .A2(n4576), .B1(n5454), .B2(n4544), .C1(n5449), 
        .C2(n4608), .ZN(n2468) );
  AOI221_X1 U4021 ( .B1(n2108), .B2(n1508), .C1(n2109), .C2(n2470), .A(n2471), 
        .ZN(n2460) );
  OAI22_X1 U4022 ( .A1(n4384), .A2(n6901), .B1(n4992), .B2(n2113), .ZN(n2471)
         );
  AOI222_X1 U4025 ( .A1(n1510), .A2(n2114), .B1(n2115), .B2(n1511), .C1(n1512), 
        .C2(n2116), .ZN(n2459) );
  INV_X1 U4029 ( .A(\UUT/jar_in [11]), .ZN(n969) );
  OAI221_X1 U4030 ( .B1(n984), .B2(n970), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2472), .A(n2473), .ZN(
        \UUT/Mcontrol/Program_counter/N24 ) );
  AOI22_X1 U4031 ( .A1(n985), .A2(\UUT/break_code[10] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [10]), .B2(n6932), .ZN(n2473) );
  OAI21_X1 U4032 ( .B1(n5762), .B2(n2260), .A(n2474), .ZN(\UUT/break_code[10] ) );
  NAND2_X1 U4033 ( .A1(n6283), .A2(n2262), .ZN(n2474) );
  INV_X1 U4035 ( .A(\UUT/branch_rega [10]), .ZN(n2472) );
  OAI222_X1 U4036 ( .A1(n5426), .A2(n5432), .B1(n5431), .B2(n615), .C1(n5424), 
        .C2(n5430), .ZN(\UUT/branch_rega [10]) );
  INV_X1 U4037 ( .A(n6239), .ZN(n5424) );
  AND4_X1 U4038 ( .A1(n2475), .A2(n2476), .A3(n2477), .A4(n2478), .ZN(n615) );
  NOR4_X1 U4039 ( .A1(n2479), .A2(n2480), .A3(n2481), .A4(n2482), .ZN(n2478)
         );
  NAND3_X1 U4040 ( .A1(n6237), .A2(n6236), .A3(n6238), .ZN(n2482) );
  OAI211_X1 U4041 ( .C1(n5462), .C2(n5313), .A(n6234), .B(n6235), .ZN(n2481)
         );
  OAI222_X1 U4042 ( .A1(n5460), .A2(n5185), .B1(n5461), .B2(n5153), .C1(n5463), 
        .C2(n5281), .ZN(n2480) );
  OAI221_X1 U4043 ( .B1(n5433), .B2(n5089), .C1(n5434), .C2(n5121), .A(n2483), 
        .ZN(n2479) );
  AOI22_X1 U4044 ( .A1(n1482), .A2(n2103), .B1(n1483), .B2(n2104), .ZN(n2483)
         );
  AOI211_X1 U4047 ( .C1(n1484), .C2(n2105), .A(n2484), .B(n2485), .ZN(n2477)
         );
  OAI22_X1 U4048 ( .A1(n5443), .A2(n4737), .B1(n5453), .B2(n4641), .ZN(n2485)
         );
  OAI222_X1 U4049 ( .A1(n5448), .A2(n4577), .B1(n5454), .B2(n4545), .C1(n5449), 
        .C2(n4609), .ZN(n2484) );
  AOI221_X1 U4051 ( .B1(n2108), .B2(n1488), .C1(n2109), .C2(n2486), .A(n2487), 
        .ZN(n2476) );
  OAI22_X1 U4052 ( .A1(n4385), .A2(n6901), .B1(n4993), .B2(n2113), .ZN(n2487)
         );
  AOI222_X1 U4055 ( .A1(n1490), .A2(n2114), .B1(n2115), .B2(n1491), .C1(n1492), 
        .C2(n2116), .ZN(n2475) );
  INV_X1 U4059 ( .A(\UUT/jar_in [10]), .ZN(n970) );
  OAI221_X1 U4060 ( .B1(n984), .B2(n971), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2488), .A(n2489), .ZN(
        \UUT/Mcontrol/Program_counter/N22 ) );
  AOI22_X1 U4061 ( .A1(n985), .A2(\UUT/break_code[9] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [9]), .B2(n983), .ZN(n2489) );
  OAI21_X1 U4062 ( .B1(n5769), .B2(n2260), .A(n2490), .ZN(\UUT/break_code[9] )
         );
  NAND2_X1 U4063 ( .A1(n6144), .A2(n2262), .ZN(n2490) );
  INV_X1 U4065 ( .A(\UUT/branch_rega [9]), .ZN(n2488) );
  OAI222_X1 U4066 ( .A1(n5335), .A2(n5432), .B1(n5431), .B2(n638), .C1(n5331), 
        .C2(n5430), .ZN(\UUT/branch_rega [9]) );
  INV_X1 U4067 ( .A(n6141), .ZN(n5331) );
  AND4_X1 U4068 ( .A1(n2491), .A2(n2492), .A3(n2493), .A4(n2494), .ZN(n638) );
  NOR4_X1 U4069 ( .A1(n2495), .A2(n2496), .A3(n2497), .A4(n2498), .ZN(n2494)
         );
  NAND3_X1 U4070 ( .A1(n6139), .A2(n6138), .A3(n6140), .ZN(n2498) );
  OAI211_X1 U4071 ( .C1(n5462), .C2(n5283), .A(n6136), .B(n6137), .ZN(n2497)
         );
  OAI222_X1 U4072 ( .A1(n5460), .A2(n5155), .B1(n5461), .B2(n5123), .C1(n5463), 
        .C2(n5251), .ZN(n2496) );
  OAI221_X1 U4073 ( .B1(n5433), .B2(n5059), .C1(n5434), .C2(n5091), .A(n2499), 
        .ZN(n2495) );
  AOI22_X1 U4074 ( .A1(n2082), .A2(n2103), .B1(n2083), .B2(n2104), .ZN(n2499)
         );
  AOI211_X1 U4077 ( .C1(n2084), .C2(n2105), .A(n2500), .B(n2501), .ZN(n2493)
         );
  OAI22_X1 U4078 ( .A1(n5443), .A2(n4707), .B1(n5453), .B2(n4611), .ZN(n2501)
         );
  OAI222_X1 U4079 ( .A1(n5448), .A2(n4547), .B1(n5454), .B2(n4515), .C1(n5449), 
        .C2(n4579), .ZN(n2500) );
  AOI221_X1 U4081 ( .B1(n2108), .B2(n2088), .C1(n2109), .C2(n2502), .A(n2503), 
        .ZN(n2492) );
  OAI22_X1 U4082 ( .A1(n4355), .A2(n6902), .B1(n4963), .B2(n2113), .ZN(n2503)
         );
  AOI222_X1 U4085 ( .A1(n2091), .A2(n2114), .B1(n2115), .B2(n2092), .C1(n2093), 
        .C2(n2116), .ZN(n2491) );
  INV_X1 U4089 ( .A(\UUT/jar_in [9]), .ZN(n971) );
  OAI221_X1 U4090 ( .B1(n984), .B2(n972), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2504), .A(n2505), .ZN(
        \UUT/Mcontrol/Program_counter/N20 ) );
  AOI22_X1 U4091 ( .A1(n985), .A2(\UUT/break_code[8] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [8]), .B2(n6932), .ZN(n2505) );
  OAI21_X1 U4092 ( .B1(n5776), .B2(n2260), .A(n2506), .ZN(\UUT/break_code[8] )
         );
  NAND2_X1 U4093 ( .A1(n6153), .A2(n2262), .ZN(n2506) );
  INV_X1 U4095 ( .A(\UUT/branch_rega [8]), .ZN(n2504) );
  INV_X1 U4097 ( .A(n6150), .ZN(n5337) );
  AND4_X1 U4098 ( .A1(n2507), .A2(n2508), .A3(n2509), .A4(n2510), .ZN(n662) );
  NOR4_X1 U4099 ( .A1(n2511), .A2(n2512), .A3(n2513), .A4(n2514), .ZN(n2510)
         );
  NAND3_X1 U4100 ( .A1(n6148), .A2(n6147), .A3(n6149), .ZN(n2514) );
  OAI211_X1 U4101 ( .C1(n5462), .C2(n5284), .A(n6145), .B(n6146), .ZN(n2513)
         );
  OAI222_X1 U4102 ( .A1(n5460), .A2(n5156), .B1(n5461), .B2(n5124), .C1(n5463), 
        .C2(n5252), .ZN(n2512) );
  OAI221_X1 U4103 ( .B1(n5433), .B2(n5060), .C1(n5434), .C2(n5092), .A(n2515), 
        .ZN(n2511) );
  AOI22_X1 U4104 ( .A1(n2062), .A2(n2103), .B1(n2063), .B2(n2104), .ZN(n2515)
         );
  AOI211_X1 U4107 ( .C1(n2064), .C2(n2105), .A(n2516), .B(n2517), .ZN(n2509)
         );
  OAI22_X1 U4108 ( .A1(n5443), .A2(n4708), .B1(n5453), .B2(n4612), .ZN(n2517)
         );
  OAI222_X1 U4109 ( .A1(n5448), .A2(n4548), .B1(n5454), .B2(n4516), .C1(n5449), 
        .C2(n4580), .ZN(n2516) );
  AOI221_X1 U4111 ( .B1(n2108), .B2(n2068), .C1(n2109), .C2(n2518), .A(n2519), 
        .ZN(n2508) );
  OAI22_X1 U4112 ( .A1(n4356), .A2(n6901), .B1(n4964), .B2(n2113), .ZN(n2519)
         );
  AOI222_X1 U4115 ( .A1(n2070), .A2(n2114), .B1(n2115), .B2(n2071), .C1(n2072), 
        .C2(n2116), .ZN(n2507) );
  INV_X1 U4119 ( .A(\UUT/jar_in [8]), .ZN(n972) );
  OAI221_X1 U4120 ( .B1(n984), .B2(n973), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2520), .A(n2521), .ZN(
        \UUT/Mcontrol/Program_counter/N18 ) );
  AOI22_X1 U4121 ( .A1(n985), .A2(\UUT/break_code[7] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [7]), .B2(n983), .ZN(n2521) );
  OAI21_X1 U4122 ( .B1(n5971), .B2(n2260), .A(n2522), .ZN(\UUT/break_code[7] )
         );
  NAND2_X1 U4123 ( .A1(n6162), .A2(n2262), .ZN(n2522) );
  INV_X1 U4125 ( .A(\UUT/branch_rega [7]), .ZN(n2520) );
  INV_X1 U4127 ( .A(n6159), .ZN(n5340) );
  NOR4_X1 U4129 ( .A1(n2527), .A2(n2528), .A3(n2529), .A4(n2530), .ZN(n2526)
         );
  NAND3_X1 U4130 ( .A1(n6157), .A2(n6156), .A3(n6158), .ZN(n2530) );
  OAI211_X1 U4131 ( .C1(n5462), .C2(n5285), .A(n6154), .B(n6155), .ZN(n2529)
         );
  OAI222_X1 U4132 ( .A1(n5460), .A2(n5157), .B1(n5461), .B2(n5125), .C1(n5463), 
        .C2(n5253), .ZN(n2528) );
  OAI221_X1 U4133 ( .B1(n5433), .B2(n5061), .C1(n5434), .C2(n5093), .A(n2531), 
        .ZN(n2527) );
  AOI22_X1 U4134 ( .A1(n2042), .A2(n2103), .B1(n2043), .B2(n2104), .ZN(n2531)
         );
  AOI211_X1 U4137 ( .C1(n2044), .C2(n2105), .A(n2532), .B(n2533), .ZN(n2525)
         );
  OAI22_X1 U4138 ( .A1(n5443), .A2(n4709), .B1(n5453), .B2(n4613), .ZN(n2533)
         );
  OAI222_X1 U4139 ( .A1(n5448), .A2(n4549), .B1(n5454), .B2(n4517), .C1(n5449), 
        .C2(n4581), .ZN(n2532) );
  AOI221_X1 U4141 ( .B1(n2108), .B2(n2048), .C1(n2109), .C2(n2534), .A(n2535), 
        .ZN(n2524) );
  OAI22_X1 U4142 ( .A1(n4357), .A2(n6901), .B1(n4965), .B2(n2113), .ZN(n2535)
         );
  AOI222_X1 U4145 ( .A1(n2050), .A2(n2114), .B1(n2115), .B2(n2051), .C1(n2052), 
        .C2(n2116), .ZN(n2523) );
  INV_X1 U4149 ( .A(\UUT/jar_in [7]), .ZN(n973) );
  OAI221_X1 U4150 ( .B1(n984), .B2(n974), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2536), .A(n2537), .ZN(
        \UUT/Mcontrol/Program_counter/N16 ) );
  AOI22_X1 U4151 ( .A1(n985), .A2(\UUT/break_code[6] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [6]), .B2(n6932), .ZN(n2537) );
  OAI21_X1 U4152 ( .B1(n6035), .B2(n2260), .A(n2538), .ZN(\UUT/break_code[6] )
         );
  NAND2_X1 U4153 ( .A1(n6171), .A2(n2262), .ZN(n2538) );
  INV_X1 U4155 ( .A(\UUT/branch_rega [6]), .ZN(n2536) );
  OAI222_X1 U4156 ( .A1(n5345), .A2(n5432), .B1(n5431), .B2(n711), .C1(n5343), 
        .C2(n5430), .ZN(\UUT/branch_rega [6]) );
  INV_X1 U4157 ( .A(n6168), .ZN(n5343) );
  AND4_X1 U4158 ( .A1(n2539), .A2(n2540), .A3(n2541), .A4(n2542), .ZN(n711) );
  NOR4_X1 U4159 ( .A1(n2543), .A2(n2544), .A3(n2545), .A4(n2546), .ZN(n2542)
         );
  NAND3_X1 U4160 ( .A1(n6166), .A2(n6165), .A3(n6167), .ZN(n2546) );
  OAI211_X1 U4161 ( .C1(n5462), .C2(n5286), .A(n6163), .B(n6164), .ZN(n2545)
         );
  OAI222_X1 U4162 ( .A1(n5460), .A2(n5158), .B1(n5461), .B2(n5126), .C1(n5463), 
        .C2(n5254), .ZN(n2544) );
  OAI221_X1 U4163 ( .B1(n5433), .B2(n5062), .C1(n5434), .C2(n5094), .A(n2547), 
        .ZN(n2543) );
  AOI22_X1 U4164 ( .A1(n2022), .A2(n2103), .B1(n2023), .B2(n2104), .ZN(n2547)
         );
  AOI211_X1 U4167 ( .C1(n2024), .C2(n2105), .A(n2548), .B(n2549), .ZN(n2541)
         );
  OAI22_X1 U4168 ( .A1(n5443), .A2(n4710), .B1(n5453), .B2(n4614), .ZN(n2549)
         );
  OAI222_X1 U4169 ( .A1(n5448), .A2(n4550), .B1(n5454), .B2(n4518), .C1(n5449), 
        .C2(n4582), .ZN(n2548) );
  AOI221_X1 U4171 ( .B1(n2108), .B2(n2028), .C1(n2109), .C2(n2550), .A(n2551), 
        .ZN(n2540) );
  OAI22_X1 U4172 ( .A1(n4358), .A2(n6902), .B1(n4966), .B2(n2113), .ZN(n2551)
         );
  AOI222_X1 U4175 ( .A1(n2030), .A2(n2114), .B1(n2115), .B2(n2031), .C1(n2032), 
        .C2(n2116), .ZN(n2539) );
  INV_X1 U4179 ( .A(\UUT/jar_in [6]), .ZN(n974) );
  OAI221_X1 U4180 ( .B1(n984), .B2(n975), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2552), .A(n2553), .ZN(
        \UUT/Mcontrol/Program_counter/N14 ) );
  AOI22_X1 U4181 ( .A1(n985), .A2(\UUT/break_code[5] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [5]), .B2(n6932), .ZN(n2553) );
  NAND2_X1 U4183 ( .A1(n6180), .A2(n2262), .ZN(n2554) );
  AND2_X1 U4184 ( .A1(n480), .A2(n6996), .ZN(n2262) );
  NOR2_X1 U4185 ( .A1(n7076), .A2(n1058), .ZN(n480) );
  NOR2_X1 U4187 ( .A1(n7076), .A2(n6996), .ZN(n2556) );
  INV_X1 U4199 ( .A(\UUT/branch_rega [5]), .ZN(n2552) );
  INV_X1 U4201 ( .A(n6177), .ZN(n5346) );
  AND4_X1 U4202 ( .A1(n2557), .A2(n2558), .A3(n2559), .A4(n2560), .ZN(n741) );
  NOR4_X1 U4203 ( .A1(n2561), .A2(n2562), .A3(n2563), .A4(n2564), .ZN(n2560)
         );
  NAND3_X1 U4204 ( .A1(n6175), .A2(n6174), .A3(n6176), .ZN(n2564) );
  OAI211_X1 U4205 ( .C1(n5462), .C2(n5287), .A(n6172), .B(n6173), .ZN(n2563)
         );
  OAI222_X1 U4206 ( .A1(n5460), .A2(n5159), .B1(n5461), .B2(n5127), .C1(n5463), 
        .C2(n5255), .ZN(n2562) );
  OAI221_X1 U4207 ( .B1(n5433), .B2(n5063), .C1(n5434), .C2(n5095), .A(n2565), 
        .ZN(n2561) );
  AOI22_X1 U4208 ( .A1(n2002), .A2(n2103), .B1(n2003), .B2(n2104), .ZN(n2565)
         );
  AOI211_X1 U4211 ( .C1(n2004), .C2(n2105), .A(n2566), .B(n2567), .ZN(n2559)
         );
  OAI22_X1 U4212 ( .A1(n5443), .A2(n4711), .B1(n5453), .B2(n4615), .ZN(n2567)
         );
  OAI222_X1 U4213 ( .A1(n5448), .A2(n4551), .B1(n5454), .B2(n4519), .C1(n5449), 
        .C2(n4583), .ZN(n2566) );
  AOI221_X1 U4215 ( .B1(n2108), .B2(n2008), .C1(n2109), .C2(n2568), .A(n2569), 
        .ZN(n2558) );
  OAI22_X1 U4216 ( .A1(n4359), .A2(n6901), .B1(n4967), .B2(n2113), .ZN(n2569)
         );
  AOI222_X1 U4219 ( .A1(n2010), .A2(n2114), .B1(n2115), .B2(n2011), .C1(n2012), 
        .C2(n2116), .ZN(n2557) );
  INV_X1 U4223 ( .A(\UUT/jar_in [5]), .ZN(n975) );
  OAI221_X1 U4224 ( .B1(n984), .B2(n976), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2570), .A(n2571), .ZN(
        \UUT/Mcontrol/Program_counter/N12 ) );
  AOI22_X1 U4225 ( .A1(n985), .A2(\UUT/break_code[4] ), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [4]), .B2(n6932), .ZN(n2571) );
  INV_X1 U4226 ( .A(n755), .ZN(\UUT/break_code[4] ) );
  AOI22_X1 U4227 ( .A1(n6190), .A2(n2425), .B1(n2426), .B2(n7202), .ZN(n755)
         );
  INV_X1 U4228 ( .A(\UUT/branch_rega [4]), .ZN(n2570) );
  OAI222_X1 U4229 ( .A1(n5351), .A2(n5432), .B1(n5431), .B2(n766), .C1(n5349), 
        .C2(n5430), .ZN(\UUT/branch_rega [4]) );
  INV_X1 U4230 ( .A(n6186), .ZN(n5349) );
  AND4_X1 U4231 ( .A1(n2572), .A2(n2573), .A3(n2574), .A4(n2575), .ZN(n766) );
  NOR4_X1 U4232 ( .A1(n2576), .A2(n2577), .A3(n2578), .A4(n2579), .ZN(n2575)
         );
  NAND3_X1 U4233 ( .A1(n6184), .A2(n6183), .A3(n6185), .ZN(n2579) );
  OAI211_X1 U4234 ( .C1(n5462), .C2(n5288), .A(n6181), .B(n6182), .ZN(n2578)
         );
  OAI222_X1 U4235 ( .A1(n5460), .A2(n5160), .B1(n5461), .B2(n5128), .C1(n5463), 
        .C2(n5256), .ZN(n2577) );
  OAI221_X1 U4236 ( .B1(n5433), .B2(n5064), .C1(n5434), .C2(n5096), .A(n2580), 
        .ZN(n2576) );
  AOI22_X1 U4237 ( .A1(n1982), .A2(n2103), .B1(n1983), .B2(n2104), .ZN(n2580)
         );
  AOI211_X1 U4240 ( .C1(n1984), .C2(n2105), .A(n2581), .B(n2582), .ZN(n2574)
         );
  OAI22_X1 U4241 ( .A1(n5443), .A2(n4712), .B1(n5453), .B2(n4616), .ZN(n2582)
         );
  OAI222_X1 U4242 ( .A1(n5448), .A2(n4552), .B1(n5454), .B2(n4520), .C1(n5449), 
        .C2(n4584), .ZN(n2581) );
  AOI221_X1 U4244 ( .B1(n2108), .B2(n1988), .C1(n2109), .C2(n2583), .A(n2584), 
        .ZN(n2573) );
  OAI22_X1 U4245 ( .A1(n4360), .A2(n6902), .B1(n4968), .B2(n2113), .ZN(n2584)
         );
  AOI222_X1 U4248 ( .A1(n1990), .A2(n2114), .B1(n2115), .B2(n1991), .C1(n1992), 
        .C2(n2116), .ZN(n2572) );
  INV_X1 U4252 ( .A(\UUT/jar_in [4]), .ZN(n976) );
  OAI221_X1 U4253 ( .B1(n984), .B2(n977), .C1(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .C2(n2585), .A(n2586), .ZN(
        \UUT/Mcontrol/Program_counter/N10 ) );
  AOI22_X1 U4254 ( .A1(n985), .A2(n7174), .B1(
        \UUT/Mcontrol/Nextpc_decoding/Bta [3]), .B2(n6932), .ZN(n2586) );
  OAI21_X1 U4258 ( .B1(n6189), .B2(n2589), .A(n2590), .ZN(n2426) );
  INV_X1 U4259 ( .A(n6215), .ZN(n2590) );
  INV_X1 U4261 ( .A(n2589), .ZN(n1132) );
  NAND2_X1 U4262 ( .A1(n5900), .A2(n6891), .ZN(n2589) );
  INV_X1 U4263 ( .A(n1058), .ZN(n5900) );
  INV_X1 U4266 ( .A(\UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(n2592) );
  INV_X1 U4267 ( .A(\UUT/branch_rega [3]), .ZN(n2585) );
  INV_X1 U4270 ( .A(n6198), .ZN(n5352) );
  AND4_X1 U4271 ( .A1(n2593), .A2(n2594), .A3(n2595), .A4(n2596), .ZN(n791) );
  NOR4_X1 U4272 ( .A1(n2597), .A2(n2598), .A3(n2599), .A4(n2600), .ZN(n2596)
         );
  NAND3_X1 U4273 ( .A1(n6196), .A2(n6195), .A3(n6197), .ZN(n2600) );
  OAI211_X1 U4274 ( .C1(n5462), .C2(n5289), .A(n6193), .B(n6194), .ZN(n2599)
         );
  OAI222_X1 U4275 ( .A1(n5460), .A2(n5161), .B1(n5461), .B2(n5129), .C1(n5463), 
        .C2(n5257), .ZN(n2598) );
  OAI221_X1 U4276 ( .B1(n5433), .B2(n5065), .C1(n5434), .C2(n5097), .A(n2601), 
        .ZN(n2597) );
  AOI22_X1 U4277 ( .A1(n1962), .A2(n2103), .B1(n1963), .B2(n2104), .ZN(n2601)
         );
  AOI211_X1 U4282 ( .C1(n1964), .C2(n2105), .A(n2602), .B(n2603), .ZN(n2595)
         );
  OAI22_X1 U4283 ( .A1(n5443), .A2(n4713), .B1(n5453), .B2(n4617), .ZN(n2603)
         );
  OAI222_X1 U4284 ( .A1(n5448), .A2(n4553), .B1(n5454), .B2(n4521), .C1(n5449), 
        .C2(n4585), .ZN(n2602) );
  AOI221_X1 U4287 ( .B1(n2108), .B2(n1968), .C1(n2109), .C2(n2604), .A(n2605), 
        .ZN(n2594) );
  OAI22_X1 U4288 ( .A1(n4361), .A2(n6902), .B1(n4969), .B2(n2113), .ZN(n2605)
         );
  INV_X1 U4295 ( .A(n6275), .ZN(n2606) );
  AOI222_X1 U4296 ( .A1(n1970), .A2(n2114), .B1(n2115), .B2(n1971), .C1(n1972), 
        .C2(n2116), .ZN(n2593) );
  AOI21_X1 U4304 ( .B1(n2607), .B2(n7375), .A(\UUT/byp_controlA[2] ), .ZN(n940) );
  INV_X1 U4305 ( .A(\UUT/regfile/N262 ), .ZN(n2607) );
  INV_X1 U4307 ( .A(\UUT/Mcontrol/st_logic/N47 ), .ZN(\UUT/byp_controlA[0] )
         );
  NAND2_X1 U4308 ( .A1(\UUT/Mcontrol/bp_logicA/memory_main ), .A2(n2608), .ZN(
        \UUT/Mcontrol/st_logic/N47 ) );
  INV_X1 U4309 ( .A(\UUT/Mcontrol/bp_logicA/exec_main ), .ZN(n2608) );
  INV_X1 U4310 ( .A(\UUT/jar_in [3]), .ZN(n977) );
  INV_X1 U4312 ( .A(n2587), .ZN(n2609) );
  OAI21_X1 U4313 ( .B1(\UUT/Mcontrol/Nextpc_decoding/N116 ), .B2(n2591), .A(
        \UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(n2587) );
  INV_X1 U4314 ( .A(\UUT/Mcontrol/st_logic/N65 ), .ZN(n2591) );
  INV_X1 U4315 ( .A(\UUT/Mcontrol/st_logic/N103 ), .ZN(n2588) );
  INV_X1 U4316 ( .A(n6891), .ZN(\UUT/Mcontrol/Operation_decoding32/N2085 ) );
  INV_X1 U4324 ( .A(\UUT/Mcontrol/Operation_decoding32/N1994 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1995 ) );
  AND4_X1 U4328 ( .A1(n4313), .A2(n4314), .A3(n4315), .A4(n4316), .ZN(
        d_select[31]) );
  NAND2_X1 U4329 ( .A1(n4317), .A2(n4318), .ZN(n4313) );
  INV_X1 U4330 ( .A(N35), .ZN(n4318) );
  AND3_X1 U4331 ( .A1(n4314), .A2(n4315), .A3(n4319), .ZN(d_select[23]) );
  OAI21_X1 U4332 ( .B1(N35), .B2(n4317), .A(n4316), .ZN(n4319) );
  INV_X1 U4333 ( .A(N31), .ZN(n4316) );
  NOR2_X1 U4334 ( .A1(N43), .A2(N42), .ZN(n4317) );
  INV_X1 U4335 ( .A(N27), .ZN(n4315) );
  INV_X1 U4336 ( .A(N22), .ZN(n4314) );
  OAI21_X1 U4337 ( .B1(N43), .B2(n4320), .A(n4321), .ZN(d_select[9]) );
  INV_X1 U4338 ( .A(N42), .ZN(n4320) );
  NAND2_X1 U4339 ( .A1(n4321), .A2(n4322), .ZN(d_select[7]) );
  INV_X1 U4340 ( .A(N43), .ZN(n4322) );
  NOR4_X1 U4341 ( .A1(N22), .A2(N27), .A3(N31), .A4(N35), .ZN(n4321) );
  OR2_X1 U4342 ( .A1(\UUT/Mcontrol/x_sampled_dmem_command[MW] ), .A2(
        \UUT/x_we ), .ZN(dmem_write) );
  AND2_X1 U4343 ( .A1(\UUT/Mcontrol/m_sampled_xrd[4] ), .A2(n5315), .ZN(
        \UUT/regfile/N358 ) );
  AND2_X1 U4344 ( .A1(\UUT/Mcontrol/m_sampled_xrd[3] ), .A2(n5315), .ZN(
        \UUT/rd_addr [3]) );
  AND2_X1 U4345 ( .A1(\UUT/Mcontrol/m_sampled_xrd[2] ), .A2(n5315), .ZN(
        \UUT/rd_addr [2]) );
  AND2_X1 U4346 ( .A1(\UUT/Mcontrol/m_sampled_xrd[1] ), .A2(n5315), .ZN(
        \UUT/rd_addr [1]) );
  OR2_X1 U4348 ( .A1(\UUT/Mcontrol/bp_logicA/memory_main ), .A2(
        \UUT/Mcontrol/bp_logicA/exec_main ), .ZN(\UUT/byp_controlA[2] ) );
  OAI222_X1 U4349 ( .A1(n5331), .A2(n99), .B1(n5333), .B2(n5334), .C1(n5335), 
        .C2(n5336), .ZN(\UUT/branch_regb [9]) );
  OAI222_X1 U4350 ( .A1(n5337), .A2(n99), .B1(n5338), .B2(n5334), .C1(n5339), 
        .C2(n5336), .ZN(\UUT/branch_regb [8]) );
  OAI222_X1 U4351 ( .A1(n5340), .A2(n5332), .B1(n5341), .B2(n5334), .C1(n5342), 
        .C2(n5336), .ZN(\UUT/branch_regb [7]) );
  OAI222_X1 U4352 ( .A1(n5343), .A2(n5332), .B1(n5344), .B2(n5334), .C1(n5345), 
        .C2(n5336), .ZN(\UUT/branch_regb [6]) );
  OAI222_X1 U4353 ( .A1(n5346), .A2(n99), .B1(n5347), .B2(n5334), .C1(n5348), 
        .C2(n5336), .ZN(\UUT/branch_regb [5]) );
  OAI222_X1 U4354 ( .A1(n5349), .A2(n5332), .B1(n5350), .B2(n5334), .C1(n5351), 
        .C2(n5336), .ZN(\UUT/branch_regb [4]) );
  OAI222_X1 U4355 ( .A1(n5352), .A2(n5332), .B1(n5353), .B2(n5334), .C1(n5354), 
        .C2(n5336), .ZN(\UUT/branch_regb [3]) );
  OAI222_X1 U4358 ( .A1(n5361), .A2(n5332), .B1(n5362), .B2(n5334), .C1(n5363), 
        .C2(n5336), .ZN(\UUT/branch_regb [2]) );
  OAI222_X1 U4360 ( .A1(n5367), .A2(n5332), .B1(n5368), .B2(n5334), .C1(n5369), 
        .C2(n5336), .ZN(\UUT/branch_regb [28]) );
  OAI222_X1 U4361 ( .A1(n5370), .A2(n5332), .B1(n5371), .B2(n5334), .C1(n5372), 
        .C2(n5336), .ZN(\UUT/branch_regb [27]) );
  OAI222_X1 U4363 ( .A1(n5376), .A2(n99), .B1(n5377), .B2(n5334), .C1(n5378), 
        .C2(n5336), .ZN(\UUT/branch_regb [25]) );
  OAI222_X1 U4364 ( .A1(n5379), .A2(n99), .B1(n5380), .B2(n5334), .C1(n5381), 
        .C2(n5336), .ZN(\UUT/branch_regb [24]) );
  OAI222_X1 U4366 ( .A1(n5385), .A2(n5332), .B1(n5386), .B2(n5334), .C1(n5387), 
        .C2(n5336), .ZN(\UUT/branch_regb [22]) );
  OAI222_X1 U4367 ( .A1(n5388), .A2(n99), .B1(n5389), .B2(n5334), .C1(n5390), 
        .C2(n5336), .ZN(\UUT/branch_regb [21]) );
  OAI222_X1 U4368 ( .A1(n5391), .A2(n99), .B1(n5392), .B2(n5334), .C1(n5393), 
        .C2(n5336), .ZN(\UUT/branch_regb [20]) );
  OAI222_X1 U4369 ( .A1(n5394), .A2(n99), .B1(n5395), .B2(n5334), .C1(n5396), 
        .C2(n5336), .ZN(\UUT/branch_regb [1]) );
  OAI222_X1 U4370 ( .A1(n5397), .A2(n99), .B1(n5398), .B2(n5334), .C1(n5399), 
        .C2(n5336), .ZN(\UUT/branch_regb [19]) );
  OAI222_X1 U4371 ( .A1(n5400), .A2(n99), .B1(n5401), .B2(n5334), .C1(n5402), 
        .C2(n5336), .ZN(\UUT/branch_regb [18]) );
  OAI222_X1 U4372 ( .A1(n5403), .A2(n99), .B1(n5404), .B2(n5334), .C1(n5405), 
        .C2(n5336), .ZN(\UUT/branch_regb [17]) );
  OAI222_X1 U4373 ( .A1(n5406), .A2(n5332), .B1(n5407), .B2(n5334), .C1(n5408), 
        .C2(n5336), .ZN(\UUT/branch_regb [16]) );
  OAI222_X1 U4374 ( .A1(n5409), .A2(n5332), .B1(n5410), .B2(n5334), .C1(n5411), 
        .C2(n5336), .ZN(\UUT/branch_regb [15]) );
  OAI222_X1 U4375 ( .A1(n5412), .A2(n5332), .B1(n5413), .B2(n5334), .C1(n5414), 
        .C2(n5336), .ZN(\UUT/branch_regb [14]) );
  OAI222_X1 U4376 ( .A1(n5415), .A2(n99), .B1(n5416), .B2(n5334), .C1(n5417), 
        .C2(n5336), .ZN(\UUT/branch_regb [13]) );
  OAI222_X1 U4377 ( .A1(n5418), .A2(n99), .B1(n5419), .B2(n5334), .C1(n5420), 
        .C2(n5336), .ZN(\UUT/branch_regb [12]) );
  OAI222_X1 U4378 ( .A1(n5421), .A2(n99), .B1(n5422), .B2(n5334), .C1(n5423), 
        .C2(n5336), .ZN(\UUT/branch_regb [11]) );
  OAI222_X1 U4379 ( .A1(n5424), .A2(n5332), .B1(n5425), .B2(n5334), .C1(n5426), 
        .C2(n5336), .ZN(\UUT/branch_regb [10]) );
  OAI222_X1 U4380 ( .A1(n5427), .A2(n99), .B1(n5428), .B2(n5334), .C1(n5429), 
        .C2(n5336), .ZN(\UUT/branch_regb [0]) );
  NAND2_X1 U4383 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(
        \UUT/Mcontrol/st_logic/N42 ), .ZN(n5332) );
  AOI22_X1 U4385 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][30] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][30] ), .ZN(n5435) );
  AOI22_X1 U4386 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][30] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][30] ), .ZN(n5440) );
  AOI22_X1 U4387 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][30] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][30] ), .ZN(n5445) );
  AOI22_X1 U4388 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][30] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][30] ), .ZN(n5450) );
  AOI22_X1 U4389 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][30] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][30] ), .ZN(n5457) );
  OAI22_X1 U4391 ( .A1(n5465), .A2(n5466), .B1(n5467), .B2(n5468), .ZN(n5464)
         );
  AOI22_X1 U4393 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][29] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][29] ), .ZN(n5469) );
  AOI22_X1 U4394 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][29] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][29] ), .ZN(n5470) );
  AOI22_X1 U4395 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][29] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][29] ), .ZN(n5471) );
  AOI22_X1 U4396 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][29] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][29] ), .ZN(n5472) );
  AOI22_X1 U4397 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][29] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][29] ), .ZN(n5473) );
  OAI222_X1 U4400 ( .A1(n5367), .A2(n5430), .B1(n5319), .B2(n5431), .C1(n5369), 
        .C2(n5432), .ZN(\UUT/branch_rega [28]) );
  AOI22_X1 U4401 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][28] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][28] ), .ZN(n5477) );
  AOI22_X1 U4402 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][28] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][28] ), .ZN(n5478) );
  AOI22_X1 U4403 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][28] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][28] ), .ZN(n5479) );
  AOI22_X1 U4404 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][28] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][28] ), .ZN(n5480) );
  AOI22_X1 U4405 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][28] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][28] ), .ZN(n5481) );
  OAI22_X1 U4407 ( .A1(n5483), .A2(n5466), .B1(n5484), .B2(n5468), .ZN(n5482)
         );
  OAI222_X1 U4408 ( .A1(n5370), .A2(n5430), .B1(n5320), .B2(n5431), .C1(n5372), 
        .C2(n5432), .ZN(\UUT/branch_rega [27]) );
  AOI22_X1 U4409 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][27] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][27] ), .ZN(n5485) );
  AOI22_X1 U4410 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][27] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][27] ), .ZN(n5486) );
  AOI22_X1 U4411 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][27] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][27] ), .ZN(n5487) );
  AOI22_X1 U4412 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][27] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][27] ), .ZN(n5488) );
  AOI22_X1 U4413 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][27] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][27] ), .ZN(n5489) );
  INV_X1 U4414 ( .A(n5490), .ZN(n5370) );
  OAI22_X1 U4415 ( .A1(n5491), .A2(n5466), .B1(n5492), .B2(n5468), .ZN(n5490)
         );
  OAI222_X1 U4416 ( .A1(n5373), .A2(n5430), .B1(n5321), .B2(n5431), .C1(n5375), 
        .C2(n5432), .ZN(\UUT/branch_rega [26]) );
  AOI22_X1 U4417 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][26] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][26] ), .ZN(n5493) );
  AOI22_X1 U4418 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][26] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][26] ), .ZN(n5494) );
  AOI22_X1 U4419 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][26] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][26] ), .ZN(n5495) );
  AOI22_X1 U4420 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][26] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][26] ), .ZN(n5496) );
  AOI22_X1 U4421 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][26] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][26] ), .ZN(n5497) );
  OAI22_X1 U4423 ( .A1(n5499), .A2(n5466), .B1(n5500), .B2(n5468), .ZN(n5498)
         );
  OAI222_X1 U4424 ( .A1(n5376), .A2(n5430), .B1(n5322), .B2(n5431), .C1(n5378), 
        .C2(n5432), .ZN(\UUT/branch_rega [25]) );
  AOI22_X1 U4425 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][25] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][25] ), .ZN(n5501) );
  AOI22_X1 U4426 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][25] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][25] ), .ZN(n5502) );
  AOI22_X1 U4427 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][25] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][25] ), .ZN(n5503) );
  AOI22_X1 U4428 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][25] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][25] ), .ZN(n5504) );
  AOI22_X1 U4429 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][25] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][25] ), .ZN(n5505) );
  OAI22_X1 U4431 ( .A1(n5507), .A2(n5466), .B1(n5508), .B2(n5468), .ZN(n5506)
         );
  OAI222_X1 U4432 ( .A1(n5379), .A2(n5430), .B1(n5323), .B2(n5431), .C1(n5381), 
        .C2(n5432), .ZN(\UUT/branch_rega [24]) );
  AOI22_X1 U4433 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][24] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][24] ), .ZN(n5509) );
  AOI22_X1 U4434 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][24] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][24] ), .ZN(n5510) );
  AOI22_X1 U4435 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][24] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][24] ), .ZN(n5511) );
  AOI22_X1 U4436 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][24] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][24] ), .ZN(n5512) );
  AOI22_X1 U4437 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][24] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][24] ), .ZN(n5513) );
  INV_X1 U4438 ( .A(n5514), .ZN(n5379) );
  OAI22_X1 U4439 ( .A1(n5515), .A2(n5466), .B1(n5516), .B2(n5468), .ZN(n5514)
         );
  AOI22_X1 U4441 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][0] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][0] ), .ZN(n5517) );
  AOI22_X1 U4442 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][0] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][0] ), .ZN(n5518) );
  AOI22_X1 U4443 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][0] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][0] ), .ZN(n5519) );
  AOI22_X1 U4444 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][0] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][0] ), .ZN(n5520) );
  AOI22_X1 U4445 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][0] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][0] ), .ZN(n5521) );
  INV_X1 U4446 ( .A(n5522), .ZN(n5427) );
  OAI222_X1 U4447 ( .A1(n5523), .A2(n5468), .B1(n5524), .B2(n5525), .C1(n5526), 
        .C2(n5466), .ZN(n5522) );
  AOI22_X1 U4448 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][9] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][9] ), .ZN(n5629) );
  AOI22_X1 U4449 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][9] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][9] ), .ZN(n5634) );
  AOI22_X1 U4450 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][9] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][9] ), .ZN(n5639) );
  AOI22_X1 U4451 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][9] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][9] ), .ZN(n5644) );
  AOI22_X1 U4452 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][9] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][9] ), .ZN(n5651) );
  AOI22_X1 U4453 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][8] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][8] ), .ZN(n5658) );
  AOI22_X1 U4454 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][8] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][8] ), .ZN(n5659) );
  AOI22_X1 U4455 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][8] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][8] ), .ZN(n5660) );
  AOI22_X1 U4456 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][8] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][8] ), .ZN(n5661) );
  AOI22_X1 U4457 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][8] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][8] ), .ZN(n5662) );
  OAI22_X1 U4458 ( .A1(n5666), .A2(n5667), .B1(n5668), .B2(n5669), .ZN(n5665)
         );
  INV_X1 U4459 ( .A(D_DATA_INBUS[31]), .ZN(n5668) );
  INV_X1 U4460 ( .A(D_DATA_INBUS[15]), .ZN(n5666) );
  AOI22_X1 U4461 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][7] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][7] ), .ZN(n5670) );
  AOI22_X1 U4462 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][7] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][7] ), .ZN(n5671) );
  AOI22_X1 U4463 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][7] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][7] ), .ZN(n5672) );
  AOI22_X1 U4464 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][7] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][7] ), .ZN(n5673) );
  AOI22_X1 U4465 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][7] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][7] ), .ZN(n5674) );
  OAI22_X1 U4466 ( .A1(n5667), .A2(n5676), .B1(n5669), .B2(n5677), .ZN(n5675)
         );
  INV_X1 U4467 ( .A(D_DATA_INBUS[30]), .ZN(n5677) );
  INV_X1 U4468 ( .A(D_DATA_INBUS[14]), .ZN(n5676) );
  INV_X1 U4469 ( .A(n5679), .ZN(n5678) );
  AOI22_X1 U4470 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[22]), 
        .B1(\UUT/Mpath/the_memhandle/N38 ), .B2(D_DATA_INBUS[14]), .ZN(n5679)
         );
  AOI22_X1 U4471 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][6] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][6] ), .ZN(n5680) );
  AOI22_X1 U4472 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][6] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][6] ), .ZN(n5681) );
  AOI22_X1 U4473 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][6] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][6] ), .ZN(n5682) );
  AOI22_X1 U4474 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][6] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][6] ), .ZN(n5683) );
  AOI22_X1 U4475 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][6] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][6] ), .ZN(n5684) );
  OAI22_X1 U4476 ( .A1(n5667), .A2(n5686), .B1(n5669), .B2(n5687), .ZN(n5685)
         );
  INV_X1 U4477 ( .A(D_DATA_INBUS[29]), .ZN(n5687) );
  INV_X1 U4478 ( .A(D_DATA_INBUS[13]), .ZN(n5686) );
  INV_X1 U4479 ( .A(n5689), .ZN(n5688) );
  AOI22_X1 U4480 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[21]), 
        .B1(\UUT/Mpath/the_memhandle/N38 ), .B2(D_DATA_INBUS[13]), .ZN(n5689)
         );
  AOI22_X1 U4481 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][5] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][5] ), .ZN(n5690) );
  AOI22_X1 U4482 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][5] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][5] ), .ZN(n5691) );
  AOI22_X1 U4483 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][5] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][5] ), .ZN(n5692) );
  AOI22_X1 U4484 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][5] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][5] ), .ZN(n5693) );
  AOI22_X1 U4485 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][5] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][5] ), .ZN(n5694) );
  OAI22_X1 U4486 ( .A1(n5667), .A2(n5696), .B1(n5669), .B2(n5697), .ZN(n5695)
         );
  INV_X1 U4487 ( .A(D_DATA_INBUS[28]), .ZN(n5697) );
  INV_X1 U4488 ( .A(D_DATA_INBUS[12]), .ZN(n5696) );
  INV_X1 U4489 ( .A(n5699), .ZN(n5698) );
  AOI22_X1 U4490 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[20]), 
        .B1(\UUT/Mpath/the_memhandle/N38 ), .B2(D_DATA_INBUS[12]), .ZN(n5699)
         );
  AOI22_X1 U4491 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][4] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][4] ), .ZN(n5700) );
  AOI22_X1 U4492 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][4] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][4] ), .ZN(n5701) );
  AOI22_X1 U4493 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][4] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][4] ), .ZN(n5702) );
  AOI22_X1 U4494 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][4] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][4] ), .ZN(n5703) );
  AOI22_X1 U4495 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][4] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][4] ), .ZN(n5704) );
  OAI22_X1 U4496 ( .A1(n5667), .A2(n5706), .B1(n5669), .B2(n5707), .ZN(n5705)
         );
  INV_X1 U4497 ( .A(D_DATA_INBUS[27]), .ZN(n5707) );
  INV_X1 U4498 ( .A(D_DATA_INBUS[11]), .ZN(n5706) );
  INV_X1 U4499 ( .A(n5709), .ZN(n5708) );
  AOI22_X1 U4500 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[19]), 
        .B1(\UUT/Mpath/the_memhandle/N38 ), .B2(D_DATA_INBUS[11]), .ZN(n5709)
         );
  AOI22_X1 U4501 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][3] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][3] ), .ZN(n5710) );
  AOI22_X1 U4502 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][3] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][3] ), .ZN(n5711) );
  AOI22_X1 U4503 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][3] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][3] ), .ZN(n5712) );
  AOI22_X1 U4504 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][3] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][3] ), .ZN(n5713) );
  AOI22_X1 U4505 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][3] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][3] ), .ZN(n5714) );
  AOI22_X1 U4506 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][31] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][31] ), .ZN(n5715) );
  AOI22_X1 U4507 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][31] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][31] ), .ZN(n5716) );
  AOI22_X1 U4508 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][31] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][31] ), .ZN(n5717) );
  AOI22_X1 U4509 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][31] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][31] ), .ZN(n5718) );
  AOI22_X1 U4510 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][31] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][31] ), .ZN(n5719) );
  AOI22_X1 U4511 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][30] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][30] ), .ZN(n5721) );
  AOI22_X1 U4512 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][30] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][30] ), .ZN(n5722) );
  AOI22_X1 U4513 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][30] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][30] ), .ZN(n5723) );
  AOI22_X1 U4514 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][30] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][30] ), .ZN(n5724) );
  AOI22_X1 U4515 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][30] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][30] ), .ZN(n5725) );
  OAI22_X1 U4516 ( .A1(n5667), .A2(n5727), .B1(n5669), .B2(n5728), .ZN(n5726)
         );
  INV_X1 U4517 ( .A(D_DATA_INBUS[26]), .ZN(n5728) );
  INV_X1 U4518 ( .A(D_DATA_INBUS[10]), .ZN(n5727) );
  INV_X1 U4519 ( .A(n5730), .ZN(n5729) );
  AOI22_X1 U4520 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[18]), 
        .B1(\UUT/Mpath/the_memhandle/N38 ), .B2(D_DATA_INBUS[10]), .ZN(n5730)
         );
  AOI22_X1 U4521 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][2] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][2] ), .ZN(n5731) );
  AOI22_X1 U4522 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][2] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][2] ), .ZN(n5732) );
  AOI22_X1 U4523 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][2] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][2] ), .ZN(n5733) );
  AOI22_X1 U4524 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][2] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][2] ), .ZN(n5734) );
  AOI22_X1 U4525 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][2] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][2] ), .ZN(n5735) );
  AOI22_X1 U4526 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][29] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][29] ), .ZN(n5736) );
  AOI22_X1 U4527 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][29] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][29] ), .ZN(n5737) );
  AOI22_X1 U4528 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][29] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][29] ), .ZN(n5738) );
  AOI22_X1 U4529 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][29] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][29] ), .ZN(n5739) );
  AOI22_X1 U4530 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][29] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][29] ), .ZN(n5740) );
  AOI22_X1 U4531 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][28] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][28] ), .ZN(n5741) );
  AOI22_X1 U4532 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][28] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][28] ), .ZN(n5742) );
  AOI22_X1 U4533 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][28] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][28] ), .ZN(n5743) );
  AOI22_X1 U4534 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][28] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][28] ), .ZN(n5744) );
  AOI22_X1 U4535 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][28] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][28] ), .ZN(n5745) );
  AOI22_X1 U4536 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][27] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][27] ), .ZN(n5746) );
  AOI22_X1 U4537 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][27] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][27] ), .ZN(n5747) );
  AOI22_X1 U4538 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][27] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][27] ), .ZN(n5748) );
  AOI22_X1 U4539 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][27] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][27] ), .ZN(n5749) );
  AOI22_X1 U4540 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][27] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][27] ), .ZN(n5750) );
  NOR2_X1 U4541 ( .A1(n5753), .A2(n5754), .ZN(n5751) );
  AOI22_X1 U4542 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][26] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][26] ), .ZN(n5755) );
  AOI22_X1 U4543 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][26] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][26] ), .ZN(n5756) );
  AOI22_X1 U4544 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][26] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][26] ), .ZN(n5757) );
  AOI22_X1 U4545 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][26] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][26] ), .ZN(n5758) );
  AOI22_X1 U4546 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][26] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][26] ), .ZN(n5759) );
  AOI22_X1 U4547 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][25] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][25] ), .ZN(n5763) );
  AOI22_X1 U4548 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][25] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][25] ), .ZN(n5764) );
  AOI22_X1 U4549 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][25] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][25] ), .ZN(n5765) );
  AOI22_X1 U4550 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][25] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][25] ), .ZN(n5766) );
  AOI22_X1 U4551 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][25] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][25] ), .ZN(n5767) );
  AOI22_X1 U4552 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][24] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][24] ), .ZN(n5770) );
  AOI22_X1 U4553 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][24] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][24] ), .ZN(n5771) );
  AOI22_X1 U4554 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][24] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][24] ), .ZN(n5772) );
  AOI22_X1 U4555 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][24] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][24] ), .ZN(n5773) );
  AOI22_X1 U4556 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][24] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][24] ), .ZN(n5774) );
  AOI22_X1 U4557 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][23] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][23] ), .ZN(n5777) );
  AOI22_X1 U4558 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][23] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][23] ), .ZN(n5778) );
  AOI22_X1 U4559 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][23] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][23] ), .ZN(n5779) );
  AOI22_X1 U4560 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][23] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][23] ), .ZN(n5780) );
  AOI22_X1 U4561 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][23] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][23] ), .ZN(n5781) );
  AOI22_X1 U4562 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][22] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][22] ), .ZN(n5782) );
  AOI22_X1 U4563 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][22] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][22] ), .ZN(n5783) );
  AOI22_X1 U4564 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][22] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][22] ), .ZN(n5784) );
  AOI22_X1 U4565 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][22] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][22] ), .ZN(n5785) );
  AOI22_X1 U4566 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][22] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][22] ), .ZN(n5786) );
  AOI22_X1 U4567 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][21] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][21] ), .ZN(n5787) );
  AOI22_X1 U4568 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][21] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][21] ), .ZN(n5788) );
  AOI22_X1 U4569 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][21] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][21] ), .ZN(n5789) );
  AOI22_X1 U4570 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][21] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][21] ), .ZN(n5790) );
  AOI22_X1 U4571 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][21] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][21] ), .ZN(n5791) );
  AOI22_X1 U4572 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][20] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][20] ), .ZN(n5792) );
  AOI22_X1 U4573 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][20] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][20] ), .ZN(n5793) );
  AOI22_X1 U4574 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][20] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][20] ), .ZN(n5794) );
  AOI22_X1 U4575 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][20] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][20] ), .ZN(n5795) );
  AOI22_X1 U4576 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][20] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][20] ), .ZN(n5796) );
  OAI22_X1 U4577 ( .A1(n5798), .A2(n5667), .B1(n5799), .B2(n5669), .ZN(n5797)
         );
  INV_X1 U4578 ( .A(D_DATA_INBUS[25]), .ZN(n5799) );
  INV_X1 U4579 ( .A(D_DATA_INBUS[9]), .ZN(n5798) );
  INV_X1 U4580 ( .A(n5801), .ZN(n5800) );
  AOI22_X1 U4581 ( .A1(\UUT/Mpath/the_memhandle/N39 ), .A2(D_DATA_INBUS[1]), 
        .B1(\UUT/Mpath/the_memhandle/N37 ), .B2(D_DATA_INBUS[17]), .ZN(n5801)
         );
  AOI22_X1 U4582 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][1] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][1] ), .ZN(n5802) );
  AOI22_X1 U4583 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][1] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][1] ), .ZN(n5803) );
  AOI22_X1 U4584 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][1] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][1] ), .ZN(n5804) );
  AOI22_X1 U4585 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][1] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][1] ), .ZN(n5805) );
  AOI22_X1 U4586 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][1] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][1] ), .ZN(n5806) );
  AOI22_X1 U4587 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][19] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][19] ), .ZN(n5807) );
  AOI22_X1 U4588 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][19] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][19] ), .ZN(n5808) );
  AOI22_X1 U4589 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][19] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][19] ), .ZN(n5809) );
  AOI22_X1 U4590 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][19] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][19] ), .ZN(n5810) );
  AOI22_X1 U4591 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][19] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][19] ), .ZN(n5811) );
  AOI22_X1 U4592 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][18] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][18] ), .ZN(n5812) );
  AOI22_X1 U4593 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][18] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][18] ), .ZN(n5813) );
  AOI22_X1 U4594 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][18] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][18] ), .ZN(n5814) );
  AOI22_X1 U4595 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][18] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][18] ), .ZN(n5815) );
  AOI22_X1 U4596 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][18] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][18] ), .ZN(n5816) );
  AOI22_X1 U4597 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][17] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][17] ), .ZN(n5817) );
  AOI22_X1 U4598 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][17] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][17] ), .ZN(n5818) );
  AOI22_X1 U4599 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][17] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][17] ), .ZN(n5819) );
  AOI22_X1 U4600 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][17] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][17] ), .ZN(n5820) );
  AOI22_X1 U4601 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][17] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][17] ), .ZN(n5821) );
  AOI22_X1 U4602 ( .A1(D_DATA_INBUS[15]), .A2(n5824), .B1(
        \UUT/Mpath/the_memhandle/N239 ), .B2(D_DATA_INBUS[31]), .ZN(n5822) );
  INV_X1 U4603 ( .A(\UUT/Mpath/the_memhandle/N239 ), .ZN(n5824) );
  AOI22_X1 U4604 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][16] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][16] ), .ZN(n5826) );
  AOI22_X1 U4605 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][16] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][16] ), .ZN(n5827) );
  AOI22_X1 U4606 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][16] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][16] ), .ZN(n5828) );
  AOI22_X1 U4607 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][16] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][16] ), .ZN(n5829) );
  AOI22_X1 U4608 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][16] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][16] ), .ZN(n5830) );
  AOI22_X1 U4609 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][15] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][15] ), .ZN(n5831) );
  AOI22_X1 U4610 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][15] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][15] ), .ZN(n5832) );
  AOI22_X1 U4611 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][15] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][15] ), .ZN(n5833) );
  AOI22_X1 U4612 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][15] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][15] ), .ZN(n5834) );
  AOI22_X1 U4613 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][15] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][15] ), .ZN(n5835) );
  AOI22_X1 U4614 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][14] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][14] ), .ZN(n5836) );
  AOI22_X1 U4615 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][14] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][14] ), .ZN(n5837) );
  AOI22_X1 U4616 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][14] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][14] ), .ZN(n5838) );
  AOI22_X1 U4617 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][14] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][14] ), .ZN(n5839) );
  AOI22_X1 U4618 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][14] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][14] ), .ZN(n5840) );
  AOI22_X1 U4619 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][13] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][13] ), .ZN(n5841) );
  AOI22_X1 U4620 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][13] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][13] ), .ZN(n5842) );
  AOI22_X1 U4621 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][13] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][13] ), .ZN(n5843) );
  AOI22_X1 U4622 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][13] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][13] ), .ZN(n5844) );
  AOI22_X1 U4623 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][13] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][13] ), .ZN(n5845) );
  AOI22_X1 U4624 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][12] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][12] ), .ZN(n5846) );
  AOI22_X1 U4625 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][12] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][12] ), .ZN(n5847) );
  AOI22_X1 U4626 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][12] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][12] ), .ZN(n5848) );
  AOI22_X1 U4627 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][12] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][12] ), .ZN(n5849) );
  AOI22_X1 U4628 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][12] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][12] ), .ZN(n5850) );
  AOI22_X1 U4629 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][11] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][11] ), .ZN(n5851) );
  AOI22_X1 U4630 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][11] ), .B1(n5636), 
        .B2(\UUT/regfile/reg_out[20][11] ), .ZN(n5852) );
  AOI22_X1 U4631 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][11] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][11] ), .ZN(n5853) );
  AOI22_X1 U4632 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][11] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][11] ), .ZN(n5854) );
  AOI22_X1 U4633 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][11] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][11] ), .ZN(n5855) );
  NOR2_X1 U4634 ( .A1(n5856), .A2(n5857), .ZN(n5626) );
  AOI221_X1 U4635 ( .B1(D_DATA_INBUS[31]), .B2(\UUT/Mpath/the_memhandle/N36 ), 
        .C1(D_DATA_INBUS[7]), .C2(\UUT/Mpath/the_memhandle/N39 ), .A(n5858), 
        .ZN(n5857) );
  INV_X1 U4636 ( .A(n5859), .ZN(n5858) );
  AOI22_X1 U4637 ( .A1(\UUT/Mpath/the_memhandle/N38 ), .A2(D_DATA_INBUS[15]), 
        .B1(\UUT/Mpath/the_memhandle/N37 ), .B2(D_DATA_INBUS[23]), .ZN(n5859)
         );
  NOR2_X1 U4638 ( .A1(n5823), .A2(n5860), .ZN(n5625) );
  NOR2_X1 U4639 ( .A1(n5861), .A2(n5823), .ZN(n5624) );
  AOI22_X1 U4640 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][10] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][10] ), .ZN(n5863) );
  AOI22_X1 U4641 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][10] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][10] ), .ZN(n5864) );
  AOI22_X1 U4642 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][10] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][10] ), .ZN(n5865) );
  AOI22_X1 U4643 ( .A1(n6356), .A2(\UUT/regfile/reg_out[29][10] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][10] ), .ZN(n5866) );
  AOI22_X1 U4644 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][10] ), .B1(n6346), 
        .B2(\UUT/regfile/reg_out[4][10] ), .ZN(n5867) );
  INV_X1 U4645 ( .A(\UUT/Mpath/the_memhandle/N34 ), .ZN(n5856) );
  OAI22_X1 U4646 ( .A1(n5869), .A2(n5667), .B1(n5870), .B2(n5669), .ZN(n5868)
         );
  NAND2_X1 U4647 ( .A1(\UUT/Mpath/the_memhandle/N74 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5669) );
  INV_X1 U4648 ( .A(D_DATA_INBUS[24]), .ZN(n5870) );
  NAND2_X1 U4649 ( .A1(\UUT/Mpath/the_memhandle/N76 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5667) );
  INV_X1 U4650 ( .A(D_DATA_INBUS[8]), .ZN(n5869) );
  OAI22_X1 U4651 ( .A1(n5862), .A2(\UUT/Mpath/the_memhandle/N243 ), .B1(
        \UUT/Mpath/the_memhandle/N72 ), .B2(n5861), .ZN(n5664) );
  INV_X1 U4652 ( .A(\UUT/Mpath/the_memhandle/N72 ), .ZN(n5862) );
  OAI21_X1 U4653 ( .B1(\UUT/Mpath/the_memhandle/N72 ), .B2(n5860), .A(n5871), 
        .ZN(n5663) );
  NAND2_X1 U4654 ( .A1(\UUT/Mpath/the_memhandle/N77 ), .A2(
        \UUT/Mpath/the_memhandle/N72 ), .ZN(n5871) );
  INV_X1 U4655 ( .A(n5861), .ZN(n5860) );
  NAND2_X1 U4656 ( .A1(\UUT/Mpath/the_memhandle/N239 ), .A2(n5825), .ZN(n5861)
         );
  INV_X1 U4657 ( .A(n5873), .ZN(n5872) );
  AOI22_X1 U4658 ( .A1(\UUT/Mpath/the_memhandle/N37 ), .A2(D_DATA_INBUS[16]), 
        .B1(\UUT/Mpath/the_memhandle/N39 ), .B2(D_DATA_INBUS[0]), .ZN(n5873)
         );
  AOI22_X1 U4659 ( .A1(n5630), .A2(\UUT/regfile/reg_out[19][0] ), .B1(n5631), 
        .B2(\UUT/regfile/reg_out[18][0] ), .ZN(n5874) );
  NAND3_X1 U4663 ( .A1(\UUT/rs2_addr [0]), .A2(n5878), .A3(n5875), .ZN(n5627)
         );
  AOI22_X1 U4665 ( .A1(n5635), .A2(\UUT/regfile/reg_out[21][0] ), .B1(n6344), 
        .B2(\UUT/regfile/reg_out[20][0] ), .ZN(n5881) );
  AND2_X1 U4666 ( .A1(n5879), .A2(n5882), .ZN(n5636) );
  NAND3_X1 U4668 ( .A1(n5876), .A2(\UUT/rs2_addr [2]), .A3(n5879), .ZN(n5633)
         );
  NAND4_X1 U4669 ( .A1(n5879), .A2(\UUT/rs2_addr [1]), .A3(\UUT/rs2_addr [0]), 
        .A4(\UUT/rs2_addr [2]), .ZN(n5632) );
  AOI22_X1 U4671 ( .A1(n5640), .A2(\UUT/regfile/reg_out[25][0] ), .B1(n5641), 
        .B2(\UUT/regfile/reg_out[24][0] ), .ZN(n5885) );
  NAND3_X1 U4674 ( .A1(n5876), .A2(\UUT/rs2_addr [4]), .A3(n5888), .ZN(n5638)
         );
  AOI22_X1 U4676 ( .A1(n6355), .A2(\UUT/regfile/reg_out[29][0] ), .B1(n5646), 
        .B2(\UUT/regfile/reg_out[28][0] ), .ZN(n5889) );
  NAND3_X1 U4679 ( .A1(n5890), .A2(\UUT/rs2_addr [4]), .A3(n5876), .ZN(n5643)
         );
  AOI22_X1 U4684 ( .A1(n5652), .A2(\UUT/regfile/reg_out[5][0] ), .B1(n6345), 
        .B2(\UUT/regfile/reg_out[4][0] ), .ZN(n5894) );
  AND3_X1 U4685 ( .A1(n5892), .A2(n5884), .A3(n5882), .ZN(n5653) );
  NAND3_X1 U4687 ( .A1(\UUT/rs2_addr [2]), .A2(n5892), .A3(n5893), .ZN(n5650)
         );
  NAND3_X1 U4688 ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/rs2_addr [2]), .A3(n5891), 
        .ZN(n5649) );
  NOR2_X1 U4692 ( .A1(n5892), .A2(n6933), .ZN(n5890) );
  INV_X1 U4698 ( .A(n5878), .ZN(\UUT/rs2_addr [1]) );
  AND2_X1 U4700 ( .A1(n5876), .A2(n5884), .ZN(n5893) );
  NOR2_X1 U4701 ( .A1(n5878), .A2(\UUT/rs2_addr [0]), .ZN(n5876) );
  NAND2_X1 U4703 ( .A1(\UUT/Mcontrol/d_sampled_finstr [17]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1873 ), .ZN(n5878) );
  NOR2_X1 U4704 ( .A1(n5892), .A2(\UUT/rs2_addr [2]), .ZN(n5888) );
  NAND2_X1 U4706 ( .A1(\UUT/Mcontrol/d_sampled_finstr [19]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1873 ), .ZN(n5892) );
  NAND2_X1 U4711 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(n5897), 
        .ZN(\UUT/rs2_addr [0]) );
  INV_X1 U4712 ( .A(\UUT/Mcontrol/st_logic/N2 ), .ZN(
        \UUT/Mcontrol/st_logic/load_stall ) );
  INV_X1 U4713 ( .A(\UUT/Mcontrol/st_logic/N8 ), .ZN(
        \UUT/Mcontrol/st_logic/branchmul_stall ) );
  INV_X1 U4714 ( .A(\UUT/Mcontrol/st_logic/N6 ), .ZN(
        \UUT/Mcontrol/st_logic/branchlw_stall ) );
  INV_X1 U4715 ( .A(\UUT/Mcontrol/st_logic/N4 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_regb ) );
  INV_X1 U4718 ( .A(\UUT/Mcontrol/st_logic/N7 ), .ZN(
        \UUT/Mcontrol/st_logic/branch_uses_main_exe_result ) );
  INV_X1 U4719 ( .A(\UUT/Mcontrol/st_logic/N10 ), .ZN(\UUT/Mcontrol/N19 ) );
  AOI21_X1 U4720 ( .B1(n7103), .B2(\UUT/Mcontrol/Operation_decoding32/N1952 ), 
        .A(n6904), .ZN(n5908) );
  NAND4_X1 U4721 ( .A1(n6994), .A2(n5914), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1907 ), .A4(n7131), .ZN(n5911) );
  NOR3_X1 U4722 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1958 ), .A2(n7180), 
        .A3(n5909), .ZN(n5914) );
  AOI21_X1 U4724 ( .B1(\UUT/Mcontrol/Operation_decoding32/N1928 ), .B2(n5916), 
        .A(\UUT/Mcontrol/Operation_decoding32/N1946 ), .ZN(n5922) );
  OAI21_X1 U4725 ( .B1(n5925), .B2(n5923), .A(n5926), .ZN(
        \UUT/Mcontrol/d_jump_type[2] ) );
  AOI21_X1 U4726 ( .B1(\UUT/Mcontrol/d_sampled_finstr [18]), .B2(n7110), .A(
        n5928), .ZN(n5925) );
  AOI21_X1 U4727 ( .B1(n5929), .B2(n5930), .A(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .ZN(n5928) );
  OAI21_X1 U4728 ( .B1(n5931), .B2(n5923), .A(n5926), .ZN(
        \UUT/Mcontrol/d_jump_type[1] ) );
  AOI21_X1 U4729 ( .B1(\UUT/Mcontrol/d_sampled_finstr [17]), .B2(n5932), .A(
        n7131), .ZN(n5931) );
  OAI21_X1 U4730 ( .B1(n5933), .B2(n5934), .A(n5926), .ZN(
        \UUT/Mcontrol/d_jump_type[0] ) );
  AOI221_X1 U4731 ( .B1(n5935), .B2(n5930), .C1(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .C2(
        \UUT/Mcontrol/d_sampled_finstr [16]), .A(n7046), .ZN(n5933) );
  INV_X1 U4732 ( .A(\UUT/Mcontrol/Operation_decoding32/N1940 ), .ZN(n5930) );
  OAI22_X1 U4733 ( .A1(n5897), .A2(n5937), .B1(
        \UUT/Mcontrol/Operation_decoding32/N1946 ), .B2(n5929), .ZN(n5935) );
  NOR2_X1 U4734 ( .A1(n5938), .A2(\UUT/Mcontrol/Operation_decoding32/N1934 ), 
        .ZN(n5929) );
  AOI21_X1 U4735 ( .B1(\UUT/Mcontrol/Operation_decoding32/N62 ), .B2(n6943), 
        .A(\UUT/Mcontrol/Operation_decoding32/N1928 ), .ZN(n5938) );
  INV_X1 U4742 ( .A(n7169), .ZN(n5945) );
  OAI211_X1 U4743 ( .C1(n5946), .C2(n5909), .A(n6879), .B(n7151), .ZN(n5947)
         );
  AOI22_X1 U4744 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][1] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][1] ), .ZN(n5950) );
  AOI22_X1 U4745 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][1] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][1] ), .ZN(n5951) );
  AOI22_X1 U4746 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][1] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][1] ), .ZN(n5952) );
  AOI22_X1 U4747 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][1] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][1] ), .ZN(n5953) );
  AOI22_X1 U4748 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][1] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][1] ), .ZN(n5954) );
  OAI222_X1 U4749 ( .A1(n5956), .A2(n5468), .B1(n5957), .B2(n5525), .C1(n5958), 
        .C2(n5466), .ZN(n5955) );
  INV_X1 U4750 ( .A(n7188), .ZN(\UUT/Mcontrol/d_instr [1]) );
  AOI22_X1 U4751 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][23] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][23] ), .ZN(n5961) );
  AOI22_X1 U4752 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][23] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][23] ), .ZN(n5962) );
  AOI22_X1 U4753 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][23] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][23] ), .ZN(n5963) );
  AOI22_X1 U4754 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][23] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][23] ), .ZN(n5964) );
  AOI22_X1 U4755 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][23] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][23] ), .ZN(n5965) );
  OAI21_X1 U4757 ( .B1(n5907), .B2(n5754), .A(n5761), .ZN(n5970) );
  AOI22_X1 U4759 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][22] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][22] ), .ZN(n5972) );
  AOI22_X1 U4760 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][22] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][22] ), .ZN(n5973) );
  AOI22_X1 U4761 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][22] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][22] ), .ZN(n5974) );
  AOI22_X1 U4762 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][22] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][22] ), .ZN(n5975) );
  AOI22_X1 U4763 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][22] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][22] ), .ZN(n5976) );
  OAI222_X1 U4764 ( .A1(n5978), .A2(n5468), .B1(n5979), .B2(n5525), .C1(n5980), 
        .C2(n5466), .ZN(n5977) );
  OAI21_X1 U4765 ( .B1(n5899), .B2(n5754), .A(n5761), .ZN(n5981) );
  AOI22_X1 U4766 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][21] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][21] ), .ZN(n5982) );
  AOI22_X1 U4767 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][21] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][21] ), .ZN(n5983) );
  AOI22_X1 U4768 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][21] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][21] ), .ZN(n5984) );
  AOI22_X1 U4769 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][21] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][21] ), .ZN(n5985) );
  AOI22_X1 U4770 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][21] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][21] ), .ZN(n5986) );
  OAI222_X1 U4771 ( .A1(n5988), .A2(n5468), .B1(n5989), .B2(n5525), .C1(n5990), 
        .C2(n5466), .ZN(n5987) );
  OAI21_X1 U4772 ( .B1(n5901), .B2(n5754), .A(n5761), .ZN(n5991) );
  AOI22_X1 U4774 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][20] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][20] ), .ZN(n5992) );
  AOI22_X1 U4775 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][20] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][20] ), .ZN(n5993) );
  AOI22_X1 U4776 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][20] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][20] ), .ZN(n5994) );
  AOI22_X1 U4777 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][20] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][20] ), .ZN(n5995) );
  AOI22_X1 U4778 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][20] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][20] ), .ZN(n5996) );
  OAI222_X1 U4779 ( .A1(n5998), .A2(n5468), .B1(n5999), .B2(n5525), .C1(n6000), 
        .C2(n5466), .ZN(n5997) );
  OAI21_X1 U4780 ( .B1(n5754), .B2(n5896), .A(n5761), .ZN(n6001) );
  OAI21_X1 U4781 ( .B1(n5720), .B2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A(n6003), .ZN(n5752) );
  AOI22_X1 U4782 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][19] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][19] ), .ZN(n6005) );
  AOI22_X1 U4783 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][19] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][19] ), .ZN(n6006) );
  AOI22_X1 U4784 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][19] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][19] ), .ZN(n6007) );
  AOI22_X1 U4785 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][19] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][19] ), .ZN(n6008) );
  AOI22_X1 U4786 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][19] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][19] ), .ZN(n6009) );
  OAI222_X1 U4787 ( .A1(n6011), .A2(n5468), .B1(n6012), .B2(n5525), .C1(n6013), 
        .C2(n5466), .ZN(n6010) );
  OAI221_X1 U4788 ( .B1(n5904), .B2(n6004), .C1(n5753), .C2(n7225), .A(n6003), 
        .ZN(n6015) );
  AOI22_X1 U4789 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][18] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][18] ), .ZN(n6018) );
  AOI22_X1 U4790 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][18] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][18] ), .ZN(n6019) );
  AOI22_X1 U4791 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][18] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][18] ), .ZN(n6020) );
  AOI22_X1 U4792 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][18] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][18] ), .ZN(n6021) );
  AOI22_X1 U4793 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][18] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][18] ), .ZN(n6022) );
  OAI222_X1 U4794 ( .A1(n6024), .A2(n5468), .B1(n6025), .B2(n5525), .C1(n6026), 
        .C2(n5466), .ZN(n6023) );
  OAI221_X1 U4795 ( .B1(n6004), .B2(n5897), .C1(n5760), .C2(n7225), .A(n6003), 
        .ZN(n6027) );
  AND2_X1 U4796 ( .A1(n6028), .A2(n6029), .ZN(n6003) );
  OR3_X1 U4797 ( .A1(n5923), .A2(n7131), .A3(n5720), .ZN(n6029) );
  NAND2_X1 U4798 ( .A1(n5934), .A2(n7021), .ZN(n6004) );
  NAND3_X1 U4800 ( .A1(n6032), .A2(n7341), .A3(n6034), .ZN(n6031) );
  INV_X1 U4811 ( .A(n7139), .ZN(\UUT/Mcontrol/d_instr [0]) );
  AOI22_X1 U4812 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][17] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][17] ), .ZN(n6039) );
  AOI22_X1 U4813 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][17] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][17] ), .ZN(n6040) );
  AOI22_X1 U4814 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][17] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][17] ), .ZN(n6041) );
  AOI22_X1 U4815 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][17] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][17] ), .ZN(n6042) );
  AOI22_X1 U4816 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][17] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][17] ), .ZN(n6043) );
  OAI222_X1 U4817 ( .A1(n6045), .A2(n5468), .B1(n6046), .B2(n5525), .C1(n6047), 
        .C2(n5466), .ZN(n6044) );
  OAI221_X1 U4818 ( .B1(n7225), .B2(n5768), .C1(n6049), .C2(n5720), .A(n6028), 
        .ZN(n6048) );
  INV_X1 U4819 ( .A(n7083), .ZN(n6049) );
  AOI22_X1 U4820 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][16] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][16] ), .ZN(n6051) );
  AOI22_X1 U4821 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][16] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][16] ), .ZN(n6052) );
  AOI22_X1 U4822 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][16] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][16] ), .ZN(n6053) );
  AOI22_X1 U4823 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][16] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][16] ), .ZN(n6054) );
  AOI22_X1 U4824 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][16] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][16] ), .ZN(n6055) );
  OAI222_X1 U4825 ( .A1(n6057), .A2(n5468), .B1(n6058), .B2(n5525), .C1(n6059), 
        .C2(n5466), .ZN(n6056) );
  OAI221_X1 U4826 ( .B1(n7168), .B2(n5902), .C1(n5775), .C2(n7225), .A(n6028), 
        .ZN(n6060) );
  AOI22_X1 U4827 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][15] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][15] ), .ZN(n6062) );
  AOI22_X1 U4828 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][15] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][15] ), .ZN(n6063) );
  AOI22_X1 U4829 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][15] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][15] ), .ZN(n6064) );
  AOI22_X1 U4830 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][15] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][15] ), .ZN(n6065) );
  AOI22_X1 U4831 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][15] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][15] ), .ZN(n6066) );
  OAI222_X1 U4832 ( .A1(n6068), .A2(n5468), .B1(n6069), .B2(n5525), .C1(n6070), 
        .C2(n5466), .ZN(n6067) );
  AOI21_X1 U4834 ( .B1(n6849), .B2(n6075), .A(n6016), .ZN(n6074) );
  NOR2_X1 U4835 ( .A1(n5720), .A2(n6996), .ZN(n6016) );
  OAI221_X1 U4836 ( .B1(n7168), .B2(n5903), .C1(n5907), .C2(n7225), .A(n6028), 
        .ZN(n6075) );
  NAND2_X1 U4837 ( .A1(n7009), .A2(\UUT/Mcontrol/d_sampled_finstr [15]), .ZN(
        n6028) );
  AOI22_X1 U4838 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][14] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][14] ), .ZN(n6076) );
  AOI22_X1 U4839 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][14] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][14] ), .ZN(n6077) );
  AOI22_X1 U4840 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][14] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][14] ), .ZN(n6078) );
  AOI22_X1 U4841 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][14] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][14] ), .ZN(n6079) );
  AOI22_X1 U4842 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][14] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][14] ), .ZN(n6080) );
  OAI222_X1 U4843 ( .A1(n6082), .A2(n5468), .B1(n6083), .B2(n5525), .C1(n6084), 
        .C2(n5466), .ZN(n6081) );
  AOI22_X1 U4845 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][13] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][13] ), .ZN(n6086) );
  AOI22_X1 U4846 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][13] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][13] ), .ZN(n6087) );
  AOI22_X1 U4847 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][13] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][13] ), .ZN(n6088) );
  AOI22_X1 U4848 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][13] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][13] ), .ZN(n6089) );
  AOI22_X1 U4849 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][13] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][13] ), .ZN(n6090) );
  OAI222_X1 U4850 ( .A1(n6092), .A2(n5468), .B1(n6093), .B2(n5525), .C1(n6094), 
        .C2(n5466), .ZN(n6091) );
  AOI21_X1 U4852 ( .B1(n6132), .B2(n7105), .A(
        \UUT/Mcontrol/Operation_decoding32/N2043 ), .ZN(n6131) );
  OAI21_X1 U4853 ( .B1(n6133), .B2(n5944), .A(n7108), .ZN(n6132) );
  INV_X1 U4855 ( .A(n6890), .ZN(n5934) );
  AOI22_X1 U4856 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][9] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][9] ), .ZN(n6136) );
  AOI22_X1 U4857 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][9] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][9] ), .ZN(n6137) );
  AOI22_X1 U4858 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][9] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][9] ), .ZN(n6138) );
  AOI22_X1 U4859 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][9] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][9] ), .ZN(n6139) );
  AOI22_X1 U4860 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][9] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][9] ), .ZN(n6140) );
  OAI222_X1 U4861 ( .A1(n6142), .A2(n5468), .B1(n6143), .B2(n5525), .C1(n6096), 
        .C2(n5466), .ZN(n6141) );
  OAI222_X1 U4862 ( .A1(n6956), .A2(n5720), .B1(n7069), .B2(n5971), .C1(n5769), 
        .C2(n7021), .ZN(n6144) );
  AOI22_X1 U4863 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][8] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][8] ), .ZN(n6145) );
  AOI22_X1 U4864 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][8] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][8] ), .ZN(n6146) );
  AOI22_X1 U4865 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][8] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][8] ), .ZN(n6147) );
  AOI22_X1 U4866 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][8] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][8] ), .ZN(n6148) );
  AOI22_X1 U4867 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][8] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][8] ), .ZN(n6149) );
  OAI222_X1 U4868 ( .A1(n6151), .A2(n5468), .B1(n6152), .B2(n5525), .C1(n6098), 
        .C2(n5466), .ZN(n6150) );
  OAI222_X1 U4869 ( .A1(n6956), .A2(n5902), .B1(n7168), .B2(n6035), .C1(n7021), 
        .C2(n5776), .ZN(n6153) );
  AOI22_X1 U4870 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][7] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][7] ), .ZN(n6154) );
  AOI22_X1 U4871 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][7] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][7] ), .ZN(n6155) );
  AOI22_X1 U4872 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][7] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][7] ), .ZN(n6156) );
  AOI22_X1 U4873 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][7] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][7] ), .ZN(n6157) );
  AOI22_X1 U4874 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][7] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][7] ), .ZN(n6158) );
  OAI222_X1 U4875 ( .A1(n6160), .A2(n5468), .B1(n6161), .B2(n5525), .C1(n6100), 
        .C2(n5466), .ZN(n6159) );
  AOI22_X1 U4877 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][6] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][6] ), .ZN(n6163) );
  AOI22_X1 U4878 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][6] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][6] ), .ZN(n6164) );
  AOI22_X1 U4879 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][6] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][6] ), .ZN(n6165) );
  AOI22_X1 U4880 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][6] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][6] ), .ZN(n6166) );
  AOI22_X1 U4881 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][6] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][6] ), .ZN(n6167) );
  OAI222_X1 U4882 ( .A1(n6169), .A2(n5468), .B1(n6170), .B2(n5525), .C1(n6102), 
        .C2(n5466), .ZN(n6168) );
  AOI22_X1 U4884 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][5] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][5] ), .ZN(n6172) );
  AOI22_X1 U4885 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][5] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][5] ), .ZN(n6173) );
  AOI22_X1 U4886 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][5] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][5] ), .ZN(n6174) );
  AOI22_X1 U4887 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][5] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][5] ), .ZN(n6175) );
  AOI22_X1 U4888 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][5] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][5] ), .ZN(n6176) );
  OAI222_X1 U4889 ( .A1(n6178), .A2(n5468), .B1(n6179), .B2(n5525), .C1(n6104), 
        .C2(n5466), .ZN(n6177) );
  AOI22_X1 U4891 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][4] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][4] ), .ZN(n6181) );
  AOI22_X1 U4892 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][4] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][4] ), .ZN(n6182) );
  AOI22_X1 U4893 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][4] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][4] ), .ZN(n6183) );
  AOI22_X1 U4894 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][4] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][4] ), .ZN(n6184) );
  AOI22_X1 U4895 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][4] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][4] ), .ZN(n6185) );
  OAI222_X1 U4896 ( .A1(n6187), .A2(n5468), .B1(n6188), .B2(n5525), .C1(n6106), 
        .C2(n5466), .ZN(n6186) );
  OAI22_X1 U4897 ( .A1(n5762), .A2(n6030), .B1(n6191), .B2(n7179), .ZN(n6190)
         );
  AOI22_X1 U4898 ( .A1(n6849), .A2(n6192), .B1(\UUT/Mcontrol/d_instr [4]), 
        .B2(n6134), .ZN(n6191) );
  OAI222_X1 U4900 ( .A1(n6017), .A2(n5762), .B1(n7069), .B2(n7210), .C1(n7221), 
        .C2(n7020), .ZN(n6192) );
  AOI22_X1 U4901 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][3] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][3] ), .ZN(n6193) );
  AOI22_X1 U4902 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][3] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][3] ), .ZN(n6194) );
  AOI22_X1 U4903 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][3] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][3] ), .ZN(n6195) );
  AOI22_X1 U4904 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][3] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][3] ), .ZN(n6196) );
  AOI22_X1 U4905 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][3] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][3] ), .ZN(n6197) );
  OAI222_X1 U4906 ( .A1(n6199), .A2(n5468), .B1(n6200), .B2(n5525), .C1(n6108), 
        .C2(n5466), .ZN(n6198) );
  OAI22_X1 U4907 ( .A1(n5769), .A2(n6030), .B1(n6202), .B2(n7179), .ZN(n6201)
         );
  OAI222_X1 U4910 ( .A1(n6017), .A2(n5769), .B1(n7060), .B2(n5329), .C1(n7022), 
        .C2(n5327), .ZN(n6203) );
  AOI22_X1 U4911 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][2] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][2] ), .ZN(n6204) );
  AOI22_X1 U4912 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][2] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][2] ), .ZN(n6205) );
  AOI22_X1 U4913 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][2] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][2] ), .ZN(n6206) );
  AOI22_X1 U4914 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][2] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][2] ), .ZN(n6207) );
  AOI22_X1 U4915 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][2] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][2] ), .ZN(n6208) );
  OAI222_X1 U4916 ( .A1(n6210), .A2(n5468), .B1(n6211), .B2(n5525), .C1(n6112), 
        .C2(n5466), .ZN(n6209) );
  NAND2_X1 U4921 ( .A1(n7100), .A2(n7049), .ZN(n6030) );
  AND2_X1 U4922 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2085 ), .A2(n5900), 
        .ZN(n6215) );
  NOR2_X1 U4923 ( .A1(n7051), .A2(\UUT/Mcontrol/Operation_decoding32/N2079 ), 
        .ZN(n6189) );
  AOI22_X1 U4924 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][12] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][12] ), .ZN(n6216) );
  AOI22_X1 U4925 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][12] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][12] ), .ZN(n6217) );
  AOI22_X1 U4926 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][12] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][12] ), .ZN(n6218) );
  AOI22_X1 U4927 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][12] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][12] ), .ZN(n6219) );
  AOI22_X1 U4928 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][12] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][12] ), .ZN(n6220) );
  OAI222_X1 U4929 ( .A1(n6222), .A2(n5468), .B1(n6223), .B2(n5525), .C1(n6125), 
        .C2(n5466), .ZN(n6221) );
  AOI22_X1 U4931 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][11] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][11] ), .ZN(n6225) );
  AOI22_X1 U4932 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][11] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][11] ), .ZN(n6226) );
  AOI22_X1 U4933 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][11] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][11] ), .ZN(n6227) );
  AOI22_X1 U4934 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][11] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][11] ), .ZN(n6228) );
  AOI22_X1 U4935 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][11] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][11] ), .ZN(n6229) );
  OAI222_X1 U4936 ( .A1(n6231), .A2(n5468), .B1(n6232), .B2(n5525), .C1(n6127), 
        .C2(n5466), .ZN(n6230) );
  AOI22_X1 U4938 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][10] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][10] ), .ZN(n6234) );
  AOI22_X1 U4939 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][10] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][10] ), .ZN(n6235) );
  AOI22_X1 U4940 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][10] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][10] ), .ZN(n6236) );
  AOI22_X1 U4941 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][10] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][10] ), .ZN(n6237) );
  AOI22_X1 U4942 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][10] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][10] ), .ZN(n6238) );
  OAI222_X1 U4943 ( .A1(n6240), .A2(n5468), .B1(n6241), .B2(n5525), .C1(n6129), 
        .C2(n5466), .ZN(n6239) );
  AOI21_X1 U4946 ( .B1(\UUT/Mcontrol/d_sampled_finstr [19]), .B2(n5932), .A(
        n7131), .ZN(n6243) );
  NAND2_X1 U4947 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1945 ), .A2(n7117), 
        .ZN(n5932) );
  INV_X1 U4948 ( .A(n5924), .ZN(n5926) );
  AOI21_X1 U4951 ( .B1(n6246), .B2(n6247), .A(n6248), .ZN(n6245) );
  INV_X1 U4953 ( .A(\UUT/Mcontrol/Nextpc_decoding/N260 ), .ZN(n6247) );
  INV_X1 U4957 ( .A(\UUT/Mcontrol/Nextpc_decoding/N248 ), .ZN(n6252) );
  INV_X1 U4961 ( .A(\UUT/Mcontrol/Nextpc_decoding/N242 ), .ZN(n6254) );
  AOI22_X1 U4963 ( .A1(n5436), .A2(\UUT/regfile/reg_out[19][31] ), .B1(n5437), 
        .B2(\UUT/regfile/reg_out[18][31] ), .ZN(n6257) );
  AOI22_X1 U4969 ( .A1(n5441), .A2(\UUT/regfile/reg_out[21][31] ), .B1(n5442), 
        .B2(\UUT/regfile/reg_out[20][31] ), .ZN(n6264) );
  NAND3_X1 U4972 ( .A1(n6259), .A2(\UUT/rs1_addr [2]), .A3(n6262), .ZN(n5439)
         );
  NAND4_X1 U4973 ( .A1(n6262), .A2(\UUT/rs1_addr [1]), .A3(\UUT/rs1_addr [0]), 
        .A4(\UUT/rs1_addr [2]), .ZN(n5438) );
  NOR2_X1 U4974 ( .A1(n6267), .A2(\UUT/rs1_addr [3]), .ZN(n6262) );
  AOI22_X1 U4975 ( .A1(n5446), .A2(\UUT/regfile/reg_out[25][31] ), .B1(n5447), 
        .B2(\UUT/regfile/reg_out[24][31] ), .ZN(n6268) );
  NAND3_X1 U4978 ( .A1(n6259), .A2(\UUT/rs1_addr [4]), .A3(n6271), .ZN(n5444)
         );
  AOI22_X1 U4980 ( .A1(n5451), .A2(\UUT/regfile/reg_out[29][31] ), .B1(n5452), 
        .B2(\UUT/regfile/reg_out[28][31] ), .ZN(n6272) );
  NOR2_X1 U4985 ( .A1(n6267), .A2(n7375), .ZN(n6270) );
  AOI22_X1 U4988 ( .A1(n5458), .A2(\UUT/regfile/reg_out[5][31] ), .B1(n5459), 
        .B2(\UUT/regfile/reg_out[4][31] ), .ZN(n6277) );
  NAND3_X1 U4991 ( .A1(\UUT/rs1_addr [2]), .A2(n6275), .A3(n6276), .ZN(n5456)
         );
  NAND3_X1 U4992 ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/rs1_addr [2]), .A3(n6274), 
        .ZN(n5455) );
  NOR3_X1 U5022 ( .A1(\UUT/Mpath/the_shift/N115 ), .A2(
        \UUT/Mpath/the_shift/N118 ), .A3(\UUT/Mpath/the_shift/N111 ), .ZN(
        n6282) );
  INV_X1 U5023 ( .A(\UUT/Mcontrol/Nextpc_decoding/N254 ), .ZN(n6249) );
  INV_X1 U5024 ( .A(\UUT/Mcontrol/Nextpc_decoding/N266 ), .ZN(n6244) );
  INV_X1 U5032 ( .A(\UUT/Mcontrol/Operation_decoding32/N1928 ), .ZN(n5937) );
  INV_X1 U5033 ( .A(\UUT/Mcontrol/Operation_decoding32/N1946 ), .ZN(n5917) );
  NOR2_X1 U5044 ( .A1(n7163), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .ZN(n5948) );
  OAI22_X1 U5045 ( .A1(n6285), .A2(n6286), .B1(n6287), .B2(n6288), .ZN(
        D_DATA_OUTBUS[9]) );
  OAI22_X1 U5046 ( .A1(n6286), .A2(n6289), .B1(n6287), .B2(n6290), .ZN(
        D_DATA_OUTBUS[8]) );
  OAI221_X1 U5047 ( .B1(n6291), .B2(n6292), .C1(n6286), .C2(n6293), .A(n6294), 
        .ZN(D_DATA_OUTBUS[31]) );
  NAND2_X1 U5048 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[31] ), .A2(n6295), 
        .ZN(n6294) );
  OAI221_X1 U5049 ( .B1(n6291), .B2(n6296), .C1(n6286), .C2(n6297), .A(n6298), 
        .ZN(D_DATA_OUTBUS[30]) );
  NAND2_X1 U5050 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[30] ), .A2(n6295), 
        .ZN(n6298) );
  OAI221_X1 U5051 ( .B1(n6291), .B2(n6299), .C1(n6286), .C2(n6300), .A(n6301), 
        .ZN(D_DATA_OUTBUS[29]) );
  NAND2_X1 U5052 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[29] ), .A2(n6295), 
        .ZN(n6301) );
  OAI221_X1 U5053 ( .B1(n6291), .B2(n6302), .C1(n6286), .C2(n6303), .A(n6304), 
        .ZN(D_DATA_OUTBUS[28]) );
  NAND2_X1 U5054 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[28] ), .A2(n6295), 
        .ZN(n6304) );
  OAI221_X1 U5055 ( .B1(n6291), .B2(n6305), .C1(n6286), .C2(n6306), .A(n6307), 
        .ZN(D_DATA_OUTBUS[27]) );
  NAND2_X1 U5056 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[27] ), .A2(n6295), 
        .ZN(n6307) );
  OAI221_X1 U5057 ( .B1(n6291), .B2(n6308), .C1(n6286), .C2(n6309), .A(n6310), 
        .ZN(D_DATA_OUTBUS[26]) );
  NAND2_X1 U5058 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[26] ), .A2(n6295), 
        .ZN(n6310) );
  OAI221_X1 U5059 ( .B1(n6288), .B2(n6291), .C1(n6285), .C2(n6286), .A(n6311), 
        .ZN(D_DATA_OUTBUS[25]) );
  NAND2_X1 U5060 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[25] ), .A2(n6295), 
        .ZN(n6311) );
  OAI221_X1 U5061 ( .B1(n6290), .B2(n6291), .C1(n6286), .C2(n6289), .A(n6312), 
        .ZN(D_DATA_OUTBUS[24]) );
  NAND2_X1 U5062 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[24] ), .A2(n6295), 
        .ZN(n6312) );
  OAI21_X1 U5063 ( .B1(n6313), .B2(n6293), .A(n6314), .ZN(D_DATA_OUTBUS[23])
         );
  NAND2_X1 U5064 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[23] ), .A2(n6295), 
        .ZN(n6314) );
  OAI21_X1 U5065 ( .B1(n6313), .B2(n6297), .A(n6315), .ZN(D_DATA_OUTBUS[22])
         );
  NAND2_X1 U5066 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[22] ), .A2(n6295), 
        .ZN(n6315) );
  OAI21_X1 U5067 ( .B1(n6313), .B2(n6300), .A(n6316), .ZN(D_DATA_OUTBUS[21])
         );
  NAND2_X1 U5068 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[21] ), .A2(n6295), 
        .ZN(n6316) );
  OAI21_X1 U5069 ( .B1(n6313), .B2(n6303), .A(n6317), .ZN(D_DATA_OUTBUS[20])
         );
  NAND2_X1 U5070 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[20] ), .A2(n6295), 
        .ZN(n6317) );
  OAI21_X1 U5071 ( .B1(n6313), .B2(n6306), .A(n6318), .ZN(D_DATA_OUTBUS[19])
         );
  NAND2_X1 U5072 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[19] ), .A2(n6295), 
        .ZN(n6318) );
  OAI21_X1 U5073 ( .B1(n6313), .B2(n6309), .A(n6319), .ZN(D_DATA_OUTBUS[18])
         );
  NAND2_X1 U5074 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[18] ), .A2(n6295), 
        .ZN(n6319) );
  OAI21_X1 U5075 ( .B1(n6313), .B2(n6285), .A(n6320), .ZN(D_DATA_OUTBUS[17])
         );
  NAND2_X1 U5076 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[17] ), .A2(n6295), 
        .ZN(n6320) );
  OAI21_X1 U5077 ( .B1(n6313), .B2(n6289), .A(n6321), .ZN(D_DATA_OUTBUS[16])
         );
  NAND2_X1 U5078 ( .A1(\UUT/Mpath/the_memhandle/smdr_out[16] ), .A2(n6295), 
        .ZN(n6321) );
  AND2_X1 U5079 ( .A1(dmem_isbyte), .A2(dmem_ishalf), .ZN(n6295) );
  AND2_X1 U5080 ( .A1(n6286), .A2(n6291), .ZN(n6313) );
  NAND2_X1 U5081 ( .A1(\UUT/Mpath/the_memhandle/N237 ), .A2(dmem_isbyte), .ZN(
        n6291) );
  OAI22_X1 U5082 ( .A1(n6286), .A2(n6293), .B1(n6287), .B2(n6292), .ZN(
        D_DATA_OUTBUS[15]) );
  OAI22_X1 U5083 ( .A1(n6286), .A2(n6297), .B1(n6287), .B2(n6296), .ZN(
        D_DATA_OUTBUS[14]) );
  OAI22_X1 U5084 ( .A1(n6286), .A2(n6300), .B1(n6287), .B2(n6299), .ZN(
        D_DATA_OUTBUS[13]) );
  OAI22_X1 U5085 ( .A1(n6286), .A2(n6303), .B1(n6287), .B2(n6302), .ZN(
        D_DATA_OUTBUS[12]) );
  OAI22_X1 U5086 ( .A1(n6286), .A2(n6306), .B1(n6287), .B2(n6305), .ZN(
        D_DATA_OUTBUS[11]) );
  OAI22_X1 U5087 ( .A1(n6286), .A2(n6309), .B1(n6287), .B2(n6308), .ZN(
        D_DATA_OUTBUS[10]) );
  INV_X1 U5088 ( .A(\UUT/Mpath/the_memhandle/N234 ), .ZN(n6286) );
  NOR2_X1 U5089 ( .A1(n6142), .A2(n6322), .ZN(D_ADDR_OUTBUS[9]) );
  INV_X1 U5090 ( .A(n6097), .ZN(n6142) );
  NOR2_X1 U5091 ( .A1(n6151), .A2(n6322), .ZN(D_ADDR_OUTBUS[8]) );
  INV_X1 U5092 ( .A(n6099), .ZN(n6151) );
  NOR2_X1 U5093 ( .A1(n6160), .A2(n6322), .ZN(D_ADDR_OUTBUS[7]) );
  INV_X1 U5094 ( .A(n6101), .ZN(n6160) );
  NOR2_X1 U5095 ( .A1(n6169), .A2(n6322), .ZN(D_ADDR_OUTBUS[6]) );
  INV_X1 U5096 ( .A(n6103), .ZN(n6169) );
  NOR2_X1 U5097 ( .A1(n6178), .A2(n6322), .ZN(D_ADDR_OUTBUS[5]) );
  INV_X1 U5098 ( .A(n6105), .ZN(n6178) );
  NOR2_X1 U5099 ( .A1(n6187), .A2(n6322), .ZN(D_ADDR_OUTBUS[4]) );
  INV_X1 U5100 ( .A(n6107), .ZN(n6187) );
  NOR2_X1 U5101 ( .A1(n6199), .A2(n6322), .ZN(D_ADDR_OUTBUS[3]) );
  INV_X1 U5102 ( .A(n6109), .ZN(n6199) );
  NOR2_X1 U5103 ( .A1(n6110), .A2(n6322), .ZN(D_ADDR_OUTBUS[31]) );
  NOR2_X1 U5104 ( .A1(n5467), .A2(n6322), .ZN(D_ADDR_OUTBUS[30]) );
  NOR2_X1 U5105 ( .A1(n6210), .A2(n6322), .ZN(D_ADDR_OUTBUS[2]) );
  INV_X1 U5106 ( .A(n6113), .ZN(n6210) );
  NOR2_X1 U5107 ( .A1(n5476), .A2(n6322), .ZN(D_ADDR_OUTBUS[29]) );
  NOR2_X1 U5108 ( .A1(n5484), .A2(n6322), .ZN(D_ADDR_OUTBUS[28]) );
  NOR2_X1 U5109 ( .A1(n5492), .A2(n6322), .ZN(D_ADDR_OUTBUS[27]) );
  NOR2_X1 U5110 ( .A1(n5500), .A2(n6322), .ZN(D_ADDR_OUTBUS[26]) );
  NOR2_X1 U5111 ( .A1(n5508), .A2(n6322), .ZN(D_ADDR_OUTBUS[25]) );
  NOR2_X1 U5112 ( .A1(n5516), .A2(n6322), .ZN(D_ADDR_OUTBUS[24]) );
  NOR2_X1 U5113 ( .A1(n5967), .A2(n6322), .ZN(D_ADDR_OUTBUS[23]) );
  INV_X1 U5114 ( .A(n6114), .ZN(n5967) );
  NOR2_X1 U5115 ( .A1(n5978), .A2(n6322), .ZN(D_ADDR_OUTBUS[22]) );
  INV_X1 U5116 ( .A(n6115), .ZN(n5978) );
  NOR2_X1 U5117 ( .A1(n5988), .A2(n6322), .ZN(D_ADDR_OUTBUS[21]) );
  INV_X1 U5118 ( .A(n6116), .ZN(n5988) );
  NOR2_X1 U5119 ( .A1(n5998), .A2(n6322), .ZN(D_ADDR_OUTBUS[20]) );
  INV_X1 U5120 ( .A(n6117), .ZN(n5998) );
  NOR2_X1 U5121 ( .A1(n5956), .A2(n6322), .ZN(D_ADDR_OUTBUS[1]) );
  INV_X1 U5122 ( .A(\UUT/daddr_out [1]), .ZN(n5956) );
  NOR2_X1 U5123 ( .A1(n6011), .A2(n6322), .ZN(D_ADDR_OUTBUS[19]) );
  INV_X1 U5124 ( .A(n6118), .ZN(n6011) );
  NOR2_X1 U5125 ( .A1(n6024), .A2(n6322), .ZN(D_ADDR_OUTBUS[18]) );
  INV_X1 U5126 ( .A(n6119), .ZN(n6024) );
  NOR2_X1 U5127 ( .A1(n6045), .A2(n6322), .ZN(D_ADDR_OUTBUS[17]) );
  INV_X1 U5128 ( .A(n6120), .ZN(n6045) );
  NOR2_X1 U5129 ( .A1(n6057), .A2(n6322), .ZN(D_ADDR_OUTBUS[16]) );
  INV_X1 U5130 ( .A(n6121), .ZN(n6057) );
  NOR2_X1 U5131 ( .A1(n6068), .A2(n6322), .ZN(D_ADDR_OUTBUS[15]) );
  INV_X1 U5132 ( .A(n6122), .ZN(n6068) );
  NOR2_X1 U5133 ( .A1(n6082), .A2(n6322), .ZN(D_ADDR_OUTBUS[14]) );
  INV_X1 U5134 ( .A(n6123), .ZN(n6082) );
  NOR2_X1 U5135 ( .A1(n6092), .A2(n6322), .ZN(D_ADDR_OUTBUS[13]) );
  INV_X1 U5136 ( .A(n6124), .ZN(n6092) );
  NOR2_X1 U5137 ( .A1(n6222), .A2(n6322), .ZN(D_ADDR_OUTBUS[12]) );
  INV_X1 U5138 ( .A(n6126), .ZN(n6222) );
  NOR2_X1 U5139 ( .A1(n6231), .A2(n6322), .ZN(D_ADDR_OUTBUS[11]) );
  INV_X1 U5140 ( .A(n6128), .ZN(n6231) );
  NOR2_X1 U5141 ( .A1(n6240), .A2(n6322), .ZN(D_ADDR_OUTBUS[10]) );
  INV_X1 U5142 ( .A(n6130), .ZN(n6240) );
  NAND2_X1 U5143 ( .A1(n6323), .A2(n6325), .ZN(n6324) );
  INV_X1 U5144 ( .A(\UUT/Mpath/the_alu/N492 ), .ZN(n6325) );
  NOR2_X1 U5145 ( .A1(n5523), .A2(n6322), .ZN(D_ADDR_OUTBUS[0]) );
  INV_X1 U5147 ( .A(\UUT/daddr_out [0]), .ZN(n5523) );
  OAI21_X1 U5148 ( .B1(\UUT/Mpath/the_alu/N492 ), .B2(n6327), .A(n6328), .ZN(
        n6326) );
  NAND2_X1 U5149 ( .A1(\UUT/Mpath/the_alu/N125 ), .A2(\UUT/Mpath/the_alu/N492 ), .ZN(n6328) );
  AOI22_X1 U5150 ( .A1(n6329), .A2(\UUT/Mpath/the_alu/N485 ), .B1(
        \UUT/Mpath/the_alu/N157 ), .B2(\UUT/Mpath/the_alu/N486 ), .ZN(n6327)
         );
  OAI21_X1 U5151 ( .B1(\UUT/Mpath/the_alu/N480 ), .B2(n6330), .A(n6331), .ZN(
        n6329) );
  NAND2_X1 U5152 ( .A1(\UUT/Mpath/the_alu/N189 ), .A2(\UUT/Mpath/the_alu/N480 ), .ZN(n6331) );
  AOI22_X1 U5153 ( .A1(\UUT/Mpath/the_alu/N221 ), .A2(\UUT/Mpath/the_alu/N474 ), .B1(\UUT/Mpath/the_alu/N473 ), .B2(\UUT/Mpath/out_regA[0] ), .ZN(n6330) );
  CLKBUF_X2 U5154 ( .A(dmem_ishalf), .Z(n6332) );
  CLKBUF_X2 U5155 ( .A(dmem_ishalf), .Z(n6333) );
  CLKBUF_X2 U5156 ( .A(dmem_ishalf), .Z(n6334) );
  CLKBUF_X2 U5157 ( .A(dmem_ishalf), .Z(n6335) );
  CLKBUF_X2 U5158 ( .A(D_ADDR_OUTBUS[1]), .Z(n6336) );
  CLKBUF_X2 U5159 ( .A(dmem_isbyte), .Z(n6337) );
  CLKBUF_X2 U5160 ( .A(dmem_isbyte), .Z(n6338) );
  CLKBUF_X2 U5161 ( .A(dmem_isbyte), .Z(N13) );
  CLKBUF_X2 U5162 ( .A(dmem_isbyte), .Z(N11) );
  CLKBUF_X2 U5163 ( .A(dmem_isbyte), .Z(N9) );
  CLKBUF_X2 U5164 ( .A(dmem_isbyte), .Z(N7) );
  CLKBUF_X2 U5165 ( .A(dmem_ishalf), .Z(N3) );
  CLKBUF_X2 U5166 ( .A(D_ADDR_OUTBUS[1]), .Z(N2) );
  CLKBUF_X2 U5167 ( .A(dmem_ishalf), .Z(N0) );
  INV_X2 U5168 ( .A(n6338), .ZN(N1) );
  INV_X2 U5169 ( .A(n6337), .ZN(N4) );
  INV_X2 U5170 ( .A(n6336), .ZN(N5) );
  INV_X2 U5171 ( .A(n6335), .ZN(N6) );
  INV_X2 U5172 ( .A(n6334), .ZN(N8) );
  INV_X2 U5173 ( .A(n6333), .ZN(N10) );
  INV_X2 U5174 ( .A(n6332), .ZN(N12) );
  ubus localbus ( .clk(CLK), .reset(\UUT/Mcontrol/int_reset ), .M1_BUSY(1'b1), 
        .M1_MR(dmem_read), .M1_MW(dmem_write), .M1_NREADY(\UUT/Mcontrol/N22 ), 
        .M1_ADDR_OUTBUS(D_ADDR_OUTBUS), .M1_DATA_INBUS(D_DATA_INBUS), 
        .M1_DATA_OUTBUS(D_DATA_OUTBUS), .S1_MR(dram_mr), .S1_MW(dram_mw), 
        .S1_NREADY(1'b1), .S1_ADDR_OUTBUS({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        \dram_addr_outbus[12] , \dram_addr_outbus[11] , \dram_addr_outbus[10] , 
        \dram_addr_outbus[9] , \dram_addr_outbus[8] , \dram_addr_outbus[7] , 
        \dram_addr_outbus[6] , \dram_addr_outbus[5] , \dram_addr_outbus[4] , 
        \dram_addr_outbus[3] , \dram_addr_outbus[2] , SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20}), .S1_DATA_INBUS({\dram_data_inbus[31] , 
        \dram_data_inbus[30] , \dram_data_inbus[29] , \dram_data_inbus[28] , 
        \dram_data_inbus[27] , \dram_data_inbus[26] , \dram_data_inbus[25] , 
        \dram_data_inbus[24] , \dram_data_inbus[23] , \dram_data_inbus[22] , 
        \dram_data_inbus[21] , \dram_data_inbus[20] , \dram_data_inbus[19] , 
        \dram_data_inbus[18] , \dram_data_inbus[17] , \dram_data_inbus[16] , 
        \dram_data_inbus[15] , \dram_data_inbus[14] , \dram_data_inbus[13] , 
        \dram_data_inbus[12] , \dram_data_inbus[11] , \dram_data_inbus[10] , 
        \dram_data_inbus[9] , \dram_data_inbus[8] , \dram_data_inbus[7] , 
        \dram_data_inbus[6] , \dram_data_inbus[5] , \dram_data_inbus[4] , 
        \dram_data_inbus[3] , \dram_data_inbus[2] , \dram_data_inbus[1] , 
        \dram_data_inbus[0] }), .S1_DATA_OUTBUS({\dram_data_outbus[31] , 
        \dram_data_outbus[30] , \dram_data_outbus[29] , \dram_data_outbus[28] , 
        \dram_data_outbus[27] , \dram_data_outbus[26] , \dram_data_outbus[25] , 
        \dram_data_outbus[24] , \dram_data_outbus[23] , \dram_data_outbus[22] , 
        \dram_data_outbus[21] , \dram_data_outbus[20] , \dram_data_outbus[19] , 
        \dram_data_outbus[18] , \dram_data_outbus[17] , \dram_data_outbus[16] , 
        \dram_data_outbus[15] , \dram_data_outbus[14] , \dram_data_outbus[13] , 
        \dram_data_outbus[12] , \dram_data_outbus[11] , \dram_data_outbus[10] , 
        \dram_data_outbus[9] , \dram_data_outbus[8] , \dram_data_outbus[7] , 
        \dram_data_outbus[6] , \dram_data_outbus[5] , \dram_data_outbus[4] , 
        \dram_data_outbus[3] , \dram_data_outbus[2] , \dram_data_outbus[1] , 
        \dram_data_outbus[0] }), .S2_BUSY(BUS_BUSY), .S2_MR(BUS_MR), .S2_MW(
        BUS_MW), .S2_NREADY(BUS_NREADY), .S2_ADDR_OUTBUS(BUS_ADDR_OUTBUS), 
        .S2_DATA_INBUS(BUS_DATA_INBUS), .S2_DATA_OUTBUS(BUS_DATA_OUTBUS), 
        .S3_NREADY(1'b1), .S3_DATA_INBUS({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .S4_NREADY(1'b1), .S4_DATA_INBUS({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  SRAM DMem ( .clk(CLK), .rdn(dram_mr), .wrn(dram_mw), .address({
        \dram_addr_outbus[12] , \dram_addr_outbus[11] , \dram_addr_outbus[10] , 
        \dram_addr_outbus[9] , \dram_addr_outbus[8] , \dram_addr_outbus[7] , 
        \dram_addr_outbus[6] , \dram_addr_outbus[5] , \dram_addr_outbus[4] , 
        \dram_addr_outbus[3] , \dram_addr_outbus[2] }), .bit_wen({d_select[31], 
        d_select[31], d_select[31], d_select[31], d_select[31], d_select[31], 
        d_select[31], d_select[31], d_select[23], d_select[23], d_select[23], 
        d_select[23], d_select[23], d_select[23], d_select[23], d_select[23], 
        d_select[9], d_select[9], d_select[9], d_select[9], d_select[9], 
        d_select[9], d_select[9], d_select[9], d_select[7], d_select[7], 
        d_select[7], d_select[7], d_select[7], d_select[7], d_select[7], 
        d_select[7]}), .data_in({\dram_data_outbus[31] , 
        \dram_data_outbus[30] , \dram_data_outbus[29] , \dram_data_outbus[28] , 
        \dram_data_outbus[27] , \dram_data_outbus[26] , \dram_data_outbus[25] , 
        \dram_data_outbus[24] , \dram_data_outbus[23] , \dram_data_outbus[22] , 
        \dram_data_outbus[21] , \dram_data_outbus[20] , \dram_data_outbus[19] , 
        \dram_data_outbus[18] , \dram_data_outbus[17] , \dram_data_outbus[16] , 
        \dram_data_outbus[15] , \dram_data_outbus[14] , \dram_data_outbus[13] , 
        \dram_data_outbus[12] , \dram_data_outbus[11] , \dram_data_outbus[10] , 
        \dram_data_outbus[9] , \dram_data_outbus[8] , \dram_data_outbus[7] , 
        \dram_data_outbus[6] , \dram_data_outbus[5] , \dram_data_outbus[4] , 
        \dram_data_outbus[3] , \dram_data_outbus[2] , \dram_data_outbus[1] , 
        \dram_data_outbus[0] }), .data_out({\dram_data_inbus[31] , 
        \dram_data_inbus[30] , \dram_data_inbus[29] , \dram_data_inbus[28] , 
        \dram_data_inbus[27] , \dram_data_inbus[26] , \dram_data_inbus[25] , 
        \dram_data_inbus[24] , \dram_data_inbus[23] , \dram_data_inbus[22] , 
        \dram_data_inbus[21] , \dram_data_inbus[20] , \dram_data_inbus[19] , 
        \dram_data_inbus[18] , \dram_data_inbus[17] , \dram_data_inbus[16] , 
        \dram_data_inbus[15] , \dram_data_inbus[14] , \dram_data_inbus[13] , 
        \dram_data_inbus[12] , \dram_data_inbus[11] , \dram_data_inbus[10] , 
        \dram_data_inbus[9] , \dram_data_inbus[8] , \dram_data_inbus[7] , 
        \dram_data_inbus[6] , \dram_data_inbus[5] , \dram_data_inbus[4] , 
        \dram_data_inbus[3] , \dram_data_inbus[2] , \dram_data_inbus[1] , 
        \dram_data_inbus[0] }) );
  SRAM IMem ( .clk(CLK), .rdn(iram_rd), .wrn(1'b1), .address({
        \UUT/Mcontrol/Program_counter/N28 , \UUT/Mcontrol/Program_counter/N26 , 
        \UUT/Mcontrol/Program_counter/N24 , \UUT/Mcontrol/Program_counter/N22 , 
        \UUT/Mcontrol/Program_counter/N20 , \UUT/Mcontrol/Program_counter/N18 , 
        \UUT/Mcontrol/Program_counter/N16 , \UUT/Mcontrol/Program_counter/N14 , 
        \UUT/Mcontrol/Program_counter/N12 , \UUT/Mcontrol/Program_counter/N10 , 
        \UUT/Mcontrol/Program_counter/N8 }), .bit_wen({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .data_out(I_DATA_INBUS) );
  up_island_DW01_add_1 \UUT/Mcontrol/Nextpc_decoding/bta_calc/add_391  ( .A({
        1'b0, \UUT/Mcontrol/f_currpc }), .B({1'b0, \UUT/break_code[23] , 
        \UUT/break_code[22] , \UUT/break_code[21] , \UUT/break_code[20] , 
        \UUT/break_code[19] , \UUT/break_code[18] , \UUT/break_code[17] , 
        \UUT/break_code[16] , \UUT/break_code[15] , \UUT/break_code[14] , 
        \UUT/break_code[13] , \UUT/break_code[12] , \UUT/break_code[11] , 
        \UUT/break_code[10] , \UUT/break_code[9] , \UUT/break_code[8] , 
        \UUT/break_code[7] , \UUT/break_code[6] , \UUT/break_code[5] , 
        \UUT/break_code[4] , n7174, n7238, \UUT/break_code[1] , 
        \UUT/break_code[0] }), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__21, 
        \UUT/Mcontrol/Nextpc_decoding/Bta }) );
  up_island_DW01_add_2 \UUT/Mcontrol/Nextpc_decoding/incr/add_391  ( .A({1'b0, 
        \UUT/Mcontrol/f_currpc }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, \UUT/jar_in }) );
  up_island_DW01_sub_1 \UUT/Mpath/the_alu/sub_96  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , n1265, n1261, \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , n1245, 
        \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[11] , n1219, n7196, 
        \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[7] , 
        \UUT/Mpath/out_regA[6] , n1321, \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .B({
        \UUT/Mpath/out_regB[31] , \UUT/Mpath/out_regB[30] , 
        \UUT/Mpath/out_regB[29] , \UUT/Mpath/out_regB[28] , 
        \UUT/Mpath/out_regB[27] , \UUT/Mpath/out_regB[26] , 
        \UUT/Mpath/out_regB[25] , \UUT/Mpath/out_regB[24] , 
        \UUT/Mpath/out_regB[23] , \UUT/Mpath/out_regB[22] , 
        \UUT/Mpath/out_regB[21] , n7094, \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n7400, n7401, n7404, 
        n7406, n7408}), .DIFF({\UUT/Mpath/the_alu/diff[31] , 
        \UUT/Mpath/the_alu/diff[30] , \UUT/Mpath/the_alu/diff[29] , 
        \UUT/Mpath/the_alu/diff[28] , \UUT/Mpath/the_alu/diff[27] , 
        \UUT/Mpath/the_alu/diff[26] , \UUT/Mpath/the_alu/diff[25] , 
        \UUT/Mpath/the_alu/diff[24] , \UUT/Mpath/the_alu/diff[23] , 
        \UUT/Mpath/the_alu/diff[22] , \UUT/Mpath/the_alu/diff[21] , 
        \UUT/Mpath/the_alu/diff[20] , \UUT/Mpath/the_alu/diff[19] , 
        \UUT/Mpath/the_alu/diff[18] , \UUT/Mpath/the_alu/diff[17] , 
        \UUT/Mpath/the_alu/diff[16] , \UUT/Mpath/the_alu/diff[15] , 
        \UUT/Mpath/the_alu/diff[14] , \UUT/Mpath/the_alu/diff[13] , 
        \UUT/Mpath/the_alu/diff[12] , \UUT/Mpath/the_alu/diff[11] , 
        \UUT/Mpath/the_alu/diff[10] , \UUT/Mpath/the_alu/diff[9] , 
        \UUT/Mpath/the_alu/diff[8] , \UUT/Mpath/the_alu/diff[7] , 
        \UUT/Mpath/the_alu/diff[6] , \UUT/Mpath/the_alu/diff[5] , 
        \UUT/Mpath/the_alu/diff[4] , \UUT/Mpath/the_alu/diff[3] , 
        \UUT/Mpath/the_alu/diff[2] , \UUT/Mpath/the_alu/diff[1] , 
        \UUT/Mpath/the_alu/diff[0] }), .CI(1'b0) );
  up_island_DW_mult_tc_1 \UUT/Mpath/the_mult/mult_186  ( .a({
        \UUT/Mpath/the_mult/x_operand1[31] , 
        \UUT/Mpath/the_mult/x_operand1[30] , 
        \UUT/Mpath/the_mult/x_operand1[29] , 
        \UUT/Mpath/the_mult/x_operand1[28] , 
        \UUT/Mpath/the_mult/x_operand1[27] , 
        \UUT/Mpath/the_mult/x_operand1[26] , 
        \UUT/Mpath/the_mult/x_operand1[25] , 
        \UUT/Mpath/the_mult/x_operand1[24] , 
        \UUT/Mpath/the_mult/x_operand1[23] , 
        \UUT/Mpath/the_mult/x_operand1[22] , 
        \UUT/Mpath/the_mult/x_operand1[21] , 
        \UUT/Mpath/the_mult/x_operand1[20] , 
        \UUT/Mpath/the_mult/x_operand1[19] , 
        \UUT/Mpath/the_mult/x_operand1[18] , 
        \UUT/Mpath/the_mult/x_operand1[17] , 
        \UUT/Mpath/the_mult/x_operand1[16] , 
        \UUT/Mpath/the_mult/x_operand1[15] , 
        \UUT/Mpath/the_mult/x_operand1[14] , 
        \UUT/Mpath/the_mult/x_operand1[13] , 
        \UUT/Mpath/the_mult/x_operand1[12] , 
        \UUT/Mpath/the_mult/x_operand1[11] , 
        \UUT/Mpath/the_mult/x_operand1[10] , 
        \UUT/Mpath/the_mult/x_operand1[9] , \UUT/Mpath/the_mult/x_operand1[8] , 
        \UUT/Mpath/the_mult/x_operand1[7] , \UUT/Mpath/the_mult/x_operand1[6] , 
        \UUT/Mpath/the_mult/x_operand1[5] , \UUT/Mpath/the_mult/x_operand1[4] , 
        \UUT/Mpath/the_mult/x_operand1[3] , \UUT/Mpath/the_mult/x_operand1[2] , 
        \UUT/Mpath/the_mult/x_operand1[1] , \UUT/Mpath/the_mult/x_operand1[0] }), .b({n6359, \UUT/Mpath/the_mult/x_operand2 [30:28], n6973, 
        \UUT/Mpath/the_mult/x_operand2 [26], n6963, 
        \UUT/Mpath/the_mult/x_operand2 [24], n7048, 
        \UUT/Mpath/the_mult/x_operand2 [22], n7053, 
        \UUT/Mpath/the_mult/x_operand2 [20], n6938, 
        \UUT/Mpath/the_mult/x_operand2 [18], n6915, 
        \UUT/Mpath/the_mult/x_operand2 [16], n6842, 
        \UUT/Mpath/the_mult/x_operand2 [14], n7006, 
        \UUT/Mpath/the_mult/x_operand2 [12], n7058, 
        \UUT/Mpath/the_mult/x_operand2 [10], n7032, 
        \UUT/Mpath/the_mult/x_operand2 [8], n6965, 
        \UUT/Mpath/the_mult/x_operand2 [6], n7080, 
        \UUT/Mpath/the_mult/x_operand2 [4], n7066, 
        \UUT/Mpath/the_mult/x_operand2 [2:0]}), .product({
        \UUT/Mpath/the_mult/x_mult_out[63] , 
        \UUT/Mpath/the_mult/x_mult_out[62] , 
        \UUT/Mpath/the_mult/x_mult_out[61] , 
        \UUT/Mpath/the_mult/x_mult_out[60] , 
        \UUT/Mpath/the_mult/x_mult_out[59] , 
        \UUT/Mpath/the_mult/x_mult_out[58] , 
        \UUT/Mpath/the_mult/x_mult_out[57] , 
        \UUT/Mpath/the_mult/x_mult_out[56] , 
        \UUT/Mpath/the_mult/x_mult_out[55] , 
        \UUT/Mpath/the_mult/x_mult_out[54] , 
        \UUT/Mpath/the_mult/x_mult_out[53] , 
        \UUT/Mpath/the_mult/x_mult_out[52] , 
        \UUT/Mpath/the_mult/x_mult_out[51] , 
        \UUT/Mpath/the_mult/x_mult_out[50] , 
        \UUT/Mpath/the_mult/x_mult_out[49] , 
        \UUT/Mpath/the_mult/x_mult_out[48] , 
        \UUT/Mpath/the_mult/x_mult_out[47] , 
        \UUT/Mpath/the_mult/x_mult_out[46] , 
        \UUT/Mpath/the_mult/x_mult_out[45] , 
        \UUT/Mpath/the_mult/x_mult_out[44] , 
        \UUT/Mpath/the_mult/x_mult_out[43] , 
        \UUT/Mpath/the_mult/x_mult_out[42] , 
        \UUT/Mpath/the_mult/x_mult_out[41] , 
        \UUT/Mpath/the_mult/x_mult_out[40] , 
        \UUT/Mpath/the_mult/x_mult_out[39] , 
        \UUT/Mpath/the_mult/x_mult_out[38] , 
        \UUT/Mpath/the_mult/x_mult_out[37] , 
        \UUT/Mpath/the_mult/x_mult_out[36] , 
        \UUT/Mpath/the_mult/x_mult_out[35] , 
        \UUT/Mpath/the_mult/x_mult_out[34] , 
        \UUT/Mpath/the_mult/x_mult_out[33] , 
        \UUT/Mpath/the_mult/x_mult_out[32] , 
        \UUT/Mpath/the_mult/x_mult_out[31] , 
        \UUT/Mpath/the_mult/x_mult_out[30] , 
        \UUT/Mpath/the_mult/x_mult_out[29] , 
        \UUT/Mpath/the_mult/x_mult_out[28] , 
        \UUT/Mpath/the_mult/x_mult_out[27] , 
        \UUT/Mpath/the_mult/x_mult_out[26] , 
        \UUT/Mpath/the_mult/x_mult_out[25] , 
        \UUT/Mpath/the_mult/x_mult_out[24] , 
        \UUT/Mpath/the_mult/x_mult_out[23] , 
        \UUT/Mpath/the_mult/x_mult_out[22] , 
        \UUT/Mpath/the_mult/x_mult_out[21] , 
        \UUT/Mpath/the_mult/x_mult_out[20] , 
        \UUT/Mpath/the_mult/x_mult_out[19] , 
        \UUT/Mpath/the_mult/x_mult_out[18] , 
        \UUT/Mpath/the_mult/x_mult_out[17] , 
        \UUT/Mpath/the_mult/x_mult_out[16] , 
        \UUT/Mpath/the_mult/x_mult_out[15] , 
        \UUT/Mpath/the_mult/x_mult_out[14] , 
        \UUT/Mpath/the_mult/x_mult_out[13] , 
        \UUT/Mpath/the_mult/x_mult_out[12] , 
        \UUT/Mpath/the_mult/x_mult_out[11] , 
        \UUT/Mpath/the_mult/x_mult_out[10] , 
        \UUT/Mpath/the_mult/x_mult_out[9] , \UUT/Mpath/the_mult/x_mult_out[8] , 
        \UUT/Mpath/the_mult/x_mult_out[7] , \UUT/Mpath/the_mult/x_mult_out[6] , 
        \UUT/Mpath/the_mult/x_mult_out[5] , \UUT/Mpath/the_mult/x_mult_out[4] , 
        \UUT/Mpath/the_mult/x_mult_out[3] , \UUT/Mpath/the_mult/x_mult_out[2] , 
        \UUT/Mpath/the_mult/x_mult_out[1] , \UUT/Mpath/the_mult/x_mult_out[0] }) );
  up_island_DW01_add_4 \UUT/Mpath/the_alu/add_95  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , n1265, n1261, \UUT/Mpath/out_regA[16] , 
        \UUT/Mpath/out_regA[15] , \UUT/Mpath/out_regA[14] , n1245, 
        \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[11] , n1219, n7196, 
        \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[7] , 
        \UUT/Mpath/out_regA[6] , \UUT/Mpath/out_regA[5] , 
        \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[3] , 
        \UUT/Mpath/out_regA[2] , \UUT/Mpath/out_regA[1] , 
        \UUT/Mpath/out_regA[0] }), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , 
        \UUT/Mpath/out_regB[20] , \UUT/Mpath/out_regB[19] , 
        \UUT/Mpath/out_regB[18] , \UUT/Mpath/out_regB[17] , 
        \UUT/Mpath/out_regB[16] , \UUT/Mpath/out_regB[15] , 
        \UUT/Mpath/out_regB[14] , \UUT/Mpath/out_regB[13] , 
        \UUT/Mpath/out_regB[12] , \UUT/Mpath/out_regB[11] , 
        \UUT/Mpath/out_regB[10] , \UUT/Mpath/out_regB[9] , 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , 
        \UUT/Mpath/out_regB[6] , \UUT/Mpath/out_regB[5] , n7399, n7401, n7403, 
        n7405, n7408}), .SUM({\UUT/Mpath/the_alu/sum[31] , 
        \UUT/Mpath/the_alu/sum[30] , \UUT/Mpath/the_alu/sum[29] , 
        \UUT/Mpath/the_alu/sum[28] , \UUT/Mpath/the_alu/sum[27] , 
        \UUT/Mpath/the_alu/sum[26] , \UUT/Mpath/the_alu/sum[25] , 
        \UUT/Mpath/the_alu/sum[24] , \UUT/Mpath/the_alu/sum[23] , 
        \UUT/Mpath/the_alu/sum[22] , \UUT/Mpath/the_alu/sum[21] , 
        \UUT/Mpath/the_alu/sum[20] , \UUT/Mpath/the_alu/sum[19] , 
        \UUT/Mpath/the_alu/sum[18] , \UUT/Mpath/the_alu/sum[17] , 
        \UUT/Mpath/the_alu/sum[16] , \UUT/Mpath/the_alu/sum[15] , 
        \UUT/Mpath/the_alu/sum[14] , \UUT/Mpath/the_alu/sum[13] , 
        \UUT/Mpath/the_alu/sum[12] , \UUT/Mpath/the_alu/sum[11] , 
        \UUT/Mpath/the_alu/sum[10] , \UUT/Mpath/the_alu/sum[9] , 
        \UUT/Mpath/the_alu/sum[8] , \UUT/Mpath/the_alu/sum[7] , 
        \UUT/Mpath/the_alu/sum[6] , \UUT/Mpath/the_alu/sum[5] , 
        \UUT/Mpath/the_alu/sum[4] , \UUT/Mpath/the_alu/sum[3] , 
        \UUT/Mpath/the_alu/sum[2] , \UUT/Mpath/the_alu/sum[1] , 
        \UUT/Mpath/the_alu/sum[0] }), .CI(1'b0) );
  up_island_DW01_add_3 \UUT/Mpath/the_mult/accumulate/add_391  ( .A({1'b0, 
        \UUT/Mpath/the_mult/acc_out[63] , \UUT/Mpath/the_mult/acc_out[62] , 
        \UUT/Mpath/the_mult/acc_out[61] , \UUT/Mpath/the_mult/acc_out[60] , 
        \UUT/Mpath/the_mult/acc_out[59] , \UUT/Mpath/the_mult/acc_out[58] , 
        \UUT/Mpath/the_mult/acc_out[57] , \UUT/Mpath/the_mult/acc_out[56] , 
        \UUT/Mpath/the_mult/acc_out[55] , \UUT/Mpath/the_mult/acc_out[54] , 
        \UUT/Mpath/the_mult/acc_out[53] , \UUT/Mpath/the_mult/acc_out[52] , 
        \UUT/Mpath/the_mult/acc_out[51] , \UUT/Mpath/the_mult/acc_out[50] , 
        \UUT/Mpath/the_mult/acc_out[49] , \UUT/Mpath/the_mult/acc_out[48] , 
        \UUT/Mpath/the_mult/acc_out[47] , \UUT/Mpath/the_mult/acc_out[46] , 
        \UUT/Mpath/the_mult/acc_out[45] , \UUT/Mpath/the_mult/acc_out[44] , 
        \UUT/Mpath/the_mult/acc_out[43] , \UUT/Mpath/the_mult/acc_out[42] , 
        \UUT/Mpath/the_mult/acc_out[41] , \UUT/Mpath/the_mult/acc_out[40] , 
        \UUT/Mpath/the_mult/acc_out[39] , \UUT/Mpath/the_mult/acc_out[38] , 
        \UUT/Mpath/the_mult/acc_out[37] , \UUT/Mpath/the_mult/acc_out[36] , 
        \UUT/Mpath/the_mult/acc_out[35] , \UUT/Mpath/the_mult/acc_out[34] , 
        \UUT/Mpath/the_mult/acc_out[33] , \UUT/Mpath/the_mult/acc_out[32] , 
        \UUT/Mpath/the_mult/acc_out[31] , \UUT/Mpath/the_mult/acc_out[30] , 
        \UUT/Mpath/the_mult/acc_out[29] , \UUT/Mpath/the_mult/acc_out[28] , 
        \UUT/Mpath/the_mult/acc_out[27] , \UUT/Mpath/the_mult/acc_out[26] , 
        \UUT/Mpath/the_mult/acc_out[25] , \UUT/Mpath/the_mult/acc_out[24] , 
        \UUT/Mpath/the_mult/acc_out[23] , \UUT/Mpath/the_mult/acc_out[22] , 
        \UUT/Mpath/the_mult/acc_out[21] , \UUT/Mpath/the_mult/acc_out[20] , 
        \UUT/Mpath/the_mult/acc_out[19] , \UUT/Mpath/the_mult/acc_out[18] , 
        \UUT/Mpath/the_mult/acc_out[17] , \UUT/Mpath/the_mult/acc_out[16] , 
        \UUT/Mpath/the_mult/acc_out[15] , \UUT/Mpath/the_mult/acc_out[14] , 
        \UUT/Mpath/the_mult/acc_out[13] , \UUT/Mpath/the_mult/acc_out[12] , 
        \UUT/Mpath/the_mult/acc_out[11] , \UUT/Mpath/the_mult/acc_out[10] , 
        \UUT/Mpath/the_mult/acc_out[9] , \UUT/Mpath/the_mult/acc_out[8] , 
        \UUT/Mpath/the_mult/acc_out[7] , \UUT/Mpath/the_mult/acc_out[6] , 
        \UUT/Mpath/the_mult/acc_out[5] , \UUT/Mpath/the_mult/acc_out[4] , 
        \UUT/Mpath/the_mult/acc_out[3] , \UUT/Mpath/the_mult/acc_out[2] , 
        \UUT/Mpath/the_mult/acc_out[1] , \UUT/Mpath/the_mult/acc_out[0] }), 
        .B({1'b0, \UUT/Mpath/the_mult/Mult_out[63] , 
        \UUT/Mpath/the_mult/Mult_out[62] , \UUT/Mpath/the_mult/Mult_out[61] , 
        \UUT/Mpath/the_mult/Mult_out[60] , \UUT/Mpath/the_mult/Mult_out[59] , 
        \UUT/Mpath/the_mult/Mult_out[58] , \UUT/Mpath/the_mult/Mult_out[57] , 
        \UUT/Mpath/the_mult/Mult_out[56] , \UUT/Mpath/the_mult/Mult_out[55] , 
        \UUT/Mpath/the_mult/Mult_out[54] , \UUT/Mpath/the_mult/Mult_out[53] , 
        \UUT/Mpath/the_mult/Mult_out[52] , \UUT/Mpath/the_mult/Mult_out[51] , 
        \UUT/Mpath/the_mult/Mult_out[50] , \UUT/Mpath/the_mult/Mult_out[49] , 
        \UUT/Mpath/the_mult/Mult_out[48] , \UUT/Mpath/the_mult/Mult_out[47] , 
        \UUT/Mpath/the_mult/Mult_out[46] , \UUT/Mpath/the_mult/Mult_out[45] , 
        \UUT/Mpath/the_mult/Mult_out[44] , \UUT/Mpath/the_mult/Mult_out[43] , 
        \UUT/Mpath/the_mult/Mult_out[42] , \UUT/Mpath/the_mult/Mult_out[41] , 
        \UUT/Mpath/the_mult/Mult_out[40] , \UUT/Mpath/the_mult/Mult_out[39] , 
        \UUT/Mpath/the_mult/Mult_out[38] , \UUT/Mpath/the_mult/Mult_out[37] , 
        \UUT/Mpath/the_mult/Mult_out[36] , \UUT/Mpath/the_mult/Mult_out[35] , 
        \UUT/Mpath/the_mult/Mult_out[34] , \UUT/Mpath/the_mult/Mult_out[33] , 
        \UUT/Mpath/the_mult/Mult_out[32] , \UUT/Mpath/the_mult/Mult_out[31] , 
        \UUT/Mpath/the_mult/Mult_out[30] , \UUT/Mpath/the_mult/Mult_out[29] , 
        \UUT/Mpath/the_mult/Mult_out[28] , \UUT/Mpath/the_mult/Mult_out[27] , 
        \UUT/Mpath/the_mult/Mult_out[26] , \UUT/Mpath/the_mult/Mult_out[25] , 
        \UUT/Mpath/the_mult/Mult_out[24] , \UUT/Mpath/the_mult/Mult_out[23] , 
        \UUT/Mpath/the_mult/Mult_out[22] , \UUT/Mpath/the_mult/Mult_out[21] , 
        \UUT/Mpath/the_mult/Mult_out[20] , \UUT/Mpath/the_mult/Mult_out[19] , 
        \UUT/Mpath/the_mult/Mult_out[18] , \UUT/Mpath/the_mult/Mult_out[17] , 
        \UUT/Mpath/the_mult/Mult_out[16] , \UUT/Mpath/the_mult/Mult_out[15] , 
        \UUT/Mpath/the_mult/Mult_out[14] , \UUT/Mpath/the_mult/Mult_out[13] , 
        \UUT/Mpath/the_mult/Mult_out[12] , \UUT/Mpath/the_mult/Mult_out[11] , 
        \UUT/Mpath/the_mult/Mult_out[10] , \UUT/Mpath/the_mult/Mult_out[9] , 
        \UUT/Mpath/the_mult/Mult_out[8] , \UUT/Mpath/the_mult/Mult_out[7] , 
        \UUT/Mpath/the_mult/Mult_out[6] , \UUT/Mpath/the_mult/Mult_out[5] , 
        \UUT/Mpath/the_mult/Mult_out[4] , \UUT/Mpath/the_mult/Mult_out[3] , 
        \UUT/Mpath/the_mult/Mult_out[2] , \UUT/Mpath/the_mult/Mult_out[1] , 
        \UUT/Mpath/the_mult/Mult_out[0] }), .SUM({SYNOPSYS_UNCONNECTED__23, 
        \UUT/Mpath/the_mult/Mad_out }), .CI(1'b0) );
  up_island_DW_rightsh_1 \UUT/Mpath/the_shift/S_SRL/srl_128  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , n7138, n7167, n1265, 
        \UUT/Mpath/out_regA[17] , n7129, n7112, n7113, n1245, n7141, n7198, 
        \UUT/Mpath/out_regA[10] , n7132, n7189, \UUT/Mpath/out_regA[7] , n7106, 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .SH({n7399, n7401, 
        n7404, n7406, n7407}), .B(\UUT/Mpath/the_shift/sh_srl ), .DATA_TC(1'b0) );
  up_island_DW_sra_1 \UUT/Mpath/the_shift/S_SRA/sra_106  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , n7138, n7167, \UUT/Mpath/out_regA[18] , 
        \UUT/Mpath/out_regA[17] , n7129, n7112, n7113, n1245, n7141, n7198, 
        \UUT/Mpath/out_regA[10] , n7132, n7189, \UUT/Mpath/out_regA[7] , n7106, 
        \UUT/Mpath/out_regA[5] , \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .SH({n7399, n7401, 
        n7402, n7405, n7408}), .B(\UUT/Mpath/the_shift/sh_sra ), .SH_TC(1'b0)
         );
  up_island_DW_rbsh_1 \UUT/Mpath/the_shift/S_ROR/ror_81  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , \UUT/Mpath/out_regA[20] , 
        \UUT/Mpath/out_regA[19] , n1265, n1261, n7129, n7112, n7113, n1245, 
        \UUT/Mpath/out_regA[12] , \UUT/Mpath/out_regA[11] , n1219, n7132, 
        \UUT/Mpath/out_regA[8] , \UUT/Mpath/out_regA[7] , 
        \UUT/Mpath/out_regA[6] , n1321, \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .SH({n7399, n7401, 
        n7403, n7405, n7407}), .B(\UUT/Mpath/the_shift/sh_ror ), .SH_TC(1'b0)
         );
  up_island_DW01_bsh_1 \UUT/Mpath/the_shift/S_ROL/rol_55  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , n7138, n7167, n1265, n1261, n7129, n7112, 
        n7113, n1245, n7141, n7198, \UUT/Mpath/out_regA[10] , n7132, n7189, 
        \UUT/Mpath/out_regA[7] , n7106, n1321, \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .SH({n7399, n7401, 
        n7402, n7405, n7407}), .B(\UUT/Mpath/the_shift/sh_rol ) );
  up_island_DW_leftsh_1 \UUT/Mpath/the_shift/S_SLL/sll_150  ( .A({
        \UUT/Mpath/out_regA[31] , \UUT/Mpath/out_regA[30] , 
        \UUT/Mpath/out_regA[29] , \UUT/Mpath/out_regA[28] , 
        \UUT/Mpath/out_regA[27] , \UUT/Mpath/out_regA[26] , 
        \UUT/Mpath/out_regA[25] , \UUT/Mpath/out_regA[24] , 
        \UUT/Mpath/out_regA[23] , \UUT/Mpath/out_regA[22] , 
        \UUT/Mpath/out_regA[21] , n7138, n7167, n1265, 
        \UUT/Mpath/out_regA[17] , n7129, n7112, n7113, n1245, n7141, 
        \UUT/Mpath/out_regA[11] , n1219, n7132, \UUT/Mpath/out_regA[8] , 
        \UUT/Mpath/out_regA[7] , n7106, n1321, \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .SH({n7400, n7401, 
        n7404, n7405, n7407}), .B(\UUT/Mpath/the_shift/sh_sll ) );
  up_island_DW_cmp_0 \UUT/Mpath/the_alu/lt_114  ( .A({\UUT/Mpath/out_regA[31] , 
        \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[29] , 
        \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[27] , 
        \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[25] , 
        \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[23] , 
        \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[21] , n7138, n7167, 
        \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[17] , n7129, n7112, 
        n7113, n1245, n7193, n7198, \UUT/Mpath/out_regA[10] , n7132, n7189, 
        \UUT/Mpath/out_regA[7] , n7106, n1321, \UUT/Mpath/out_regA[4] , 
        \UUT/Mpath/out_regA[3] , \UUT/Mpath/out_regA[2] , 
        \UUT/Mpath/out_regA[1] , \UUT/Mpath/out_regA[0] }), .B({
        \UUT/Mpath/out_regB[31] , \UUT/Mpath/out_regB[30] , 
        \UUT/Mpath/out_regB[29] , \UUT/Mpath/out_regB[28] , 
        \UUT/Mpath/out_regB[27] , \UUT/Mpath/out_regB[26] , 
        \UUT/Mpath/out_regB[25] , \UUT/Mpath/out_regB[24] , 
        \UUT/Mpath/out_regB[23] , \UUT/Mpath/out_regB[22] , 
        \UUT/Mpath/out_regB[21] , n7194, n7190, n7135, n7197, n7136, n7125, 
        n7140, n7122, n7134, n7107, n7137, n7128, \UUT/Mpath/out_regB[8] , 
        \UUT/Mpath/out_regB[7] , n7099, n7114, n7399, n7401, n7403, n7405, 
        n7408}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(
        \UUT/Mpath/the_alu/N91 ) );
  up_island_DW_cmp_1 \UUT/Mpath/the_alu/lt_120  ( .A({\UUT/Mpath/out_regA[31] , 
        \UUT/Mpath/out_regA[30] , \UUT/Mpath/out_regA[29] , 
        \UUT/Mpath/out_regA[28] , \UUT/Mpath/out_regA[27] , 
        \UUT/Mpath/out_regA[26] , \UUT/Mpath/out_regA[25] , 
        \UUT/Mpath/out_regA[24] , \UUT/Mpath/out_regA[23] , 
        \UUT/Mpath/out_regA[22] , \UUT/Mpath/out_regA[21] , n7138, n7167, 
        \UUT/Mpath/out_regA[18] , \UUT/Mpath/out_regA[17] , n7129, n7112, 
        n7113, n1245, n7193, n7198, \UUT/Mpath/out_regA[10] , n7132, n7189, 
        \UUT/Mpath/out_regA[7] , n7106, \UUT/Mpath/out_regA[5] , 
        \UUT/Mpath/out_regA[4] , \UUT/Mpath/out_regA[3] , 
        \UUT/Mpath/out_regA[2] , \UUT/Mpath/out_regA[1] , 
        \UUT/Mpath/out_regA[0] }), .B({\UUT/Mpath/out_regB[31] , 
        \UUT/Mpath/out_regB[30] , \UUT/Mpath/out_regB[29] , 
        \UUT/Mpath/out_regB[28] , \UUT/Mpath/out_regB[27] , 
        \UUT/Mpath/out_regB[26] , \UUT/Mpath/out_regB[25] , 
        \UUT/Mpath/out_regB[24] , \UUT/Mpath/out_regB[23] , 
        \UUT/Mpath/out_regB[22] , \UUT/Mpath/out_regB[21] , n7194, n7190, 
        n7135, n7197, n7136, n7125, n7140, n7122, n7134, n7107, n7137, n7128, 
        \UUT/Mpath/out_regB[8] , \UUT/Mpath/out_regB[7] , n7099, n7114, n7399, 
        n7401, n7403, n7405, n7408}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(\UUT/Mpath/the_alu/N93 ) );
  up_island_DW01_cmp6_1 r723 ( .A({n7303, n7324, n7178, n7166, 
        \UUT/branch_rega [27:21], n7267, \UUT/branch_rega [19:0]}), .B(
        \UUT/branch_regb ), .TC(1'b0), .EQ(\UUT/Mcontrol/Nextpc_decoding/N22 ), 
        .NE(\UUT/Mcontrol/Nextpc_decoding/N25 ) );
  DFFR_X2 \UUT/Mcontrol/ir_fd/data_out_reg[26]  ( .D(n4239), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [26]), .QN(n2763)
         );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[7]  ( .D(n3546), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[7] ), .QN(
        \UUT/Mpath/the_alu/N69 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[0]  ( .D(n3785), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[0] ), .QN(
        \UUT/Mpath/the_alu/N83 ) );
  DFFR_X2 \UUT/Mpath/the_mult/multb/data_out_reg[1]  ( .D(n3779), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [1])
         );
  DFFR_X2 \UUT/Mpath/the_mult/multb/data_out_reg[29]  ( .D(n2873), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [29])
         );
  DFFS_X2 \UUT/Mcontrol/Program_counter/out_pc_reg[9]  ( .D(n4166), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [9]), .QN(
        n2712) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[2]  ( .D(n3746), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[2] ), .QN(
        \UUT/Mpath/the_alu/N79 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[17]  ( .D(n3148), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[17] ), .QN(
        \UUT/Mpath/the_alu/N49 ) );
  DFFR_X2 \UUT/Mpath/regA/data_out_reg[29]  ( .D(n4121), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[29] ), .QN(
        \UUT/Mpath/the_alu/N25 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[5]  ( .D(n3626), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[5] ), .QN(
        \UUT/Mpath/the_alu/N73 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[11]  ( .D(n3388), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[11] ), .QN(
        \UUT/Mpath/the_alu/N61 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[9]  ( .D(n3466), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[9] ), .QN(
        \UUT/Mpath/the_alu/N65 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[12]  ( .D(n3348), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[12] ), .QN(
        \UUT/Mpath/the_alu/N59 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[8]  ( .D(n3506), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[8] ), .QN(
        \UUT/Mpath/the_alu/N67 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[19]  ( .D(n3068), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[19] ), .QN(
        \UUT/Mpath/the_alu/N45 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[18]  ( .D(n3108), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[18] ), .QN(
        \UUT/Mpath/the_alu/N47 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[14]  ( .D(n3263), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[14] ), .QN(
        \UUT/Mpath/the_alu/N56 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[20]  ( .D(n3028), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[20] ), .QN(
        \UUT/Mpath/the_alu/N43 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[10]  ( .D(n3422), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[10] ), .QN(
        \UUT/Mpath/the_alu/N64 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[18]  ( .D(n3103), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[18] ), .QN(
        \UUT/Mpath/the_alu/N48 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[12]  ( .D(n3343), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[12] ), .QN(
        \UUT/Mpath/the_alu/N60 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[16]  ( .D(n3188), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[16] ), .QN(
        \UUT/Mpath/the_alu/N51 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[13]  ( .D(n3308), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[13] ), .QN(
        \UUT/Mpath/the_alu/N57 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[13]  ( .D(n3303), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[13] ), .QN(
        \UUT/Mpath/the_alu/N58 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[10]  ( .D(n3427), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[10] ), .QN(
        \UUT/Mpath/the_alu/N63 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[5]  ( .D(n3621), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[5] ), .QN(
        \UUT/Mpath/the_alu/N74 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[14]  ( .D(n3268), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[14] ), .QN(
        \UUT/Mpath/the_alu/N55 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[15]  ( .D(n3228), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[15] ), .QN(
        \UUT/Mpath/the_alu/N53 ) );
  DFFR_X1 \UUT/Mpath/regA/data_out_reg[6]  ( .D(n3586), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regA[6] ), .QN(
        \UUT/Mpath/the_alu/N71 ) );
  DFFR_X1 \UUT/Mpath/regB/data_out_reg[6]  ( .D(n3581), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[6] ), .QN(
        \UUT/Mpath/the_alu/N72 ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[15]  ( .D(n3221), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [15]), 
        .QN(n6841) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[5]  ( .D(n3620), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7079) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[3]  ( .D(n3700), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7065) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[11]  ( .D(n3382), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7057) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[21]  ( .D(n2981), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7052) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[23]  ( .D(n2868), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7047) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[27]  ( .D(n4240), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [27]), .QN(n2764)
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[9]  ( .D(n3460), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7031) );
  DFFR_X2 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[57]  ( .D(n4305), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[57] ) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[13]  ( .D(n3301), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n7005) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[27]  ( .D(n2884), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6972) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[7]  ( .D(n3540), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6964) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[25]  ( .D(n2896), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6962) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[28]  ( .D(n4241), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [28]), .QN(n2765)
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[19]  ( .D(n3061), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6937) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[22]  ( .D(n2941), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [22])
         );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[17]  ( .D(n3141), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6914) );
  DFFR_X2 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[3]  ( .D(n3702), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/acc_out[35] ), 
        .QN(n5597) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[23]  ( .D(n4159), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [23]), .QN(
        n2710) );
  DFFS_X2 \UUT/Mcontrol/Program_counter/out_pc_reg[6]  ( .D(n3579), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [6]), .QN(
        n2687) );
  DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[15]  ( .D(n3222), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/f_currpc [15]), .QN(
        n2663) );
  DFFR_X2 \UUT/Mpath/the_mult/multb/data_out_reg[30]  ( .D(n2870), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [30])
         );
  DFFR_X2 \UUT/Mpath/regB/data_out_reg[30]  ( .D(n2871), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/out_regB[30] ), .QN(
        \UUT/Mpath/the_alu/N24 ) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[SIGN]  ( .D(n4236), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), .QN(n1099) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MR]  ( .D(n4234), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(n1095) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MH]  ( .D(n4233), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(n1090) );
  DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MB]  ( .D(n4232), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .QN(n1083) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[0]  ( .D(n4158), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n995), .QN(n5524) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[1]  ( .D(n4156), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n896), .QN(n5957) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[2]  ( .D(n4155), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n830), .QN(n6211) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[3]  ( .D(n4154), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n801), .QN(n6200) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[4]  ( .D(n4153), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n776), .QN(n6188) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[5]  ( .D(n4152), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n751), .QN(n6179) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[0]  ( .D(n3783), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n839), .QN(n5590) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[6]  ( .D(n4151), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n726), .QN(n6170) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[31]  ( .D(n4076), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n108), .QN(n5542) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[29]  ( .D(n2876), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n120), .QN(n5548) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[26]  ( .D(n2894), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n172), .QN(n5554) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[23]  ( .D(n3855), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n862), .QN(n5560) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[20]  ( .D(n3026), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n356), .QN(n5566) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[17]  ( .D(n3146), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n431), .QN(n5574) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[14]  ( .D(n3266), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n515), .QN(n5580) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[11]  ( .D(n3386), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n588), .QN(n5586) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[8]  ( .D(n3504), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n658), .QN(n5530) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[5]  ( .D(n3624), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n737), .QN(n5536) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[2]  ( .D(n3744), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n812), .QN(n5546) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[7]  ( .D(n4150), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n696), .QN(n6161) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[6]  ( .D(n3584), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n707), .QN(n5534) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[30]  ( .D(n4126), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n923), .QN(n5544) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[28]  ( .D(n2882), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n138), .QN(n5550) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[27]  ( .D(n2888), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n155), .QN(n5552) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[25]  ( .D(n2900), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n188), .QN(n5556) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[24]  ( .D(n2906), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n211), .QN(n5558) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[22]  ( .D(n2946), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n308), .QN(n5562) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[21]  ( .D(n2986), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n333), .QN(n5564) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[19]  ( .D(n3066), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n383), .QN(n5570) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[18]  ( .D(n3106), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n407), .QN(n5572) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[16]  ( .D(n3186), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n460), .QN(n5576) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[15]  ( .D(n3226), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n488), .QN(n5578) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[13]  ( .D(n3306), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n539), .QN(n5582) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[12]  ( .D(n3346), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n564), .QN(n5584) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[10]  ( .D(n3425), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n611), .QN(n5588) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[9]  ( .D(n3464), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n634), .QN(n5528) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[7]  ( .D(n3544), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n682), .QN(n5532) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[4]  ( .D(n3664), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n762), .QN(n5538) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[3]  ( .D(n3704), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n787), .QN(n5540) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[1]  ( .D(n3819), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(n850), .QN(n5568) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[8]  ( .D(n4149), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n671), .QN(n6152) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[9]  ( .D(n4148), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n647), .QN(n6143) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[10]  ( .D(n4147), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n624), .QN(n6241) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[11]  ( .D(n4146), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n601), .QN(n6232) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[12]  ( .D(n4145), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n577), .QN(n6223) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[13]  ( .D(n4144), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n552), .QN(n6093) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[14]  ( .D(n4143), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n528), .QN(n6083) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[15]  ( .D(n4142), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n504), .QN(n6069) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[16]  ( .D(n4141), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n472), .QN(n6058) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[17]  ( .D(n4140), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n443), .QN(n6046) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[18]  ( .D(n4139), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n419), .QN(n6025) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[19]  ( .D(n4138), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n395), .QN(n6012) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[20]  ( .D(n4137), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n368), .QN(n5999) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[21]  ( .D(n4136), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n345), .QN(n5989) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[22]  ( .D(n4135), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n321), .QN(n5979) );
  DFFR_X1 \UUT/Mpath/JAR/data_out_reg[23]  ( .D(n4134), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n954), .QN(n5968) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[31]  ( .D(n4103), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4522) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[30]  ( .D(n4068), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4523) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[29]  ( .D(n4037), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4525) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[28]  ( .D(n4006), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4526) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[27]  ( .D(n3975), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4527) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[26]  ( .D(n3944), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4528) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[25]  ( .D(n3913), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4529) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[24]  ( .D(n2933), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4530) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[23]  ( .D(n3882), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4531) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[22]  ( .D(n2973), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4532) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[21]  ( .D(n3013), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4533) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[20]  ( .D(n3053), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4534) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[19]  ( .D(n3093), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4536) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[18]  ( .D(n3133), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4537) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[17]  ( .D(n3173), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4538) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[16]  ( .D(n3213), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4539) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[15]  ( .D(n3253), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4540) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[14]  ( .D(n3293), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4541) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[13]  ( .D(n3333), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4542) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[12]  ( .D(n3373), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4543) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[11]  ( .D(n3413), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4544) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[10]  ( .D(n3452), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4545) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[9]  ( .D(n3491), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4515) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[8]  ( .D(n3531), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4516) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[7]  ( .D(n3571), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4517) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[6]  ( .D(n3611), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4518) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[5]  ( .D(n3651), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4519) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[4]  ( .D(n3691), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4520) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[3]  ( .D(n3731), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4521) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[2]  ( .D(n3771), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4524) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[1]  ( .D(n3846), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4535) );
  DFFR_X1 \UUT/regfile/rx_3/data_out_reg[0]  ( .D(n3810), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4546) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[31]  ( .D(n4100), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4618) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[30]  ( .D(n4065), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4619) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[29]  ( .D(n4034), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4621) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[28]  ( .D(n4003), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4622) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[27]  ( .D(n3972), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4623) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[26]  ( .D(n3941), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4624) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[25]  ( .D(n3910), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4625) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[24]  ( .D(n2930), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4626) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[23]  ( .D(n3879), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4627) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[22]  ( .D(n2970), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4628) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[21]  ( .D(n3010), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4629) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[20]  ( .D(n3050), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4630) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[19]  ( .D(n3090), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4632) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[18]  ( .D(n3130), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4633) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[17]  ( .D(n3170), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4634) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[16]  ( .D(n3210), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4635) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[15]  ( .D(n3250), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4636) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[14]  ( .D(n3290), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4637) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[13]  ( .D(n3330), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4638) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[12]  ( .D(n3370), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4639) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[11]  ( .D(n3410), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4640) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[10]  ( .D(n3449), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4641) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[9]  ( .D(n3488), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4611) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[8]  ( .D(n3528), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4612) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[7]  ( .D(n3568), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4613) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[6]  ( .D(n3608), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4614) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[5]  ( .D(n3648), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4615) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[4]  ( .D(n3688), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4616) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[3]  ( .D(n3728), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4617) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[2]  ( .D(n3768), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4620) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[1]  ( .D(n3843), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4631) );
  DFFR_X1 \UUT/regfile/rx_2/data_out_reg[0]  ( .D(n3807), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4642) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[31]  ( .D(n4089), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1947), .QN(n4970) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[30]  ( .D(n4054), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1927), .QN(n4971) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[29]  ( .D(n4023), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1887), .QN(n4973) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[28]  ( .D(n3992), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1867), .QN(n4974) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[27]  ( .D(n3961), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1847), .QN(n4975) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[26]  ( .D(n3930), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1827), .QN(n4976) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[25]  ( .D(n3899), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1807), .QN(n4977) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[24]  ( .D(n2919), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1787), .QN(n4978) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[23]  ( .D(n3868), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1767), .QN(n4979) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[22]  ( .D(n2959), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1747), .QN(n4980) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[21]  ( .D(n2999), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1727), .QN(n4981) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[20]  ( .D(n3039), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1707), .QN(n4982) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[19]  ( .D(n3079), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1667), .QN(n4984) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[18]  ( .D(n3119), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1647), .QN(n4985) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[17]  ( .D(n3159), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1627), .QN(n4986) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[16]  ( .D(n3199), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1607), .QN(n4987) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[15]  ( .D(n3239), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1587), .QN(n4988) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[14]  ( .D(n3279), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1567), .QN(n4989) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[13]  ( .D(n3319), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1547), .QN(n4990) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[12]  ( .D(n3359), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1527), .QN(n4991) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[11]  ( .D(n3399), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1507), .QN(n4992) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[10]  ( .D(n3438), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1487), .QN(n4993) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[9]  ( .D(n3477), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2087), .QN(n4963) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[8]  ( .D(n3517), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2067), .QN(n4964) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[7]  ( .D(n3557), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2047), .QN(n4965) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[6]  ( .D(n3597), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2027), .QN(n4966) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[5]  ( .D(n3637), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2007), .QN(n4967) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[4]  ( .D(n3677), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1987), .QN(n4968) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[3]  ( .D(n3717), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1967), .QN(n4969) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[2]  ( .D(n3757), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1907), .QN(n4972) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[1]  ( .D(n3832), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1687), .QN(n4983) );
  DFFR_X1 \UUT/regfile/rx_1/data_out_reg[0]  ( .D(n3796), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1461), .QN(n4994) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[20]  ( .D(n3060), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5393) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[19]  ( .D(n3100), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5399) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[18]  ( .D(n3140), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5402) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[17]  ( .D(n3180), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5405) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[16]  ( .D(n3220), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5408) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[15]  ( .D(n3260), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5411) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[14]  ( .D(n3300), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5414) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[13]  ( .D(n3340), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5417) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[12]  ( .D(n3380), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5420) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[11]  ( .D(n3420), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5423) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[10]  ( .D(n3459), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5426) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[9]  ( .D(n3498), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5335) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[8]  ( .D(n3538), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5339) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[7]  ( .D(n3578), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5342) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[6]  ( .D(n3618), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5345) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[5]  ( .D(n3658), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5348) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[4]  ( .D(n3698), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5351) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[3]  ( .D(n3738), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5354) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[2]  ( .D(n3778), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5363) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[1]  ( .D(n4112), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5396) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[0]  ( .D(n4163), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5429) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[21]  ( .D(n3020), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5390) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[26]  ( .D(n4116), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5375) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[27]  ( .D(n4118), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5372) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[23]  ( .D(n4133), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5384) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[22]  ( .D(n2980), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5387) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[28]  ( .D(n4120), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5369) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[24]  ( .D(n2940), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5381) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[29]  ( .D(n4122), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5366) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[9]  ( .D(n2845), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6288) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[8]  ( .D(n2844), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .QN(n6290) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[15]  ( .D(n2851), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6292) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[14]  ( .D(n2850), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6296) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[13]  ( .D(n2849), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6299) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[12]  ( .D(n2848), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6302) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[11]  ( .D(n2847), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6305) );
  DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[10]  ( .D(n2846), .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .QN(n6308) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[25]  ( .D(n4114), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5378) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[31]  ( .D(n4131), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5357) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[31]  ( .D(n4107), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1952), .QN(n4394) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[30]  ( .D(n4072), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1932), .QN(n4395) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[29]  ( .D(n4041), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1892), .QN(n4397) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[28]  ( .D(n4010), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1872), .QN(n4398) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[27]  ( .D(n3979), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1852), .QN(n4399) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[26]  ( .D(n3948), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1832), .QN(n4400) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[25]  ( .D(n3917), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1812), .QN(n4401) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[24]  ( .D(n2937), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1792), .QN(n4402) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[23]  ( .D(n3886), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1772), .QN(n4403) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[22]  ( .D(n2977), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1752), .QN(n4404) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[21]  ( .D(n3017), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1732), .QN(n4405) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[20]  ( .D(n3057), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1712), .QN(n4406) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[19]  ( .D(n3097), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1672), .QN(n4408) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[18]  ( .D(n3137), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1652), .QN(n4409) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[17]  ( .D(n3177), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1632), .QN(n4410) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[16]  ( .D(n3217), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1612), .QN(n4411) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[15]  ( .D(n3257), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1592), .QN(n4412) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[14]  ( .D(n3297), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1572), .QN(n4413) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[13]  ( .D(n3337), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1552), .QN(n4414) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[12]  ( .D(n3377), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1532), .QN(n4415) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[11]  ( .D(n3417), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1512), .QN(n4416) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[10]  ( .D(n3456), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1492), .QN(n4417) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[9]  ( .D(n3495), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2093), .QN(n4387) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[8]  ( .D(n3535), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2072), .QN(n4388) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[7]  ( .D(n3575), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2052), .QN(n4389) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[6]  ( .D(n3615), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2032), .QN(n4390) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[5]  ( .D(n3655), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2012), .QN(n4391) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[4]  ( .D(n3695), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1992), .QN(n4392) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[3]  ( .D(n3735), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1972), .QN(n4393) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[2]  ( .D(n3775), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1912), .QN(n4396) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[1]  ( .D(n3850), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1692), .QN(n4407) );
  DFFR_X1 \UUT/regfile/rx_7/data_out_reg[0]  ( .D(n3814), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1471), .QN(n4418) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[31]  ( .D(n4106), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1950), .QN(n4426) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[30]  ( .D(n4071), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1930), .QN(n4427) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[29]  ( .D(n4040), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1890), .QN(n4429) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[28]  ( .D(n4009), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1870), .QN(n4430) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[27]  ( .D(n3978), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1850), .QN(n4431) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[26]  ( .D(n3947), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1830), .QN(n4432) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[25]  ( .D(n3916), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1810), .QN(n4433) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[24]  ( .D(n2936), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1790), .QN(n4434) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[23]  ( .D(n3885), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1770), .QN(n4435) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[22]  ( .D(n2976), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1750), .QN(n4436) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[21]  ( .D(n3016), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1730), .QN(n4437) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[20]  ( .D(n3056), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1710), .QN(n4438) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[19]  ( .D(n3096), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1670), .QN(n4440) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[18]  ( .D(n3136), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1650), .QN(n4441) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[17]  ( .D(n3176), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1630), .QN(n4442) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[16]  ( .D(n3216), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1610), .QN(n4443) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[15]  ( .D(n3256), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1590), .QN(n4444) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[14]  ( .D(n3296), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1570), .QN(n4445) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[13]  ( .D(n3336), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1550), .QN(n4446) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[12]  ( .D(n3376), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1530), .QN(n4447) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[11]  ( .D(n3416), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1510), .QN(n4448) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[10]  ( .D(n3455), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1490), .QN(n4449) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[9]  ( .D(n3494), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2091), .QN(n4419) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[8]  ( .D(n3534), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2070), .QN(n4420) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[7]  ( .D(n3574), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2050), .QN(n4421) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[6]  ( .D(n3614), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2030), .QN(n4422) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[5]  ( .D(n3654), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2010), .QN(n4423) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[4]  ( .D(n3694), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1990), .QN(n4424) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[3]  ( .D(n3734), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1970), .QN(n4425) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[2]  ( .D(n3774), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1910), .QN(n4428) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[1]  ( .D(n3849), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1690), .QN(n4439) );
  DFFR_X1 \UUT/regfile/rx_6/data_out_reg[0]  ( .D(n3813), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1467), .QN(n4450) );
  DFFR_X1 \UUT/Mpath/regM/data_out_reg[30]  ( .D(n4129), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5360) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[31]  ( .D(n4080), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5258) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[30]  ( .D(n4045), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5259) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[29]  ( .D(n4014), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5261) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[28]  ( .D(n3983), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5262) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[27]  ( .D(n3952), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5263) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[26]  ( .D(n3921), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5264) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[25]  ( .D(n3890), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5265) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[24]  ( .D(n2910), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5266) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[23]  ( .D(n3859), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5267) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[22]  ( .D(n2950), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5268) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[21]  ( .D(n2990), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5269) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[20]  ( .D(n3030), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5270) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[19]  ( .D(n3070), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5272) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[18]  ( .D(n3110), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5273) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[17]  ( .D(n3150), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5274) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[16]  ( .D(n3190), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5275) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[15]  ( .D(n3230), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5276) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[14]  ( .D(n3270), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5277) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[13]  ( .D(n3310), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5278) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[12]  ( .D(n3350), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5279) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[11]  ( .D(n3390), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5280) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[10]  ( .D(n3429), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5281) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[9]  ( .D(n3468), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5251) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[8]  ( .D(n3508), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5252) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[7]  ( .D(n3548), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5253) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[6]  ( .D(n3588), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5254) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[5]  ( .D(n3628), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5255) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[4]  ( .D(n3668), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5256) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[3]  ( .D(n3708), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5257) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[2]  ( .D(n3748), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5260) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[1]  ( .D(n3823), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5271) );
  DFFR_X1 \UUT/regfile/rx_11/data_out_reg[0]  ( .D(n3787), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5282) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[31]  ( .D(n4079), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5290) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[30]  ( .D(n4044), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5291) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[29]  ( .D(n4013), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5293) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[28]  ( .D(n3982), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5294) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[27]  ( .D(n3951), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5295) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[26]  ( .D(n3920), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5296) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[25]  ( .D(n3889), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5297) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[24]  ( .D(n2909), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5298) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[23]  ( .D(n3858), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5299) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[22]  ( .D(n2949), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5300) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[21]  ( .D(n2989), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5301) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[20]  ( .D(n3029), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5302) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[19]  ( .D(n3069), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5304) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[18]  ( .D(n3109), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5305) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[17]  ( .D(n3149), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5306) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[16]  ( .D(n3189), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5307) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[15]  ( .D(n3229), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5308) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[14]  ( .D(n3269), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5309) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[13]  ( .D(n3309), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5310) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[12]  ( .D(n3349), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5311) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[11]  ( .D(n3389), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5312) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[10]  ( .D(n3428), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5313) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[9]  ( .D(n3467), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5283) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[8]  ( .D(n3507), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5284) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[7]  ( .D(n3547), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5285) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[6]  ( .D(n3587), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5286) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[5]  ( .D(n3627), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5287) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[4]  ( .D(n3667), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5288) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[3]  ( .D(n3707), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5289) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[2]  ( .D(n3747), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5292) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[1]  ( .D(n3822), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5303) );
  DFFR_X1 \UUT/regfile/rx_10/data_out_reg[0]  ( .D(n3786), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5314) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[31]  ( .D(n4109), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1951), .QN(n4330) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[30]  ( .D(n4074), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1931), .QN(n4331) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[29]  ( .D(n4043), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1891), .QN(n4333) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[28]  ( .D(n4012), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1871), .QN(n4334) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[27]  ( .D(n3981), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1851), .QN(n4335) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[26]  ( .D(n3950), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1831), .QN(n4336) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[25]  ( .D(n3919), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1811), .QN(n4337) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[24]  ( .D(n2939), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1791), .QN(n4338) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[23]  ( .D(n3888), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1771), .QN(n4339) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[22]  ( .D(n2979), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1751), .QN(n4340) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[21]  ( .D(n3019), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1731), .QN(n4341) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[20]  ( .D(n3059), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1711), .QN(n4342) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[19]  ( .D(n3099), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1671), .QN(n4344) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[18]  ( .D(n3139), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1651), .QN(n4345) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[17]  ( .D(n3179), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1631), .QN(n4346) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[16]  ( .D(n3219), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1611), .QN(n4347) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[15]  ( .D(n3259), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1591), .QN(n4348) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[14]  ( .D(n3299), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1571), .QN(n4349) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[13]  ( .D(n3339), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1551), .QN(n4350) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[12]  ( .D(n3379), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1531), .QN(n4351) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[11]  ( .D(n3419), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1511), .QN(n4352) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[10]  ( .D(n3458), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1491), .QN(n4353) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[9]  ( .D(n3497), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2092), .QN(n4323) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[8]  ( .D(n3537), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2071), .QN(n4324) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[7]  ( .D(n3577), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2051), .QN(n4325) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[6]  ( .D(n3617), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2031), .QN(n4326) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[5]  ( .D(n3657), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2011), .QN(n4327) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[4]  ( .D(n3697), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1991), .QN(n4328) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[3]  ( .D(n3737), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1971), .QN(n4329) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[2]  ( .D(n3777), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1911), .QN(n4332) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[1]  ( .D(n3852), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1691), .QN(n4343) );
  DFFR_X1 \UUT/regfile/rx_9/data_out_reg[0]  ( .D(n3816), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1470), .QN(n4354) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[31]  ( .D(n4108), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4362) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[30]  ( .D(n4073), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4363) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[29]  ( .D(n4042), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4365) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[28]  ( .D(n4011), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4366) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[27]  ( .D(n3980), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4367) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[26]  ( .D(n3949), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4368) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[25]  ( .D(n3918), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4369) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[24]  ( .D(n2938), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4370) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[23]  ( .D(n3887), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4371) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[22]  ( .D(n2978), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4372) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[21]  ( .D(n3018), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4373) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[20]  ( .D(n3058), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4374) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[19]  ( .D(n3098), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4376) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[18]  ( .D(n3138), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4377) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[17]  ( .D(n3178), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4378) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[16]  ( .D(n3218), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4379) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[15]  ( .D(n3258), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4380) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[14]  ( .D(n3298), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4381) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[13]  ( .D(n3338), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4382) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[12]  ( .D(n3378), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4383) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[11]  ( .D(n3418), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4384) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[10]  ( .D(n3457), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4385) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[9]  ( .D(n3496), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4355) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[8]  ( .D(n3536), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4356) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[7]  ( .D(n3576), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4357) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[6]  ( .D(n3616), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4358) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[5]  ( .D(n3656), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4359) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[4]  ( .D(n3696), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4360) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[3]  ( .D(n3736), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4361) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[2]  ( .D(n3776), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4364) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[1]  ( .D(n3851), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4375) );
  DFFR_X1 \UUT/regfile/rx_8/data_out_reg[0]  ( .D(n3815), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4386) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[31]  ( .D(n4084), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5130) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[30]  ( .D(n4049), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5131) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[29]  ( .D(n4018), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5133) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[28]  ( .D(n3987), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5134) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[27]  ( .D(n3956), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5135) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[26]  ( .D(n3925), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5136) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[25]  ( .D(n3894), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5137) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[24]  ( .D(n2914), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5138) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[23]  ( .D(n3863), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5139) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[22]  ( .D(n2954), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5140) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[21]  ( .D(n2994), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5141) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[20]  ( .D(n3034), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5142) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[19]  ( .D(n3074), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5144) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[18]  ( .D(n3114), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5145) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[17]  ( .D(n3154), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5146) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[16]  ( .D(n3194), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5147) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[15]  ( .D(n3234), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5148) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[14]  ( .D(n3274), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5149) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[13]  ( .D(n3314), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5150) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[12]  ( .D(n3354), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5151) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[11]  ( .D(n3394), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5152) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[10]  ( .D(n3433), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5153) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[9]  ( .D(n3472), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5123) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[8]  ( .D(n3512), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5124) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[7]  ( .D(n3552), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5125) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[6]  ( .D(n3592), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5126) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[5]  ( .D(n3632), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5127) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[4]  ( .D(n3672), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5128) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[3]  ( .D(n3712), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5129) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[2]  ( .D(n3752), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5132) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[1]  ( .D(n3827), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5143) );
  DFFR_X1 \UUT/regfile/rx_15/data_out_reg[0]  ( .D(n3791), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5154) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[31]  ( .D(n4083), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5162) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[30]  ( .D(n4048), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5163) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[29]  ( .D(n4017), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5165) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[28]  ( .D(n3986), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5166) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[27]  ( .D(n3955), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5167) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[26]  ( .D(n3924), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5168) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[25]  ( .D(n3893), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5169) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[24]  ( .D(n2913), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5170) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[23]  ( .D(n3862), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5171) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[22]  ( .D(n2953), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5172) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[21]  ( .D(n2993), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5173) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[20]  ( .D(n3033), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5174) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[19]  ( .D(n3073), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5176) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[18]  ( .D(n3113), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5177) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[17]  ( .D(n3153), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5178) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[16]  ( .D(n3193), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5179) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[15]  ( .D(n3233), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5180) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[14]  ( .D(n3273), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5181) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[13]  ( .D(n3313), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5182) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[12]  ( .D(n3353), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5183) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[11]  ( .D(n3393), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5184) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[10]  ( .D(n3432), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5185) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[9]  ( .D(n3471), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5155) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[8]  ( .D(n3511), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5156) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[7]  ( .D(n3551), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5157) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[6]  ( .D(n3591), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5158) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[5]  ( .D(n3631), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5159) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[4]  ( .D(n3671), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5160) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[3]  ( .D(n3711), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5161) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[2]  ( .D(n3751), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5164) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[1]  ( .D(n3826), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5175) );
  DFFR_X1 \UUT/regfile/rx_14/data_out_reg[0]  ( .D(n3790), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5186) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[31]  ( .D(n4082), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2219), .QN(n5194) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[30]  ( .D(n4047), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2206), .QN(n5195) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[29]  ( .D(n4016), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2193), .QN(n5197) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[28]  ( .D(n3985), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2180), .QN(n5198) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[27]  ( .D(n3954), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2167), .QN(n5199) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[26]  ( .D(n3923), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2154), .QN(n5200) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[25]  ( .D(n3892), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2141), .QN(n5201) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[24]  ( .D(n2912), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2128), .QN(n5202) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[23]  ( .D(n3861), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2277), .QN(n5203) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[22]  ( .D(n2952), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2290), .QN(n5204) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[21]  ( .D(n2992), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2303), .QN(n5205) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[20]  ( .D(n3032), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2316), .QN(n5206) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[19]  ( .D(n3072), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2342), .QN(n5208) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[18]  ( .D(n3112), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2355), .QN(n5209) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[17]  ( .D(n3152), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2368), .QN(n5210) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[16]  ( .D(n3192), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2381), .QN(n5211) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[15]  ( .D(n3232), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2394), .QN(n5212) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[14]  ( .D(n3272), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2407), .QN(n5213) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[13]  ( .D(n3312), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2420), .QN(n5214) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[12]  ( .D(n3352), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2454), .QN(n5215) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[11]  ( .D(n3392), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2470), .QN(n5216) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[10]  ( .D(n3431), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2486), .QN(n5217) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[9]  ( .D(n3470), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2502), .QN(n5187) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[8]  ( .D(n3510), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2518), .QN(n5188) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[7]  ( .D(n3550), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2534), .QN(n5189) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[6]  ( .D(n3590), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2550), .QN(n5190) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[5]  ( .D(n3630), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2568), .QN(n5191) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[4]  ( .D(n3670), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2583), .QN(n5192) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[3]  ( .D(n3710), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2604), .QN(n5193) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[2]  ( .D(n3750), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2438), .QN(n5196) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[1]  ( .D(n3825), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2329), .QN(n5207) );
  DFFR_X1 \UUT/regfile/rx_13/data_out_reg[0]  ( .D(n3789), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2110), .QN(n5218) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[31]  ( .D(n4081), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1948), .QN(n5226) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[30]  ( .D(n4046), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1928), .QN(n5227) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[29]  ( .D(n4015), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1888), .QN(n5229) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[28]  ( .D(n3984), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1868), .QN(n5230) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[27]  ( .D(n3953), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1848), .QN(n5231) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[26]  ( .D(n3922), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1828), .QN(n5232) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[25]  ( .D(n3891), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1808), .QN(n5233) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[24]  ( .D(n2911), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1788), .QN(n5234) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[23]  ( .D(n3860), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1768), .QN(n5235) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[22]  ( .D(n2951), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1748), .QN(n5236) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[21]  ( .D(n2991), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1728), .QN(n5237) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[20]  ( .D(n3031), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1708), .QN(n5238) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[19]  ( .D(n3071), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1668), .QN(n5240) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[18]  ( .D(n3111), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1648), .QN(n5241) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[17]  ( .D(n3151), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1628), .QN(n5242) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[16]  ( .D(n3191), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1608), .QN(n5243) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[15]  ( .D(n3231), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1588), .QN(n5244) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[14]  ( .D(n3271), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1568), .QN(n5245) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[13]  ( .D(n3311), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1548), .QN(n5246) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[12]  ( .D(n3351), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1528), .QN(n5247) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[11]  ( .D(n3391), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1508), .QN(n5248) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[10]  ( .D(n3430), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1488), .QN(n5249) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[9]  ( .D(n3469), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2088), .QN(n5219) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[8]  ( .D(n3509), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2068), .QN(n5220) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[7]  ( .D(n3549), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2048), .QN(n5221) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[6]  ( .D(n3589), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2028), .QN(n5222) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[5]  ( .D(n3629), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2008), .QN(n5223) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[4]  ( .D(n3669), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1988), .QN(n5224) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[3]  ( .D(n3709), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1968), .QN(n5225) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[2]  ( .D(n3749), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1908), .QN(n5228) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[1]  ( .D(n3824), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1688), .QN(n5239) );
  DFFR_X1 \UUT/regfile/rx_12/data_out_reg[0]  ( .D(n3788), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1463), .QN(n5250) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[31]  ( .D(n4086), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5066) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[30]  ( .D(n4051), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5067) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[29]  ( .D(n4020), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5069) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[28]  ( .D(n3989), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5070) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[27]  ( .D(n3958), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5071) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[26]  ( .D(n3927), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5072) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[25]  ( .D(n3896), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5073) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[24]  ( .D(n2916), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5074) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[23]  ( .D(n3865), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5075) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[22]  ( .D(n2956), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5076) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[21]  ( .D(n2996), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5077) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[20]  ( .D(n3036), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5078) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[19]  ( .D(n3076), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5080) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[18]  ( .D(n3116), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5081) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[17]  ( .D(n3156), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5082) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[16]  ( .D(n3196), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5083) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[15]  ( .D(n3236), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5084) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[14]  ( .D(n3276), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5085) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[13]  ( .D(n3316), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5086) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[12]  ( .D(n3356), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5087) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[11]  ( .D(n3396), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5088) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[10]  ( .D(n3435), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5089) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[9]  ( .D(n3474), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5059) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[8]  ( .D(n3514), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5060) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[7]  ( .D(n3554), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5061) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[6]  ( .D(n3594), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5062) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[5]  ( .D(n3634), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5063) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[4]  ( .D(n3674), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5064) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[3]  ( .D(n3714), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5065) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[2]  ( .D(n3754), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5068) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[1]  ( .D(n3829), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5079) );
  DFFR_X1 \UUT/regfile/rx_17/data_out_reg[0]  ( .D(n3793), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5090) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[31]  ( .D(n4085), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5098) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[30]  ( .D(n4050), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5099) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[29]  ( .D(n4019), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5101) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[28]  ( .D(n3988), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5102) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[27]  ( .D(n3957), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5103) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[26]  ( .D(n3926), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5104) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[25]  ( .D(n3895), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5105) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[24]  ( .D(n2915), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5106) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[23]  ( .D(n3864), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5107) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[22]  ( .D(n2955), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5108) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[21]  ( .D(n2995), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5109) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[20]  ( .D(n3035), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5110) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[19]  ( .D(n3075), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5112) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[18]  ( .D(n3115), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5113) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[17]  ( .D(n3155), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5114) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[16]  ( .D(n3195), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5115) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[15]  ( .D(n3235), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5116) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[14]  ( .D(n3275), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5117) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[13]  ( .D(n3315), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5118) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[12]  ( .D(n3355), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5119) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[11]  ( .D(n3395), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5120) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[10]  ( .D(n3434), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5121) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[9]  ( .D(n3473), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5091) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[8]  ( .D(n3513), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5092) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[7]  ( .D(n3553), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5093) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[6]  ( .D(n3593), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5094) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[5]  ( .D(n3633), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5095) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[4]  ( .D(n3673), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5096) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[3]  ( .D(n3713), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5097) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[2]  ( .D(n3753), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5100) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[1]  ( .D(n3828), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5111) );
  DFFR_X1 \UUT/regfile/rx_16/data_out_reg[0]  ( .D(n3792), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5122) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[31]  ( .D(n4097), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4714) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[30]  ( .D(n4062), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4715) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[29]  ( .D(n4031), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4717) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[28]  ( .D(n4000), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4718) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[27]  ( .D(n3969), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4719) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[26]  ( .D(n3938), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4720) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[25]  ( .D(n3907), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4721) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[24]  ( .D(n2927), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4722) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[23]  ( .D(n3876), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4723) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[22]  ( .D(n2967), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4724) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[21]  ( .D(n3007), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4725) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[20]  ( .D(n3047), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4726) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[19]  ( .D(n3087), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4728) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[18]  ( .D(n3127), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4729) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[17]  ( .D(n3167), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4730) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[16]  ( .D(n3207), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4731) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[15]  ( .D(n3247), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4732) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[14]  ( .D(n3287), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4733) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[13]  ( .D(n3327), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4734) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[12]  ( .D(n3367), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4735) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[11]  ( .D(n3407), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4736) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[10]  ( .D(n3446), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4737) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[9]  ( .D(n3485), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4707) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[8]  ( .D(n3525), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4708) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[7]  ( .D(n3565), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4709) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[6]  ( .D(n3605), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4710) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[5]  ( .D(n3645), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4711) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[4]  ( .D(n3685), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4712) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[3]  ( .D(n3725), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4713) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[2]  ( .D(n3765), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4716) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[1]  ( .D(n3840), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4727) );
  DFFR_X1 \UUT/regfile/rx_27/data_out_reg[0]  ( .D(n3804), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4738) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[31]  ( .D(n4096), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1944), .QN(n4746) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[30]  ( .D(n4061), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1924), .QN(n4747) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[29]  ( .D(n4030), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1884), .QN(n4749) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[28]  ( .D(n3999), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1864), .QN(n4750) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[27]  ( .D(n3968), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1844), .QN(n4751) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[26]  ( .D(n3937), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1824), .QN(n4752) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[25]  ( .D(n3906), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1804), .QN(n4753) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[24]  ( .D(n2926), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1784), .QN(n4754) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[23]  ( .D(n3875), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1764), .QN(n4755) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[22]  ( .D(n2966), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1744), .QN(n4756) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[21]  ( .D(n3006), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1724), .QN(n4757) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[20]  ( .D(n3046), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1704), .QN(n4758) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[19]  ( .D(n3086), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1664), .QN(n4760) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[18]  ( .D(n3126), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1644), .QN(n4761) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[17]  ( .D(n3166), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1624), .QN(n4762) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[16]  ( .D(n3206), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1604), .QN(n4763) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[15]  ( .D(n3246), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1584), .QN(n4764) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[14]  ( .D(n3286), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1564), .QN(n4765) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[13]  ( .D(n3326), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1544), .QN(n4766) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[12]  ( .D(n3366), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1524), .QN(n4767) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[11]  ( .D(n3406), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1504), .QN(n4768) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[10]  ( .D(n3445), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1484), .QN(n4769) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[9]  ( .D(n3484), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2084), .QN(n4739) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[8]  ( .D(n3524), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2064), .QN(n4740) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[7]  ( .D(n3564), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2044), .QN(n4741) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[6]  ( .D(n3604), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2024), .QN(n4742) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[5]  ( .D(n3644), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2004), .QN(n4743) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[4]  ( .D(n3684), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1984), .QN(n4744) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[3]  ( .D(n3724), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1964), .QN(n4745) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[2]  ( .D(n3764), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1904), .QN(n4748) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[1]  ( .D(n3839), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1684), .QN(n4759) );
  DFFR_X1 \UUT/regfile/rx_26/data_out_reg[0]  ( .D(n3803), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1456), .QN(n4770) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[31]  ( .D(n4093), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1942), .QN(n4842) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[30]  ( .D(n4058), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1922), .QN(n4843) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[29]  ( .D(n4027), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1882), .QN(n4845) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[28]  ( .D(n3996), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1862), .QN(n4846) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[27]  ( .D(n3965), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1842), .QN(n4847) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[26]  ( .D(n3934), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1822), .QN(n4848) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[25]  ( .D(n3903), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1802), .QN(n4849) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[24]  ( .D(n2923), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1782), .QN(n4850) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[23]  ( .D(n3872), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1762), .QN(n4851) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[22]  ( .D(n2963), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1742), .QN(n4852) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[21]  ( .D(n3003), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1722), .QN(n4853) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[20]  ( .D(n3043), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1702), .QN(n4854) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[19]  ( .D(n3083), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1662), .QN(n4856) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[18]  ( .D(n3123), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1642), .QN(n4857) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[17]  ( .D(n3163), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1622), .QN(n4858) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[16]  ( .D(n3203), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1602), .QN(n4859) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[15]  ( .D(n3243), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1582), .QN(n4860) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[14]  ( .D(n3283), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1562), .QN(n4861) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[13]  ( .D(n3323), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1542), .QN(n4862) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[12]  ( .D(n3363), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1522), .QN(n4863) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[11]  ( .D(n3403), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1502), .QN(n4864) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[10]  ( .D(n3442), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1482), .QN(n4865) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[9]  ( .D(n3481), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2082), .QN(n4835) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[8]  ( .D(n3521), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2062), .QN(n4836) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[7]  ( .D(n3561), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2042), .QN(n4837) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[6]  ( .D(n3601), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2022), .QN(n4838) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[5]  ( .D(n3641), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2002), .QN(n4839) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[4]  ( .D(n3681), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1982), .QN(n4840) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[3]  ( .D(n3721), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1962), .QN(n4841) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[2]  ( .D(n3761), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1902), .QN(n4844) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[1]  ( .D(n3836), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1682), .QN(n4855) );
  DFFR_X1 \UUT/regfile/rx_23/data_out_reg[0]  ( .D(n3800), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1452), .QN(n4866) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[31]  ( .D(n4092), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1943), .QN(n4874) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[30]  ( .D(n4057), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1923), .QN(n4875) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[29]  ( .D(n4026), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1883), .QN(n4877) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[28]  ( .D(n3995), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1863), .QN(n4878) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[27]  ( .D(n3964), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1843), .QN(n4879) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[26]  ( .D(n3933), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1823), .QN(n4880) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[25]  ( .D(n3902), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1803), .QN(n4881) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[24]  ( .D(n2922), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1783), .QN(n4882) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[23]  ( .D(n3871), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1763), .QN(n4883) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[22]  ( .D(n2962), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1743), .QN(n4884) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[21]  ( .D(n3002), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1723), .QN(n4885) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[20]  ( .D(n3042), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1703), .QN(n4886) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[19]  ( .D(n3082), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1663), .QN(n4888) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[18]  ( .D(n3122), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1643), .QN(n4889) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[17]  ( .D(n3162), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1623), .QN(n4890) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[16]  ( .D(n3202), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1603), .QN(n4891) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[15]  ( .D(n3242), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1583), .QN(n4892) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[14]  ( .D(n3282), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1563), .QN(n4893) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[13]  ( .D(n3322), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1543), .QN(n4894) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[12]  ( .D(n3362), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1523), .QN(n4895) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[11]  ( .D(n3402), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1503), .QN(n4896) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[10]  ( .D(n3441), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1483), .QN(n4897) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[9]  ( .D(n3480), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2083), .QN(n4867) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[8]  ( .D(n3520), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2063), .QN(n4868) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[7]  ( .D(n3560), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2043), .QN(n4869) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[6]  ( .D(n3600), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2023), .QN(n4870) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[5]  ( .D(n3640), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n2003), .QN(n4871) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[4]  ( .D(n3680), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1983), .QN(n4872) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[3]  ( .D(n3720), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1963), .QN(n4873) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[2]  ( .D(n3760), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1903), .QN(n4876) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[1]  ( .D(n3835), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1683), .QN(n4887) );
  DFFR_X1 \UUT/regfile/rx_22/data_out_reg[0]  ( .D(n3799), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(n1454), .QN(n4898) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[31]  ( .D(n4102), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4554) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[30]  ( .D(n4067), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4555) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[29]  ( .D(n4036), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4557) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[28]  ( .D(n4005), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4558) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[27]  ( .D(n3974), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4559) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[26]  ( .D(n3943), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4560) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[25]  ( .D(n3912), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4561) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[24]  ( .D(n2932), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4562) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[23]  ( .D(n3881), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4563) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[22]  ( .D(n2972), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4564) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[21]  ( .D(n3012), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4565) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[20]  ( .D(n3052), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4566) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[19]  ( .D(n3092), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4568) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[18]  ( .D(n3132), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4569) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[17]  ( .D(n3172), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4570) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[16]  ( .D(n3212), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4571) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[15]  ( .D(n3252), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4572) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[14]  ( .D(n3292), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4573) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[13]  ( .D(n3332), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4574) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[12]  ( .D(n3372), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4575) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[11]  ( .D(n3412), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4576) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[10]  ( .D(n3451), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4577) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[9]  ( .D(n3490), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4547) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[8]  ( .D(n3530), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4548) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[7]  ( .D(n3570), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4549) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[6]  ( .D(n3610), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4550) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[5]  ( .D(n3650), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4551) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[4]  ( .D(n3690), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4552) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[3]  ( .D(n3730), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4553) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[2]  ( .D(n3770), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4556) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[1]  ( .D(n3845), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4567) );
  DFFR_X1 \UUT/regfile/rx_31/data_out_reg[0]  ( .D(n3809), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4578) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[31]  ( .D(n4101), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4586) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[30]  ( .D(n4066), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4587) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[29]  ( .D(n4035), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4589) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[28]  ( .D(n4004), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4590) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[27]  ( .D(n3973), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4591) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[26]  ( .D(n3942), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4592) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[25]  ( .D(n3911), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4593) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[24]  ( .D(n2931), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4594) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[23]  ( .D(n3880), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4595) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[22]  ( .D(n2971), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4596) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[21]  ( .D(n3011), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4597) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[20]  ( .D(n3051), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4598) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[19]  ( .D(n3091), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4600) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[18]  ( .D(n3131), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4601) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[17]  ( .D(n3171), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4602) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[16]  ( .D(n3211), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4603) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[15]  ( .D(n3251), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4604) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[14]  ( .D(n3291), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4605) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[13]  ( .D(n3331), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4606) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[12]  ( .D(n3371), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4607) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[11]  ( .D(n3411), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4608) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[10]  ( .D(n3450), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4609) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[9]  ( .D(n3489), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4579) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[8]  ( .D(n3529), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4580) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[7]  ( .D(n3569), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4581) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[6]  ( .D(n3609), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4582) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[5]  ( .D(n3649), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4583) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[4]  ( .D(n3689), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4584) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[3]  ( .D(n3729), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4585) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[2]  ( .D(n3769), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4588) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[1]  ( .D(n3844), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4599) );
  DFFR_X1 \UUT/regfile/rx_30/data_out_reg[0]  ( .D(n3808), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n4610) );
  DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[0]  ( .D(n4244), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/m_sampled_xrd[0] ), .QN(
        n1112) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[0]  ( .D(n4248), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[0] ), .QN(n840) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[4]  ( .D(n4204), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[4] ), .QN(n1052) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[5]  ( .D(n4209), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[5] ), .QN(n1060) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[2]  ( .D(n4194), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[2] ), .QN(n1040) );
  DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[1]  ( .D(n4188), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/x_mul_command[1] ), .QN(n1032) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[1]  ( .D(n4249), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[1] ), .QN(n851) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[2]  ( .D(n4250), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[2] ), .QN(n813) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[3]  ( .D(n4251), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[3] ), .QN(n788) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[3]  ( .D(n4178), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[3] ), .QN(n1022) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[2]  ( .D(n4176), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[2] ), .QN(n1020) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[1]  ( .D(n4174), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[1] ), .QN(n1014) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[0]  ( .D(n4245), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[0] ), .QN(n1111) );
  DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[4]  ( .D(n4180), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/x_rd[4] ), .QN(n1024) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[4]  ( .D(n4252), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[4] ), .QN(n763) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[5]  ( .D(n4253), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[5] ), .QN(n738) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[6]  ( .D(n4254), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[6] ), .QN(n708) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[7]  ( .D(n4255), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[7] ), .QN(n683) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[8]  ( .D(n4256), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[8] ), .QN(n659) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[9]  ( .D(n4257), .CK(
        CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[9] ), .QN(n635) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[10]  ( .D(n4258), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[10] ), .QN(n612) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[11]  ( .D(n4259), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[11] ), .QN(n589) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[13]  ( .D(n4261), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[13] ), .QN(n540) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[12]  ( .D(n4260), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[12] ), .QN(n565) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[14]  ( .D(n4262), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[14] ), .QN(n516) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[15]  ( .D(n4263), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[15] ), .QN(n489) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[16]  ( .D(n4264), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[16] ), .QN(n461) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[17]  ( .D(n4265), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[17] ), .QN(n432) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[18]  ( .D(n4266), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[18] ), .QN(n408) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[19]  ( .D(n4267), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[19] ), .QN(n384) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[20]  ( .D(n4268), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[20] ), .QN(n357) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[21]  ( .D(n4269), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[21] ), .QN(n334) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[26]  ( .D(n4274), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[26] ), .QN(n173) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[27]  ( .D(n4275), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[27] ), .QN(n156) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[28]  ( .D(n4276), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[28] ), .QN(n139) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[25]  ( .D(n4273), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[25] ), .QN(n189) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[23]  ( .D(n4271), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[23] ), .QN(n863) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[22]  ( .D(n4270), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[22] ), .QN(n309) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[29]  ( .D(n4277), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[29] ), .QN(n116) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[24]  ( .D(n4272), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[24] ), .QN(n212) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[25]  ( .D(n4231), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [25]), 
        .QN(n5753) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[24]  ( .D(n4230), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5760) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[23]  ( .D(n4229), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .QN(n5768) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[22]  ( .D(n4228), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [22]), 
        .QN(n5775) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[21]  ( .D(n4227), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [21]), 
        .QN(n5907) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[20]  ( .D(n4226), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [20]), 
        .QN(n5899) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[19]  ( .D(n4225), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [19]), 
        .QN(n5901) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[18]  ( .D(n4224), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [18]), 
        .QN(n5896) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[17]  ( .D(n4223), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [17]), 
        .QN(n5904) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[16]  ( .D(n4222), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [16]), 
        .QN(n5897) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[15]  ( .D(n4221), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [15]), 
        .QN(n5720) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[14]  ( .D(n4220), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [14]), 
        .QN(n5902) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[13]  ( .D(n4219), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [13]), 
        .QN(n5903) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[12]  ( .D(n4218), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [12]), 
        .QN(n5905) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[11]  ( .D(n4217), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [11]), 
        .QN(n5906) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[10]  ( .D(n4216), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [10]), 
        .QN(n5762) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[9]  ( .D(n4215), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [9]), 
        .QN(n5769) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[8]  ( .D(n4214), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_sampled_finstr [8]), 
        .QN(n5776) );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[7]  ( .D(n4213), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [7]), .QN(n5971)
         );
  DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[6]  ( .D(n4212), .CK(CLK), .RN(
        \UUT/Mcontrol/int_reset ), .Q(\UUT/Mcontrol/d_instr [6]), .QN(n6035)
         );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[32]  ( .D(n4280), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[32] ), .QN(n837) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[30]  ( .D(n4278), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[30] ), .QN(n921) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[31]  ( .D(n4279), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[31] ), .QN(n873) );
  DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[33]  ( .D(n4281), 
        .CK(CLK), .RN(\UUT/Mcontrol/int_reset ), .Q(
        \UUT/Mpath/the_mult/Mult_out[33] ), .QN(n848) );
  DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[20]  ( .D(n3027), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[20] ), 
        .QN(n359) );
  DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[31]  ( .D(n2869), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand2 [31]), 
        .QN(n6358) );
  DFFS_X2 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MR]  ( .D(n4169), .CK(CLK), 
        .SN(\UUT/Mcontrol/int_reset ), .Q(\UUT/m_mem_command[MR] ), .QN(n5623)
         );
  DFFR_X2 \UUT/Mpath/the_mult/multa/data_out_reg[0]  ( .D(n3784), .CK(CLK), 
        .RN(\UUT/Mcontrol/int_reset ), .Q(\UUT/Mpath/the_mult/x_operand1[0] )
         );
  NAND2_X4 U5175 ( .A1(n5893), .A2(n5888), .ZN(n5656) );
  NAND3_X4 U5176 ( .A1(n5883), .A2(n2090), .A3(n5895), .ZN(n1466) );
  AND4_X2 U5177 ( .A1(\UUT/Mcontrol/N22 ), .A2(n932), .A3(n5315), .A4(n933), 
        .ZN(n109) );
  INV_X1 U5178 ( .A(\UUT/branch_rega [4]), .ZN(n7365) );
  INV_X1 U5179 ( .A(\UUT/branch_rega [4]), .ZN(n7352) );
  INV_X1 U5180 ( .A(\UUT/branch_rega [4]), .ZN(n7348) );
  NOR3_X2 U5181 ( .A1(n451), .A2(n7391), .A3(n203), .ZN(n96) );
  OR2_X1 U5182 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N263 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N264 ) );
  OR2_X1 U5183 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N115 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N116 ) );
  OR2_X1 U5184 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N257 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N258 ) );
  OR2_X1 U5185 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N251 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N252 ) );
  OR2_X1 U5186 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N123 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N124 ) );
  OR2_X1 U5187 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N245 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N246 ) );
  INV_X1 U5188 ( .A(\UUT/Mcontrol/d_jump_type[1] ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N224 ) );
  OR2_X1 U5189 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N106 ), .ZN(\UUT/Mcontrol/st_logic/N107 ) );
  OR2_X1 U5190 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N61 ), .ZN(\UUT/Mcontrol/st_logic/N62 ) );
  OR2_X1 U5191 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N68 ), .ZN(\UUT/Mcontrol/st_logic/N69 ) );
  INV_X1 U5192 ( .A(\UUT/Mcontrol/d_jump_type[1] ), .ZN(
        \UUT/Mcontrol/st_logic/N90 ) );
  OR2_X1 U5193 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N86 ), .ZN(\UUT/Mcontrol/st_logic/N87 ) );
  OR2_X1 U5194 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N74 ), .ZN(\UUT/Mcontrol/st_logic/N75 ) );
  NOR3_X2 U5195 ( .A1(n2591), .A2(\UUT/Mcontrol/Nextpc_decoding/N116 ), .A3(
        n2592), .ZN(n985) );
  NOR2_X2 U5196 ( .A1(n1210), .A2(n499), .ZN(n285) );
  OAI222_X1 U5197 ( .A1(n50), .A2(n94), .B1(n805), .B2(n302), .C1(
        \UUT/Mpath/the_alu/N80 ), .C2(\UUT/Mcontrol/N22 ), .ZN(n3741) );
  NAND2_X2 U5198 ( .A1(\UUT/Mcontrol/N22 ), .A2(n835), .ZN(n94) );
  CLKBUF_X2 U5199 ( .A(n83), .Z(n6340) );
  OAI21_X1 U5200 ( .B1(\UUT/Mpath/the_mult/N227 ), .B2(
        \UUT/Mpath/the_mult/N223 ), .A(\UUT/Mcontrol/N22 ), .ZN(n83) );
  OR3_X1 U5201 ( .A1(\UUT/Mpath/the_shift/N115 ), .A2(
        \UUT/Mpath/the_shift/N118 ), .A3(n1440), .ZN(n6341) );
  INV_X1 U5202 ( .A(n6341), .ZN(n6342) );
  INV_X1 U5203 ( .A(n6341), .ZN(n6343) );
  AND3_X2 U5204 ( .A1(\UUT/Mcontrol/N22 ), .A2(n929), .A3(n5315), .ZN(n117) );
  AND3_X2 U5205 ( .A1(\UUT/Mcontrol/N22 ), .A2(n936), .A3(n5315), .ZN(n105) );
  AND2_X4 U5206 ( .A1(n5886), .A2(n5895), .ZN(n1469) );
  INV_X2 U5207 ( .A(n5455), .ZN(n2116) );
  INV_X4 U5208 ( .A(n5649), .ZN(n1472) );
  AND2_X4 U5209 ( .A1(n5875), .A2(n5876), .ZN(n5631) );
  AND2_X1 U5210 ( .A1(n5879), .A2(n5882), .ZN(n6344) );
  NOR2_X4 U5211 ( .A1(n5884), .A2(\UUT/rs2_addr [3]), .ZN(n5879) );
  AND2_X1 U5212 ( .A1(n5883), .A2(n5877), .ZN(n5882) );
  CLKBUF_X1 U5213 ( .A(n5653), .Z(n6345) );
  CLKBUF_X1 U5214 ( .A(n5653), .Z(n6346) );
  AND3_X4 U5215 ( .A1(\UUT/rs2_addr [4]), .A2(n5877), .A3(n5886), .ZN(n5641)
         );
  AND3_X4 U5216 ( .A1(\UUT/rs2_addr [3]), .A2(\UUT/rs2_addr [4]), .A3(n5882), 
        .ZN(n5646) );
  NAND3_X1 U5217 ( .A1(n6933), .A2(n5878), .A3(n5891), .ZN(n6347) );
  INV_X1 U5218 ( .A(n6347), .ZN(n6348) );
  INV_X1 U5219 ( .A(n6347), .ZN(n6349) );
  NAND2_X4 U5220 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(\UUT/byp_controlB[0] ), 
        .ZN(n5336) );
  INV_X2 U5221 ( .A(n5439), .ZN(n2104) );
  INV_X4 U5222 ( .A(n5633), .ZN(n1455) );
  NAND2_X4 U5223 ( .A1(n5893), .A2(n5890), .ZN(n5654) );
  AND3_X4 U5224 ( .A1(n6266), .A2(n2606), .A3(n6278), .ZN(n2109) );
  AND3_X4 U5225 ( .A1(n5882), .A2(n2090), .A3(n5884), .ZN(n1462) );
  INV_X2 U5226 ( .A(\UUT/N3 ), .ZN(n6322) );
  OR2_X1 U5227 ( .A1(\UUT/N76 ), .A2(\UUT/N77 ), .ZN(\UUT/N3 ) );
  AND4_X2 U5228 ( .A1(\UUT/Mcontrol/N22 ), .A2(n924), .A3(n5315), .A4(n925), 
        .ZN(n121) );
  INV_X2 U5229 ( .A(n877), .ZN(n880) );
  OR2_X2 U5230 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/regfile/N269 ), .ZN(n102) );
  OR2_X4 U5231 ( .A1(\UUT/Mcontrol/bp_logicB/memory_main ), .A2(
        \UUT/Mcontrol/bp_logicB/exec_main ), .ZN(\UUT/byp_controlB[2] ) );
  INV_X2 U5232 ( .A(n688), .ZN(n679) );
  INV_X2 U5233 ( .A(n868), .ZN(n871) );
  INV_X2 U5234 ( .A(n713), .ZN(n704) );
  INV_X2 U5235 ( .A(n856), .ZN(n859) );
  INV_X2 U5236 ( .A(n844), .ZN(n847) );
  INV_X2 U5237 ( .A(n743), .ZN(n734) );
  INV_X2 U5238 ( .A(n768), .ZN(n759) );
  INV_X2 U5239 ( .A(n818), .ZN(n809) );
  INV_X2 U5240 ( .A(n466), .ZN(n455) );
  INV_X2 U5241 ( .A(n793), .ZN(n784) );
  INV_X2 U5242 ( .A(n314), .ZN(n305) );
  INV_X2 U5243 ( .A(n177), .ZN(n169) );
  INV_X2 U5244 ( .A(n160), .ZN(n152) );
  INV_X2 U5245 ( .A(n339), .ZN(n330) );
  INV_X2 U5246 ( .A(n362), .ZN(n353) );
  INV_X2 U5247 ( .A(n143), .ZN(n135) );
  INV_X2 U5248 ( .A(n216), .ZN(n208) );
  INV_X2 U5249 ( .A(n389), .ZN(n380) );
  INV_X2 U5250 ( .A(n413), .ZN(n404) );
  INV_X2 U5251 ( .A(n193), .ZN(n185) );
  INV_X2 U5252 ( .A(n128), .ZN(n114) );
  INV_X2 U5253 ( .A(n437), .ZN(n428) );
  CLKBUF_X1 U5254 ( .A(n124), .Z(n6350) );
  NAND2_X2 U5255 ( .A1(\UUT/Mcontrol/N22 ), .A2(n940), .ZN(n218) );
  INV_X4 U5256 ( .A(n5638), .ZN(n1457) );
  INV_X4 U5257 ( .A(n5444), .ZN(n2105) );
  AND3_X1 U5258 ( .A1(n5877), .A2(n5878), .A3(n5875), .ZN(n6351) );
  INV_X1 U5259 ( .A(n6351), .ZN(n6352) );
  INV_X1 U5260 ( .A(n6351), .ZN(n6353) );
  NAND3_X2 U5261 ( .A1(n5888), .A2(\UUT/rs2_addr [1]), .A3(n5895), .ZN(n5657)
         );
  NAND3_X2 U5262 ( .A1(n5887), .A2(n5890), .A3(\UUT/rs2_addr [1]), .ZN(n5642)
         );
  NOR2_X4 U5263 ( .A1(n5884), .A2(n5877), .ZN(n5887) );
  INV_X2 U5264 ( .A(n997), .ZN(n287) );
  NAND3_X4 U5265 ( .A1(n5877), .A2(n5884), .A3(n5886), .ZN(n1465) );
  INV_X4 U5266 ( .A(n5456), .ZN(n2114) );
  INV_X2 U5267 ( .A(n5650), .ZN(n1468) );
  INV_X4 U5268 ( .A(n5632), .ZN(n1453) );
  INV_X2 U5269 ( .A(n5438), .ZN(n2103) );
  AND2_X4 U5270 ( .A1(n5891), .A2(n5883), .ZN(n5652) );
  AND2_X4 U5271 ( .A1(n5886), .A2(n5887), .ZN(n5640) );
  AND2_X2 U5272 ( .A1(n5888), .A2(n5878), .ZN(n5886) );
  NAND3_X4 U5273 ( .A1(\UUT/rs2_addr [1]), .A2(n5890), .A3(n5895), .ZN(n5655)
         );
  AND2_X2 U5274 ( .A1(n928), .A2(n926), .ZN(n119) );
  NAND3_X1 U5275 ( .A1(n5887), .A2(\UUT/rs2_addr [3]), .A3(n5883), .ZN(n6354)
         );
  INV_X1 U5276 ( .A(n6354), .ZN(n6355) );
  INV_X1 U5277 ( .A(n6354), .ZN(n6356) );
  AND3_X4 U5278 ( .A1(n6266), .A2(\UUT/rs1_addr [0]), .A3(n6262), .ZN(n5441)
         );
  NAND2_X2 U5279 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/Mcontrol/st_logic/N42 ), .ZN(n99) );
  AND3_X4 U5280 ( .A1(n5883), .A2(\UUT/rs2_addr [0]), .A3(n5879), .ZN(n5635)
         );
  NAND3_X2 U5281 ( .A1(\UUT/Mpath/the_mult/N285 ), .A2(n928), .A3(
        \UUT/Mpath/the_mult/N313 ), .ZN(n103) );
  OR2_X1 U5282 ( .A1(\UUT/Mpath/the_mult/m_mul_command[0] ), .A2(
        \UUT/Mpath/the_mult/N284 ), .ZN(\UUT/Mpath/the_mult/N285 ) );
  OR2_X1 U5283 ( .A1(\UUT/Mpath/the_mult/N292 ), .A2(\UUT/Mpath/the_mult/N298 ), .ZN(\UUT/Mpath/the_mult/N313 ) );
  NAND3_X2 U5284 ( .A1(\UUT/Mpath/the_mult/N255 ), .A2(n928), .A3(
        \UUT/Mpath/the_mult/N311 ), .ZN(n115) );
  OR2_X1 U5285 ( .A1(\UUT/Mpath/the_mult/N231 ), .A2(\UUT/Mpath/the_mult/N254 ), .ZN(\UUT/Mpath/the_mult/N255 ) );
  OR2_X1 U5286 ( .A1(\UUT/Mpath/the_mult/N262 ), .A2(\UUT/Mpath/the_mult/N268 ), .ZN(\UUT/Mpath/the_mult/N311 ) );
  NAND3_X4 U5287 ( .A1(\UUT/rs2_addr [1]), .A2(n5887), .A3(n5888), .ZN(n5637)
         );
  NAND3_X4 U5288 ( .A1(n6933), .A2(n5892), .A3(n5893), .ZN(n5647) );
  AND2_X2 U5289 ( .A1(n928), .A2(n934), .ZN(n107) );
  INV_X2 U5290 ( .A(n872), .ZN(n100) );
  NAND2_X2 U5291 ( .A1(\UUT/byp_controlB[2] ), .A2(\UUT/byp_controlB[0] ), 
        .ZN(n101) );
  INV_X2 U5292 ( .A(n48), .ZN(n46) );
  NAND2_X2 U5293 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1098), .ZN(n48) );
  NOR3_X4 U5294 ( .A1(n997), .A2(\UUT/Mpath/N128 ), .A3(n998), .ZN(n320) );
  OR2_X1 U5295 ( .A1(\UUT/Mpath/N112 ), .A2(\UUT/Mpath/N127 ), .ZN(
        \UUT/Mpath/N128 ) );
  INV_X2 U5296 ( .A(n83), .ZN(n125) );
  NOR2_X4 U5297 ( .A1(n1208), .A2(\UUT/Mpath/the_mult/N216 ), .ZN(n291) );
  NOR2_X4 U5298 ( .A1(n6340), .A2(n5430), .ZN(n129) );
  NOR2_X4 U5299 ( .A1(n7382), .A2(n5430), .ZN(n221) );
  NOR2_X4 U5300 ( .A1(n7382), .A2(n5432), .ZN(n220) );
  NOR2_X4 U5301 ( .A1(n6340), .A2(n5432), .ZN(n127) );
  CLKBUF_X2 U5302 ( .A(n293), .Z(n6357) );
  INV_X4 U5303 ( .A(n6358), .ZN(n6359) );
  OR3_X1 U5304 ( .A1(\UUT/regfile/N433 ), .A2(n7392), .A3(n882), .ZN(n6360) );
  INV_X2 U5305 ( .A(n6360), .ZN(n6361) );
  INV_X2 U5306 ( .A(n257), .ZN(n6362) );
  INV_X2 U5307 ( .A(n6361), .ZN(n259) );
  INV_X2 U5308 ( .A(n256), .ZN(n257) );
  OR3_X1 U5309 ( .A1(\UUT/regfile/N421 ), .A2(n7392), .A3(n884), .ZN(n6363) );
  INV_X2 U5310 ( .A(n6363), .ZN(n6364) );
  INV_X2 U5311 ( .A(n261), .ZN(n6365) );
  INV_X2 U5312 ( .A(n6364), .ZN(n255) );
  INV_X2 U5313 ( .A(n260), .ZN(n261) );
  INV_X2 U5314 ( .A(n263), .ZN(n6366) );
  INV_X2 U5315 ( .A(n253), .ZN(n6367) );
  INV_X2 U5316 ( .A(n262), .ZN(n263) );
  INV_X2 U5317 ( .A(n252), .ZN(n253) );
  INV_X2 U5318 ( .A(n251), .ZN(n6368) );
  INV_X2 U5319 ( .A(n265), .ZN(n6369) );
  INV_X2 U5320 ( .A(n250), .ZN(n251) );
  INV_X2 U5321 ( .A(n264), .ZN(n265) );
  INV_X2 U5322 ( .A(n267), .ZN(n6370) );
  INV_X2 U5323 ( .A(n249), .ZN(n6371) );
  INV_X2 U5324 ( .A(n266), .ZN(n267) );
  INV_X2 U5325 ( .A(n248), .ZN(n249) );
  INV_X2 U5326 ( .A(n247), .ZN(n6372) );
  INV_X2 U5327 ( .A(n269), .ZN(n6373) );
  INV_X2 U5328 ( .A(n246), .ZN(n247) );
  INV_X2 U5329 ( .A(n268), .ZN(n269) );
  INV_X2 U5330 ( .A(n271), .ZN(n6374) );
  INV_X2 U5331 ( .A(n245), .ZN(n6375) );
  INV_X2 U5332 ( .A(n270), .ZN(n271) );
  INV_X2 U5333 ( .A(n244), .ZN(n245) );
  INV_X2 U5334 ( .A(n243), .ZN(n6376) );
  INV_X2 U5335 ( .A(n273), .ZN(n6377) );
  INV_X2 U5336 ( .A(n242), .ZN(n243) );
  INV_X2 U5337 ( .A(n272), .ZN(n273) );
  INV_X2 U5338 ( .A(n275), .ZN(n6378) );
  INV_X2 U5339 ( .A(n241), .ZN(n6379) );
  INV_X2 U5340 ( .A(n274), .ZN(n275) );
  INV_X2 U5341 ( .A(n240), .ZN(n241) );
  INV_X2 U5342 ( .A(n239), .ZN(n6380) );
  INV_X2 U5343 ( .A(n277), .ZN(n6381) );
  INV_X2 U5344 ( .A(n238), .ZN(n239) );
  INV_X2 U5345 ( .A(n276), .ZN(n277) );
  INV_X2 U5346 ( .A(n237), .ZN(n6382) );
  INV_X2 U5347 ( .A(n281), .ZN(n6383) );
  INV_X2 U5348 ( .A(n279), .ZN(n6384) );
  INV_X2 U5349 ( .A(n233), .ZN(n6385) );
  INV_X2 U5350 ( .A(n236), .ZN(n237) );
  INV_X2 U5351 ( .A(n280), .ZN(n281) );
  INV_X2 U5352 ( .A(n278), .ZN(n279) );
  INV_X2 U5353 ( .A(n232), .ZN(n233) );
  OR3_X1 U5354 ( .A1(\UUT/regfile/N342 ), .A2(n7391), .A3(n883), .ZN(n6386) );
  INV_X2 U5355 ( .A(n6386), .ZN(n6387) );
  OR3_X1 U5356 ( .A1(\UUT/regfile/N367 ), .A2(n7391), .A3(n883), .ZN(n6388) );
  INV_X2 U5357 ( .A(n6388), .ZN(n6389) );
  INV_X2 U5358 ( .A(n231), .ZN(n6390) );
  INV_X2 U5359 ( .A(n283), .ZN(n6391) );
  INV_X2 U5360 ( .A(n6387), .ZN(n227) );
  INV_X2 U5361 ( .A(n6389), .ZN(n235) );
  INV_X2 U5362 ( .A(n230), .ZN(n231) );
  INV_X2 U5363 ( .A(n282), .ZN(n283) );
  OR3_X1 U5364 ( .A1(\UUT/regfile/N330 ), .A2(n7391), .A3(n881), .ZN(n6392) );
  INV_X2 U5365 ( .A(n6392), .ZN(n6393) );
  OR3_X1 U5366 ( .A1(\UUT/regfile/N348 ), .A2(n7391), .A3(n884), .ZN(n6394) );
  INV_X2 U5367 ( .A(n6394), .ZN(n6395) );
  INV_X2 U5368 ( .A(n225), .ZN(n6396) );
  AOI211_X4 U5369 ( .C1(n573), .C2(n498), .A(n499), .B(n574), .ZN(n561) );
  INV_X2 U5370 ( .A(n6393), .ZN(n223) );
  INV_X2 U5371 ( .A(n6395), .ZN(n229) );
  INV_X2 U5372 ( .A(n224), .ZN(n225) );
  AOI211_X4 U5373 ( .C1(n497), .C2(n498), .A(n499), .B(n500), .ZN(n485) );
  AOI211_X4 U5374 ( .C1(n548), .C2(n498), .A(n499), .B(n549), .ZN(n536) );
  AOI211_X4 U5375 ( .C1(n524), .C2(n498), .A(n499), .B(n525), .ZN(n512) );
  AOI211_X4 U5376 ( .C1(n597), .C2(n498), .A(n499), .B(n598), .ZN(n585) );
  CLKBUF_X2 U5377 ( .A(n289), .Z(n6397) );
  AOI211_X4 U5378 ( .C1(n620), .C2(n498), .A(n499), .B(n621), .ZN(n608) );
  AOI211_X4 U5379 ( .C1(n667), .C2(n498), .A(n499), .B(n668), .ZN(n655) );
  AOI211_X4 U5380 ( .C1(n643), .C2(n498), .A(n499), .B(n644), .ZN(n631) );
  INV_X2 U5381 ( .A(n7169), .ZN(\UUT/Mcontrol/Operation_decoding32/N2060 ) );
  AOI21_X1 U5382 ( .B1(\UUT/Mcontrol/Nextpc_decoding/N32 ), .B2(
        \UUT/Mcontrol/Nextpc_decoding/N230 ), .A(
        \UUT/Mcontrol/Nextpc_decoding/N236 ), .ZN(n6256) );
  INV_X4 U5383 ( .A(n7341), .ZN(n6017) );
  INV_X2 U5384 ( .A(\UUT/Mcontrol/d_instr [26]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1922 ) );
  INV_X2 U5385 ( .A(\UUT/rs1_addr [3]), .ZN(n6275) );
  NOR2_X2 U5386 ( .A1(n5760), .A2(n6279), .ZN(\UUT/rs1_addr [3]) );
  AND4_X2 U5387 ( .A1(n2156), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(n5320)
         );
  NAND2_X1 U5388 ( .A1(n1006), .A2(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
        .ZN(n6827) );
  AND2_X1 U5389 ( .A1(\UUT/jar_in [16]), .A2(n6867), .ZN(n6828) );
  AND2_X1 U5390 ( .A1(n300), .A2(\UUT/branch_rega [16]), .ZN(n6829) );
  AND2_X1 U5391 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [16]), .A2(n301), .ZN(
        n6830) );
  NOR3_X1 U5392 ( .A1(n6828), .A2(n6829), .A3(n6830), .ZN(n449) );
  NOR2_X1 U5393 ( .A1(n556), .A2(\UUT/Mcontrol/Nextpc_decoding/N125 ), .ZN(
        n300) );
  INV_X1 U5394 ( .A(n7356), .ZN(n6831) );
  NAND2_X1 U5395 ( .A1(n6832), .A2(n6833), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N200 ) );
  AND2_X1 U5396 ( .A1(n7261), .A2(n7260), .ZN(n6832) );
  NOR2_X1 U5397 ( .A1(n6843), .A2(n6831), .ZN(n6833) );
  OAI222_X2 U5398 ( .A1(n5967), .A2(n5468), .B1(n5968), .B2(n5525), .C1(n5969), 
        .C2(n5466), .ZN(n5966) );
  AND2_X4 U5399 ( .A1(\UUT/Mpath/the_alu/N486 ), .A2(n2230), .ZN(n6834) );
  INV_X4 U5400 ( .A(n6834), .ZN(n1304) );
  NOR2_X1 U5401 ( .A1(n7165), .A2(n7161), .ZN(n7219) );
  AND2_X2 U5402 ( .A1(n1334), .A2(n1335), .ZN(n6100) );
  BUF_X1 U5403 ( .A(\UUT/Mcontrol/d_sampled_finstr [30]), .Z(n7192) );
  OR2_X1 U5404 ( .A1(\UUT/Alu_command[OP][4] ), .A2(\UUT/Alu_command[OP][5] ), 
        .ZN(\UUT/Mpath/the_alu/N517 ) );
  OR2_X1 U5405 ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(\UUT/Alu_command[OP][5] ), 
        .ZN(\UUT/Mpath/the_alu/N505 ) );
  OR2_X1 U5406 ( .A1(\UUT/Mpath/the_alu/N453 ), .A2(\UUT/Alu_command[OP][5] ), 
        .ZN(\UUT/Mpath/the_alu/N511 ) );
  OAI22_X2 U5407 ( .A1(\UUT/Mpath/the_alu/N520 ), .A2(n2240), .B1(
        \UUT/Mpath/the_alu/N526 ), .B2(\UUT/Mpath/the_alu/N468 ), .ZN(n1216)
         );
  AND2_X2 U5408 ( .A1(n6878), .A2(\UUT/Mcontrol/st_logic/N108 ), .ZN(n6877) );
  INV_X2 U5409 ( .A(\UUT/Mcontrol/st_logic/N10 ), .ZN(n1013) );
  CLKBUF_X1 U5410 ( .A(\UUT/Mpath/the_mult/x_mult_out[30] ), .Z(n6835) );
  AND3_X2 U5411 ( .A1(n6837), .A2(n6836), .A3(n7150), .ZN(n6034) );
  NOR2_X1 U5412 ( .A1(n7152), .A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
        .ZN(n6836) );
  NOR2_X1 U5413 ( .A1(n1373), .A2(n7208), .ZN(n6837) );
  OR2_X2 U5414 ( .A1(\UUT/Mcontrol/N22 ), .A2(n930), .ZN(n6838) );
  NAND2_X1 U5415 ( .A1(n6838), .A2(n1201), .ZN(n4310) );
  AOI222_X2 U5416 ( .A1(n6397), .A2(n901), .B1(n291), .B2(n902), .C1(
        \UUT/Mpath/the_mult/x_mult_out[25] ), .C2(n6357), .ZN(n900) );
  NAND2_X2 U5417 ( .A1(n7338), .A2(n7339), .ZN(n7238) );
  INV_X1 U5418 ( .A(n1203), .ZN(n86) );
  NAND2_X2 U5419 ( .A1(n7372), .A2(n7371), .ZN(n7222) );
  OAI222_X4 U5420 ( .A1(n5399), .A2(n5432), .B1(n5431), .B2(n387), .C1(n5397), 
        .C2(n5430), .ZN(\UUT/branch_rega [19]) );
  INV_X1 U5421 ( .A(n6034), .ZN(n6037) );
  OAI22_X2 U5422 ( .A1(n5776), .A2(n6030), .B1(n6213), .B2(n7179), .ZN(n6212)
         );
  OAI21_X2 U5423 ( .B1(n5915), .B2(n5936), .A(n6890), .ZN(n6050) );
  NAND2_X2 U5424 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1933 ), .A2(n7118), 
        .ZN(n7104) );
  OAI222_X1 U5425 ( .A1(n98), .A2(n5332), .B1(n100), .B2(n101), .C1(n5359), 
        .C2(n102), .ZN(n6840) );
  INV_X8 U5426 ( .A(n6841), .ZN(n6842) );
  OAI222_X1 U5427 ( .A1(n98), .A2(n99), .B1(n100), .B2(n101), .C1(n5359), .C2(
        n102), .ZN(n93) );
  INV_X1 U5428 ( .A(n7090), .ZN(n7091) );
  OR2_X1 U5429 ( .A1(\UUT/branch_rega [18]), .A2(\UUT/branch_rega [17]), .ZN(
        n7376) );
  INV_X1 U5430 ( .A(n7376), .ZN(n7377) );
  OR2_X1 U5431 ( .A1(n6844), .A2(\UUT/branch_rega [24]), .ZN(n6843) );
  INV_X1 U5432 ( .A(n7346), .ZN(n6844) );
  NAND2_X1 U5433 ( .A1(n7360), .A2(n7361), .ZN(n6845) );
  NAND2_X1 U5434 ( .A1(n1294), .A2(n7362), .ZN(n6846) );
  AND2_X1 U5435 ( .A1(n6845), .A2(n6846), .ZN(n7359) );
  OR2_X1 U5436 ( .A1(n477), .A2(n296), .ZN(n6847) );
  OR2_X1 U5437 ( .A1(n297), .A2(n2663), .ZN(n6848) );
  NAND3_X1 U5438 ( .A1(n6847), .A2(n6848), .A3(n478), .ZN(n3222) );
  INV_X1 U5439 ( .A(n6111), .ZN(n7360) );
  INV_X1 U5440 ( .A(n5466), .ZN(n7361) );
  OAI222_X1 U5441 ( .A1(n7359), .A2(n5332), .B1(n5356), .B2(n5334), .C1(n5357), 
        .C2(n5336), .ZN(\UUT/branch_regb [31]) );
  AOI221_X1 U5442 ( .B1(n479), .B2(n480), .C1(n6892), .C2(n482), .A(n456), 
        .ZN(n477) );
  OAI221_X1 U5443 ( .B1(n6110), .B2(n286), .C1(n6111), .C2(n287), .A(n1204), 
        .ZN(n878) );
  NOR2_X2 U5444 ( .A1(n7121), .A2(n6955), .ZN(n1204) );
  NOR2_X1 U5445 ( .A1(n984), .A2(n556), .ZN(n6867) );
  INV_X4 U5446 ( .A(\UUT/branch_rega [22]), .ZN(n7356) );
  NOR2_X1 U5447 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N205 ), .A2(
        \UUT/branch_rega [16]), .ZN(n6928) );
  NAND2_X1 U5448 ( .A1(n6897), .A2(n6898), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N205 ) );
  OR2_X1 U5449 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2016 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2017 ) );
  INV_X1 U5450 ( .A(\UUT/Mcontrol/Operation_decoding32/N1973 ), .ZN(n6853) );
  AND2_X2 U5451 ( .A1(n6002), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .ZN(n6849) );
  INV_X2 U5452 ( .A(n6849), .ZN(n6134) );
  BUF_X2 U5453 ( .A(n6849), .Z(n6995) );
  BUF_X2 U5454 ( .A(n6995), .Z(n6996) );
  OR2_X2 U5455 ( .A1(n6851), .A2(n6903), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2066 ) );
  OR2_X2 U5456 ( .A1(n7030), .A2(\UUT/Mcontrol/Operation_decoding32/N1989 ), 
        .ZN(n6903) );
  BUF_X1 U5457 ( .A(n7237), .Z(n6850) );
  OR2_X1 U5458 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2050 ), .A2(n7216), 
        .ZN(n6893) );
  OR2_X2 U5459 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2050 ), .A2(
        \UUT/Mcontrol/d_instr [29]), .ZN(n6851) );
  CLKBUF_X1 U5460 ( .A(n6888), .Z(n6852) );
  BUF_X1 U5461 ( .A(n7150), .Z(n6879) );
  AND2_X1 U5462 ( .A1(n6881), .A2(n7154), .ZN(n6854) );
  AND2_X2 U5463 ( .A1(n6881), .A2(n6853), .ZN(n7070) );
  OR2_X2 U5464 ( .A1(n7192), .A2(n7201), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1947 ) );
  INV_X1 U5465 ( .A(n6852), .ZN(n5909) );
  INV_X1 U5466 ( .A(n7216), .ZN(\UUT/Mcontrol/d_instr [29]) );
  CLKBUF_X1 U5467 ( .A(\UUT/Mcontrol/d_instr [31]), .Z(n6855) );
  AND2_X2 U5468 ( .A1(n6882), .A2(\UUT/Mcontrol/Operation_decoding32/N1877 ), 
        .ZN(n6856) );
  NAND2_X1 U5469 ( .A1(n6856), .A2(n6857), .ZN(n7118) );
  AND2_X1 U5470 ( .A1(n6858), .A2(n2765), .ZN(n6857) );
  INV_X1 U5471 ( .A(\UUT/Mcontrol/Operation_decoding32/N1922 ), .ZN(n6858) );
  NOR2_X2 U5472 ( .A1(n7222), .A2(n6859), .ZN(n7332) );
  NAND2_X1 U5473 ( .A1(n6860), .A2(n7312), .ZN(n6859) );
  NOR2_X1 U5474 ( .A1(n7223), .A2(n7001), .ZN(n6860) );
  AND2_X1 U5475 ( .A1(n6867), .A2(\UUT/jar_in [23]), .ZN(n6861) );
  NOR2_X1 U5476 ( .A1(n6861), .A2(n6862), .ZN(n7149) );
  OR2_X1 U5477 ( .A1(n6863), .A2(n7340), .ZN(n6862) );
  INV_X1 U5478 ( .A(n7326), .ZN(n6863) );
  AND2_X1 U5479 ( .A1(\UUT/Mpath/the_alu/sum[20] ), .A2(n7213), .ZN(n6864) );
  AND2_X1 U5480 ( .A1(\UUT/Mpath/the_alu/N137 ), .A2(n6834), .ZN(n6865) );
  AND2_X1 U5481 ( .A1(n1218), .A2(n1273), .ZN(n6866) );
  NOR3_X1 U5482 ( .A1(n6864), .A2(n6865), .A3(n6866), .ZN(n1272) );
  NOR2_X1 U5483 ( .A1(n984), .A2(n556), .ZN(n299) );
  NOR2_X2 U5484 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2015 ), .A2(n6939), 
        .ZN(n6970) );
  NOR2_X2 U5485 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1947 ), .A2(n6906), 
        .ZN(n7064) );
  CLKBUF_X1 U5486 ( .A(n6874), .Z(n6869) );
  OR2_X2 U5487 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2050 ), .A2(
        \UUT/Mcontrol/d_instr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2081 ) );
  CLKBUF_X1 U5488 ( .A(n5900), .Z(n6868) );
  NOR2_X1 U5489 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1965 ), .A2(n6881), 
        .ZN(n6882) );
  NAND2_X1 U5490 ( .A1(n7185), .A2(n6997), .ZN(n6870) );
  INV_X2 U5491 ( .A(n6870), .ZN(\UUT/Mcontrol/Operation_decoding32/N2043 ) );
  NAND2_X1 U5492 ( .A1(n6974), .A2(n6975), .ZN(n6871) );
  INV_X1 U5493 ( .A(n6879), .ZN(n6872) );
  OR2_X1 U5494 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2016 ), .A2(n7111), 
        .ZN(n7150) );
  NAND2_X1 U5495 ( .A1(n7172), .A2(\UUT/Mcontrol/Operation_decoding32/N2066 ), 
        .ZN(n6873) );
  NAND2_X1 U5496 ( .A1(n7172), .A2(\UUT/Mcontrol/Operation_decoding32/N2066 ), 
        .ZN(n1373) );
  OR2_X1 U5497 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2002 ), .A2(n7216), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1984 ) );
  NOR2_X1 U5498 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2015 ), .A2(n7044), 
        .ZN(n6874) );
  INV_X4 U5499 ( .A(n2764), .ZN(n7044) );
  INV_X1 U5500 ( .A(n7377), .ZN(n6896) );
  OAI222_X4 U5501 ( .A1(n5405), .A2(n5432), .B1(n5431), .B2(n435), .C1(n5403), 
        .C2(n5430), .ZN(\UUT/branch_rega [17]) );
  OR2_X2 U5502 ( .A1(n7216), .A2(\UUT/Mcontrol/d_instr [28]), .ZN(n6906) );
  OR2_X2 U5503 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1977 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1978 ) );
  NAND2_X1 U5504 ( .A1(n7028), .A2(n7029), .ZN(n6875) );
  NAND2_X1 U5505 ( .A1(n7028), .A2(n7029), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1994 ) );
  NOR2_X2 U5506 ( .A1(\UUT/Mcontrol/st_logic/N112 ), .A2(
        \UUT/Mcontrol/st_logic/N96 ), .ZN(n6876) );
  AND2_X1 U5507 ( .A1(n6876), .A2(\UUT/Mcontrol/st_logic/N101 ), .ZN(n6878) );
  OR2_X2 U5508 ( .A1(n6895), .A2(n6939), .ZN(n6894) );
  NOR2_X1 U5509 ( .A1(n6873), .A2(n7208), .ZN(n6880) );
  NOR2_X2 U5510 ( .A1(n6893), .A2(n6894), .ZN(n7185) );
  AND2_X2 U5511 ( .A1(n7349), .A2(n7350), .ZN(n7366) );
  AND2_X2 U5512 ( .A1(n7331), .A2(n7332), .ZN(n7350) );
  OAI222_X4 U5513 ( .A1(n5390), .A2(n5432), .B1(n5431), .B2(n337), .C1(n5388), 
        .C2(n5430), .ZN(\UUT/branch_rega [21]) );
  AOI21_X1 U5514 ( .B1(n6251), .B2(n6252), .A(n6253), .ZN(n6250) );
  INV_X1 U5515 ( .A(\UUT/Mcontrol/st_logic/branch_uses_main_exe_result ), .ZN(
        \UUT/Mcontrol/st_logic/N41 ) );
  INV_X1 U5516 ( .A(\UUT/Mcontrol/st_logic/branchmul_stall ), .ZN(
        \UUT/Mcontrol/st_logic/N14 ) );
  INV_X1 U5517 ( .A(\UUT/Mcontrol/Operation_decoding32/N1921 ), .ZN(n6881) );
  OR2_X2 U5518 ( .A1(n6873), .A2(n6892), .ZN(n7051) );
  OR2_X1 U5519 ( .A1(n7044), .A2(\UUT/Mcontrol/d_instr [26]), .ZN(n6883) );
  NOR2_X1 U5520 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N134 ), .A2(
        \UUT/branch_rega [22]), .ZN(n6884) );
  NAND2_X1 U5521 ( .A1(n6884), .A2(n6885), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N137 ) );
  AND2_X1 U5522 ( .A1(n6886), .A2(n7367), .ZN(n6885) );
  INV_X1 U5523 ( .A(\UUT/branch_rega [20]), .ZN(n6886) );
  INV_X1 U5524 ( .A(n7164), .ZN(n6887) );
  AND2_X2 U5525 ( .A1(n6032), .A2(n7008), .ZN(n6888) );
  AND2_X1 U5526 ( .A1(n6970), .A2(n6889), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2025 ) );
  AND2_X1 U5527 ( .A1(n7044), .A2(n2763), .ZN(n6889) );
  CLKBUF_X1 U5528 ( .A(n6135), .Z(n6890) );
  NOR2_X1 U5529 ( .A1(n7180), .A2(n6904), .ZN(n6135) );
  AND4_X1 U5530 ( .A1(n2292), .A2(n2293), .A3(n2294), .A4(n2295), .ZN(n337) );
  INV_X1 U5531 ( .A(\UUT/branch_rega [21]), .ZN(n7367) );
  AND3_X4 U5532 ( .A1(\UUT/rs1_addr [1]), .A2(\UUT/rs1_addr [0]), .A3(n6258), 
        .ZN(n5436) );
  OR2_X2 U5533 ( .A1(n7154), .A2(\UUT/Mcontrol/Operation_decoding32/N2083 ), 
        .ZN(n6891) );
  AND2_X2 U5534 ( .A1(n1364), .A2(n1365), .ZN(n5990) );
  NOR2_X4 U5535 ( .A1(n7370), .A2(\UUT/rs1_addr [0]), .ZN(n6259) );
  NAND3_X4 U5536 ( .A1(n6273), .A2(\UUT/rs1_addr [4]), .A3(n6259), .ZN(n5449)
         );
  AND2_X4 U5537 ( .A1(n6258), .A2(n6259), .ZN(n5437) );
  AND2_X4 U5538 ( .A1(n6259), .A2(n6267), .ZN(n6276) );
  NAND2_X1 U5539 ( .A1(n6970), .A2(n6971), .ZN(n7059) );
  OR2_X1 U5540 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1955 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1956 ) );
  AND2_X1 U5541 ( .A1(n7154), .A2(\UUT/Mcontrol/Operation_decoding32/N1921 ), 
        .ZN(n6971) );
  NOR2_X1 U5542 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2088 ), .ZN(n7014) );
  CLKBUF_X1 U5543 ( .A(n7208), .Z(n6892) );
  OR2_X2 U5544 ( .A1(n1124), .A2(n7169), .ZN(n7208) );
  INV_X1 U5545 ( .A(\UUT/Mcontrol/Operation_decoding32/N1921 ), .ZN(n6895) );
  NOR2_X1 U5546 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N200 ), .A2(
        \UUT/branch_rega [21]), .ZN(n6897) );
  NOR2_X1 U5547 ( .A1(n7309), .A2(n6896), .ZN(n6898) );
  NOR2_X2 U5548 ( .A1(n7219), .A2(n7218), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N32 ) );
  INV_X2 U5549 ( .A(n2112), .ZN(n6899) );
  INV_X1 U5550 ( .A(n6899), .ZN(n6900) );
  INV_X2 U5551 ( .A(n6899), .ZN(n6902) );
  INV_X4 U5552 ( .A(n6899), .ZN(n6901) );
  INV_X2 U5553 ( .A(n194), .ZN(n184) );
  NOR2_X1 U5554 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1962 ), .ZN(n6904) );
  NAND2_X1 U5555 ( .A1(n6905), .A2(n2765), .ZN(n7073) );
  NOR2_X1 U5556 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1947 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1877 ), .ZN(n6905) );
  CLKBUF_X1 U5557 ( .A(\UUT/branch_rega [29]), .Z(n7178) );
  OR2_X2 U5558 ( .A1(\UUT/branch_rega [29]), .A2(\UUT/branch_rega [28]), .ZN(
        n7186) );
  OAI21_X2 U5559 ( .B1(n7203), .B2(n2260), .A(n2554), .ZN(\UUT/break_code[5] )
         );
  OAI21_X2 U5560 ( .B1(n6071), .B2(n2556), .A(n6868), .ZN(n2260) );
  OAI21_X1 U5561 ( .B1(n5915), .B2(n5936), .A(n6890), .ZN(n6908) );
  OAI21_X1 U5562 ( .B1(n5915), .B2(n5936), .A(n6890), .ZN(n6907) );
  OR2_X1 U5563 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N127 ), .A2(n7178), .ZN(
        n6909) );
  NOR2_X1 U5564 ( .A1(n6909), .A2(n6910), .ZN(n7156) );
  OR2_X1 U5565 ( .A1(n6911), .A2(n7077), .ZN(n6910) );
  INV_X1 U5566 ( .A(n7045), .ZN(n6911) );
  INV_X1 U5567 ( .A(n6999), .ZN(n6912) );
  NOR2_X1 U5568 ( .A1(n7023), .A2(n6913), .ZN(n7355) );
  NAND2_X1 U5569 ( .A1(n7353), .A2(n6912), .ZN(n6913) );
  NOR3_X2 U5570 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2001 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2007 ), .A3(
        \UUT/Mcontrol/Operation_decoding32/N1995 ), .ZN(n5913) );
  AND2_X2 U5571 ( .A1(\UUT/rs1_addr [3]), .A2(\UUT/rs1_addr [2]), .ZN(n6273)
         );
  OR2_X2 U5572 ( .A1(n7192), .A2(n7201), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1965 ) );
  AND2_X1 U5573 ( .A1(n7015), .A2(n7016), .ZN(n7180) );
  INV_X2 U5574 ( .A(n5892), .ZN(\UUT/rs2_addr [3]) );
  OR2_X2 U5575 ( .A1(\UUT/branch_rega [20]), .A2(\UUT/branch_rega [21]), .ZN(
        n7266) );
  INV_X1 U5576 ( .A(n5987), .ZN(n5388) );
  AOI22_X2 U5577 ( .A1(n107), .A2(n108), .B1(\UUT/Mpath/the_mult/Mad_out [63]), 
        .B2(n109), .ZN(n106) );
  AND4_X2 U5578 ( .A1(n1913), .A2(n1914), .A3(n1915), .A4(n1916), .ZN(n5359)
         );
  INV_X8 U5579 ( .A(n6914), .ZN(n6915) );
  INV_X1 U5580 ( .A(n7275), .ZN(n6916) );
  NAND2_X1 U5581 ( .A1(n6917), .A2(n6918), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N134 ) );
  AND2_X1 U5582 ( .A1(n7277), .A2(n7276), .ZN(n6917) );
  NOR2_X2 U5583 ( .A1(n7299), .A2(n6916), .ZN(n6918) );
  AND3_X2 U5584 ( .A1(n7375), .A2(n7370), .A3(n6258), .ZN(n6919) );
  INV_X32 U5585 ( .A(n6919), .ZN(n5434) );
  AND4_X1 U5586 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n5356)
         );
  NOR2_X4 U5587 ( .A1(n6933), .A2(\UUT/rs2_addr [1]), .ZN(n5883) );
  AND2_X2 U5588 ( .A1(n6921), .A2(n6922), .ZN(n6920) );
  NAND2_X1 U5589 ( .A1(\UUT/Mcontrol/st_logic/N45 ), .A2(
        \UUT/Mcontrol/st_logic/N46 ), .ZN(n6921) );
  NAND2_X1 U5590 ( .A1(\UUT/Mcontrol/st_logic/N50 ), .A2(
        \UUT/Mcontrol/st_logic/N51 ), .ZN(n6922) );
  INV_X2 U5591 ( .A(n5627), .ZN(n6923) );
  INV_X1 U5592 ( .A(n6923), .ZN(n6924) );
  INV_X4 U5593 ( .A(n6923), .ZN(n6925) );
  NOR4_X1 U5594 ( .A1(n2212), .A2(n2213), .A3(n2214), .A4(n2215), .ZN(n2211)
         );
  NAND3_X2 U5595 ( .A1(n6271), .A2(\UUT/rs1_addr [1]), .A3(n6278), .ZN(n5463)
         );
  NAND3_X2 U5596 ( .A1(\UUT/rs1_addr [1]), .A2(n6270), .A3(n6271), .ZN(n5443)
         );
  INV_X1 U5597 ( .A(\UUT/Mcontrol/st_logic/N76 ), .ZN(
        \UUT/Mcontrol/st_logic/N77 ) );
  OR2_X1 U5598 ( .A1(\UUT/Mcontrol/d_jump_type[0] ), .A2(
        \UUT/Mcontrol/st_logic/N75 ), .ZN(\UUT/Mcontrol/st_logic/N76 ) );
  AND2_X2 U5599 ( .A1(n6262), .A2(n6265), .ZN(n5442) );
  AND3_X4 U5600 ( .A1(\UUT/rs1_addr [4]), .A2(n7375), .A3(n6269), .ZN(n5447)
         );
  INV_X1 U5601 ( .A(\UUT/Mcontrol/st_logic/N82 ), .ZN(
        \UUT/Mcontrol/st_logic/N83 ) );
  OR2_X1 U5602 ( .A1(\UUT/Mcontrol/st_logic/N65 ), .A2(
        \UUT/Mcontrol/st_logic/N81 ), .ZN(\UUT/Mcontrol/st_logic/N82 ) );
  AND3_X4 U5603 ( .A1(\UUT/rs2_addr [1]), .A2(\UUT/rs2_addr [0]), .A3(n5875), 
        .ZN(n5630) );
  AND2_X2 U5604 ( .A1(n5879), .A2(n6933), .ZN(n5875) );
  NAND2_X4 U5605 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [20]), .ZN(n5884) );
  OR2_X4 U5606 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1893 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1899 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1873 ) );
  INV_X2 U5607 ( .A(n5884), .ZN(\UUT/rs2_addr [4]) );
  OR2_X4 U5608 ( .A1(\UUT/BYP_BRANCH_MUXB/N4 ), .A2(\UUT/regfile/N269 ), .ZN(
        n5334) );
  BUF_X2 U5609 ( .A(n7237), .Z(n7205) );
  OR2_X1 U5610 ( .A1(n7237), .A2(n7228), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1889 ) );
  OR2_X2 U5611 ( .A1(n7025), .A2(\UUT/Mcontrol/Operation_decoding32/N1952 ), 
        .ZN(n5936) );
  NAND2_X1 U5612 ( .A1(n5948), .A2(n6872), .ZN(n6927) );
  AND2_X2 U5613 ( .A1(n6927), .A2(n6880), .ZN(n6038) );
  NAND2_X1 U5614 ( .A1(n6928), .A2(n6929), .ZN(n7165) );
  AND2_X1 U5615 ( .A1(n6987), .A2(n7308), .ZN(n6929) );
  CLKBUF_X1 U5616 ( .A(n301), .Z(n6930) );
  INV_X1 U5617 ( .A(n983), .ZN(n6931) );
  INV_X2 U5618 ( .A(n6931), .ZN(n6932) );
  AND2_X2 U5619 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1873 ), .A2(n5896), 
        .ZN(n6933) );
  INV_X4 U5620 ( .A(n6933), .ZN(\UUT/rs2_addr [2]) );
  INV_X4 U5621 ( .A(\UUT/branch_rega [8]), .ZN(n7282) );
  INV_X4 U5622 ( .A(\UUT/branch_rega [8]), .ZN(n7304) );
  OR2_X2 U5623 ( .A1(\UUT/branch_rega [8]), .A2(\UUT/branch_rega [7]), .ZN(
        n7378) );
  INV_X4 U5624 ( .A(\UUT/branch_rega [12]), .ZN(n7347) );
  INV_X4 U5625 ( .A(\UUT/branch_rega [12]), .ZN(n7311) );
  INV_X2 U5626 ( .A(n5643), .ZN(n6934) );
  INV_X1 U5627 ( .A(n6934), .ZN(n6935) );
  INV_X2 U5628 ( .A(n6934), .ZN(n6936) );
  AND2_X4 U5629 ( .A1(n983), .A2(n297), .ZN(n301) );
  INV_X8 U5630 ( .A(n6937), .ZN(n6938) );
  BUF_X4 U5631 ( .A(\UUT/Mcontrol/d_instr [28]), .Z(n6939) );
  NOR2_X1 U5632 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N142 ), .A2(
        \UUT/branch_rega [14]), .ZN(n6940) );
  AND2_X1 U5633 ( .A1(n6940), .A2(n6941), .ZN(n7302) );
  AND2_X1 U5634 ( .A1(n6942), .A2(n7344), .ZN(n6941) );
  INV_X1 U5635 ( .A(n7010), .ZN(n6942) );
  NOR2_X1 U5636 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1919 ), .ZN(n6943) );
  OR2_X1 U5637 ( .A1(n7044), .A2(\UUT/Mcontrol/Operation_decoding32/N1918 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1919 ) );
  OR2_X1 U5638 ( .A1(n5492), .A2(n286), .ZN(n6944) );
  OR2_X1 U5639 ( .A1(n5491), .A2(n287), .ZN(n6945) );
  NAND3_X1 U5640 ( .A1(n6944), .A2(n6945), .A3(n908), .ZN(n161) );
  NAND2_X4 U5641 ( .A1(n6397), .A2(n909), .ZN(n6946) );
  NAND2_X1 U5642 ( .A1(n291), .A2(n910), .ZN(n6947) );
  NAND2_X1 U5643 ( .A1(\UUT/Mpath/the_mult/x_mult_out[27] ), .A2(n6357), .ZN(
        n6948) );
  AND3_X1 U5644 ( .A1(n6946), .A2(n6947), .A3(n6948), .ZN(n908) );
  INV_X1 U5645 ( .A(n161), .ZN(n151) );
  OR2_X1 U5646 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N262 ) );
  OR2_X1 U5647 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N98 ) );
  OR2_X1 U5648 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N60 ) );
  OR2_X1 U5649 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N114 ) );
  OR2_X1 U5650 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N244 ) );
  OR2_X1 U5651 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N232 ) );
  OR2_X1 U5652 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N250 ) );
  OR2_X1 U5653 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N238 ) );
  OR2_X1 U5654 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N226 ) );
  OR2_X1 U5655 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N256 ) );
  OR2_X1 U5656 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/Nextpc_decoding/N122 ) );
  OR2_X1 U5657 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N67 ) );
  OR2_X1 U5658 ( .A1(\UUT/Mcontrol/st_logic/N103 ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N105 ) );
  BUF_X1 U5659 ( .A(\UUT/Mcontrol/Operation_decoding32/N1989 ), .Z(n7033) );
  OR2_X1 U5660 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N85 ) );
  OR2_X1 U5661 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N92 ) );
  OR2_X1 U5662 ( .A1(n5484), .A2(n286), .ZN(n6949) );
  OR2_X1 U5663 ( .A1(n5483), .A2(n287), .ZN(n6950) );
  NAND3_X1 U5664 ( .A1(n6949), .A2(n6950), .A3(n912), .ZN(n144) );
  AND2_X1 U5665 ( .A1(n6397), .A2(n913), .ZN(n6951) );
  AND2_X1 U5666 ( .A1(n291), .A2(n914), .ZN(n6952) );
  AND2_X2 U5667 ( .A1(\UUT/Mpath/the_mult/x_mult_out[28] ), .A2(n6357), .ZN(
        n6953) );
  NOR3_X2 U5668 ( .A1(n6951), .A2(n6952), .A3(n6953), .ZN(n912) );
  INV_X1 U5669 ( .A(n1413), .ZN(n5484) );
  INV_X1 U5670 ( .A(n144), .ZN(n134) );
  OR2_X2 U5671 ( .A1(\UUT/Mcontrol/d_instr [31]), .A2(n7205), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1977 ) );
  OAI21_X2 U5672 ( .B1(n6037), .B2(n6888), .A(n6038), .ZN(n5959) );
  OR2_X1 U5673 ( .A1(\UUT/Mcontrol/d_jump_type[1] ), .A2(
        \UUT/Mcontrol/st_logic/N80 ), .ZN(\UUT/Mcontrol/st_logic/N81 ) );
  OR2_X1 U5674 ( .A1(\UUT/Mcontrol/st_logic/N58 ), .A2(
        \UUT/Mcontrol/st_logic/N79 ), .ZN(\UUT/Mcontrol/st_logic/N80 ) );
  NAND3_X2 U5675 ( .A1(n6996), .A2(n7019), .A3(n5920), .ZN(n5924) );
  NOR2_X1 U5676 ( .A1(n7119), .A2(n7120), .ZN(n6954) );
  INV_X1 U5677 ( .A(n6954), .ZN(n6955) );
  AND2_X1 U5678 ( .A1(\UUT/Mpath/the_mult/x_mult_out[31] ), .A2(n6357), .ZN(
        n7121) );
  CLKBUF_X1 U5679 ( .A(n6017), .Z(n6956) );
  OAI222_X4 U5680 ( .A1(n6017), .A2(n5906), .B1(n7069), .B2(n5327), .C1(n7203), 
        .C2(n7021), .ZN(n6180) );
  OAI222_X4 U5681 ( .A1(n6956), .A2(n5897), .B1(n7168), .B2(n5776), .C1(n7021), 
        .C2(n5762), .ZN(n6283) );
  OAI222_X4 U5682 ( .A1(n6956), .A2(n5896), .B1(n7168), .B2(n5762), .C1(n7021), 
        .C2(n5905), .ZN(n6224) );
  OR2_X1 U5683 ( .A1(n5500), .A2(n286), .ZN(n6957) );
  OR2_X1 U5684 ( .A1(n5499), .A2(n287), .ZN(n6958) );
  NAND3_X1 U5685 ( .A1(n6957), .A2(n6958), .A3(n904), .ZN(n178) );
  NAND2_X4 U5686 ( .A1(n6397), .A2(n905), .ZN(n6959) );
  NAND2_X1 U5687 ( .A1(n291), .A2(n906), .ZN(n6960) );
  NAND2_X1 U5688 ( .A1(\UUT/Mpath/the_mult/x_mult_out[26] ), .A2(n6357), .ZN(
        n6961) );
  AND3_X1 U5689 ( .A1(n6959), .A2(n6960), .A3(n6961), .ZN(n904) );
  INV_X1 U5690 ( .A(n178), .ZN(n168) );
  INV_X8 U5691 ( .A(n6962), .ZN(n6963) );
  OAI221_X1 U5692 ( .B1(n531), .B2(n296), .C1(n297), .C2(n2669), .A(n533), 
        .ZN(n3302) );
  NAND3_X4 U5693 ( .A1(\UUT/rs1_addr [0]), .A2(n7370), .A3(n6258), .ZN(n5433)
         );
  INV_X8 U5694 ( .A(n6964), .ZN(n6965) );
  INV_X2 U5695 ( .A(n878), .ZN(n948) );
  CLKBUF_X1 U5696 ( .A(\UUT/break_code[0] ), .Z(n6966) );
  AND2_X1 U5697 ( .A1(n2765), .A2(n6967), .ZN(n7015) );
  NOR2_X1 U5698 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1965 ), .A2(n7216), 
        .ZN(n6967) );
  OR2_X1 U5699 ( .A1(n7192), .A2(n7201), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1923 ) );
  CLKBUF_X1 U5700 ( .A(n6002), .Z(n6968) );
  OR2_X1 U5701 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1924 ), .A2(n6969), 
        .ZN(n7082) );
  OR2_X1 U5702 ( .A1(n6983), .A2(\UUT/Mcontrol/d_instr [26]), .ZN(n6969) );
  INV_X1 U5703 ( .A(n7101), .ZN(n1103) );
  INV_X8 U5704 ( .A(n6972), .ZN(n6973) );
  NOR2_X1 U5705 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N2015 ), 
        .ZN(n6974) );
  NOR2_X1 U5706 ( .A1(n7003), .A2(n7044), .ZN(n6975) );
  NAND2_X1 U5707 ( .A1(n1006), .A2(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
        .ZN(n1124) );
  BUF_X1 U5708 ( .A(n2763), .Z(n6976) );
  OR2_X1 U5709 ( .A1(\UUT/Mcontrol/d_sampled_finstr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2056 ), .ZN(n6977) );
  OR2_X1 U5710 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2056 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2057 ) );
  NOR2_X1 U5711 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1924 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .ZN(n6978) );
  NAND2_X1 U5712 ( .A1(n6978), .A2(n6979), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1927 ) );
  AND2_X1 U5713 ( .A1(n6980), .A2(n2765), .ZN(n6979) );
  INV_X1 U5714 ( .A(n7154), .ZN(n6980) );
  NAND2_X1 U5715 ( .A1(n6981), .A2(n7002), .ZN(n7026) );
  NOR2_X1 U5716 ( .A1(n6887), .A2(\UUT/Mcontrol/d_instr [31]), .ZN(n6981) );
  INV_X1 U5717 ( .A(n6968), .ZN(n6982) );
  OR2_X2 U5718 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1924 ), .A2(n6983), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1932 ) );
  NAND2_X1 U5719 ( .A1(n7044), .A2(n2765), .ZN(n6983) );
  NAND2_X1 U5720 ( .A1(n2765), .A2(n7044), .ZN(n7027) );
  OR2_X1 U5721 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1924 ), .A2(n6984), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1945 ) );
  NAND2_X1 U5722 ( .A1(n6985), .A2(n6976), .ZN(n6984) );
  AND2_X1 U5723 ( .A1(n2765), .A2(\UUT/Mcontrol/Operation_decoding32/N1921 ), 
        .ZN(n6985) );
  INV_X1 U5724 ( .A(n7264), .ZN(n6986) );
  NOR2_X1 U5725 ( .A1(n7035), .A2(n6986), .ZN(n6987) );
  CLKBUF_X1 U5726 ( .A(n1097), .Z(n6988) );
  OR2_X4 U5727 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1979 ), .A2(n6989), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1981 ) );
  NAND2_X1 U5728 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(n7171), 
        .ZN(n6989) );
  INV_X1 U5729 ( .A(n7040), .ZN(n6990) );
  NOR2_X4 U5730 ( .A1(n6991), .A2(n6977), .ZN(n7169) );
  NAND2_X1 U5731 ( .A1(n7171), .A2(n6990), .ZN(n6991) );
  INV_X4 U5732 ( .A(\UUT/branch_rega [7]), .ZN(n7306) );
  INV_X4 U5733 ( .A(\UUT/branch_rega [7]), .ZN(n7312) );
  INV_X4 U5734 ( .A(n7378), .ZN(n7379) );
  NOR2_X1 U5735 ( .A1(n6992), .A2(n7033), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2007 ) );
  NAND2_X1 U5736 ( .A1(n6874), .A2(n6976), .ZN(n6992) );
  OR2_X2 U5737 ( .A1(n7002), .A2(\UUT/Mcontrol/Operation_decoding32/N1923 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1924 ) );
  NAND2_X1 U5738 ( .A1(n6997), .A2(n6993), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1987 ) );
  NOR2_X1 U5739 ( .A1(n7044), .A2(\UUT/Mcontrol/Operation_decoding32/N1985 ), 
        .ZN(n6993) );
  CLKBUF_X1 U5740 ( .A(n6943), .Z(n6994) );
  NAND2_X1 U5741 ( .A1(n6939), .A2(n6869), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2005 ) );
  BUF_X2 U5742 ( .A(n2763), .Z(n6997) );
  NAND2_X1 U5743 ( .A1(n7002), .A2(n6998), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1955 ) );
  NOR2_X1 U5744 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1923 ), .A2(n6939), 
        .ZN(n6998) );
  CLKBUF_X1 U5745 ( .A(\UUT/Mcontrol/d_sampled_finstr [29]), .Z(n7002) );
  NAND2_X1 U5746 ( .A1(n7000), .A2(n7343), .ZN(n6999) );
  NOR2_X1 U5747 ( .A1(\UUT/branch_rega [22]), .A2(n7266), .ZN(n7000) );
  INV_X1 U5748 ( .A(n7158), .ZN(n7001) );
  OR2_X2 U5749 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2027 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1989 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2016 ) );
  INV_X1 U5750 ( .A(n7171), .ZN(n7003) );
  CLKBUF_X1 U5751 ( .A(n7173), .Z(n7004) );
  INV_X8 U5752 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U5753 ( .A1(n6853), .A2(n6854), .ZN(n7008) );
  INV_X1 U5754 ( .A(n7021), .ZN(n7009) );
  CLKBUF_X2 U5755 ( .A(n7022), .Z(n7021) );
  BUF_X1 U5756 ( .A(n7022), .Z(n7020) );
  NAND2_X1 U5757 ( .A1(n7011), .A2(n7159), .ZN(n7010) );
  AND2_X2 U5758 ( .A1(n7092), .A2(n7039), .ZN(n7011) );
  NAND2_X1 U5759 ( .A1(n7201), .A2(n6850), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2050 ) );
  CLKBUF_X1 U5760 ( .A(\UUT/Mcontrol/Operation_decoding32/N2007 ), .Z(n7012)
         );
  NAND2_X4 U5761 ( .A1(n7154), .A2(n7014), .ZN(n7013) );
  INV_X4 U5762 ( .A(n7013), .ZN(\UUT/Mcontrol/Operation_decoding32/N2079 ) );
  AND2_X1 U5763 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(n6997), 
        .ZN(n7016) );
  OR2_X1 U5764 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1922 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1950 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1951 ) );
  OR2_X1 U5765 ( .A1(n5467), .A2(n286), .ZN(n7017) );
  OR2_X1 U5766 ( .A1(n5465), .A2(n287), .ZN(n7018) );
  NAND3_X2 U5767 ( .A1(n7017), .A2(n7018), .A3(n942), .ZN(n939) );
  AND2_X2 U5768 ( .A1(n1438), .A2(n1439), .ZN(n5465) );
  AND3_X2 U5769 ( .A1(n7290), .A2(n7289), .A3(n7288), .ZN(n942) );
  CLKBUF_X1 U5770 ( .A(n7022), .Z(n7019) );
  NAND2_X1 U5771 ( .A1(n7154), .A2(n7070), .ZN(n7022) );
  INV_X2 U5772 ( .A(\UUT/Mcontrol/d_instr [26]), .ZN(n7154) );
  NAND2_X1 U5773 ( .A1(n7157), .A2(n7156), .ZN(n7023) );
  NOR2_X1 U5774 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1918 ), .A2(n6883), 
        .ZN(n7024) );
  NOR2_X1 U5775 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1956 ), .ZN(n7025) );
  OR2_X2 U5776 ( .A1(n7026), .A2(n7027), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1999 ) );
  AND2_X1 U5777 ( .A1(\UUT/Mpath/out_regA[0] ), .A2(n7408), .ZN(
        \UUT/Mpath/the_alu/N125 ) );
  OR2_X1 U5778 ( .A1(\UUT/Mpath/out_regA[0] ), .A2(n7408), .ZN(
        \UUT/Mpath/the_alu/N157 ) );
  NOR2_X1 U5779 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1989 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2027 ), .ZN(n7028) );
  NOR2_X1 U5780 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(n6997), 
        .ZN(n7029) );
  NAND2_X1 U5781 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(n6997), 
        .ZN(n7030) );
  INV_X8 U5782 ( .A(n7031), .ZN(n7032) );
  OR2_X2 U5783 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2002 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2027 ) );
  INV_X1 U5784 ( .A(\UUT/branch_rega [10]), .ZN(n7034) );
  NAND2_X1 U5785 ( .A1(n7072), .A2(n7034), .ZN(n7035) );
  NAND2_X1 U5786 ( .A1(n7067), .A2(n7103), .ZN(n7036) );
  OR2_X2 U5787 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2002 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2015 ) );
  INV_X4 U5788 ( .A(n7370), .ZN(\UUT/rs1_addr [1]) );
  NAND3_X2 U5789 ( .A1(n6270), .A2(n6273), .A3(\UUT/rs1_addr [1]), .ZN(n5448)
         );
  AND3_X4 U5790 ( .A1(\UUT/rs1_addr [3]), .A2(\UUT/rs1_addr [4]), .A3(n6265), 
        .ZN(n5452) );
  INV_X1 U5791 ( .A(n7100), .ZN(n7037) );
  INV_X1 U5792 ( .A(n7059), .ZN(n7100) );
  INV_X4 U5793 ( .A(\UUT/branch_rega [13]), .ZN(n7344) );
  INV_X4 U5794 ( .A(\UUT/branch_rega [13]), .ZN(n7320) );
  NAND2_X1 U5795 ( .A1(\UUT/Mcontrol/d_instr [28]), .A2(n7038), .ZN(n7043) );
  AND2_X1 U5796 ( .A1(\UUT/Mcontrol/d_instr [27]), .A2(n2763), .ZN(n7038) );
  INV_X1 U5797 ( .A(\UUT/Mcontrol/d_instr [28]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1989 ) );
  INV_X1 U5798 ( .A(n7244), .ZN(n7039) );
  NAND2_X1 U5799 ( .A1(\UUT/Mcontrol/d_instr [28]), .A2(n2764), .ZN(n7040) );
  INV_X1 U5800 ( .A(n1094), .ZN(n7041) );
  NAND2_X1 U5801 ( .A1(\UUT/Mcontrol/d_instr [29]), .A2(n7042), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1962 ) );
  NOR2_X1 U5802 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1965 ), .A2(n7133), 
        .ZN(n7042) );
  NAND2_X1 U5803 ( .A1(n6970), .A2(n7044), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2023 ) );
  INV_X4 U5804 ( .A(\UUT/Mcontrol/d_instr [27]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1921 ) );
  NOR2_X1 U5805 ( .A1(\UUT/branch_rega [26]), .A2(\UUT/branch_rega [27]), .ZN(
        n7045) );
  CLKBUF_X1 U5806 ( .A(n7036), .Z(n7046) );
  INV_X8 U5807 ( .A(n7047), .ZN(n7048) );
  AND2_X2 U5808 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1884 ), .A2(
        \UUT/Mcontrol/d_instr [2]), .ZN(n7142) );
  CLKBUF_X1 U5809 ( .A(n6870), .Z(n7049) );
  OR2_X1 U5810 ( .A1(n7270), .A2(\UUT/branch_rega [24]), .ZN(n7050) );
  INV_X8 U5811 ( .A(n7052), .ZN(n7053) );
  NAND2_X4 U5812 ( .A1(n6397), .A2(n290), .ZN(n7054) );
  NAND2_X1 U5813 ( .A1(n291), .A2(n292), .ZN(n7055) );
  NAND2_X1 U5814 ( .A1(\UUT/Mpath/the_mult/x_mult_out[24] ), .A2(n6357), .ZN(
        n7056) );
  AND3_X1 U5815 ( .A1(n7054), .A2(n7055), .A3(n7056), .ZN(n288) );
  OAI221_X1 U5816 ( .B1(n5516), .B2(n286), .C1(n5515), .C2(n287), .A(n288), 
        .ZN(n217) );
  NOR3_X2 U5817 ( .A1(\UUT/Mpath/the_alu/N486 ), .A2(n6324), .A3(
        \UUT/Mpath/the_alu/N480 ), .ZN(n2228) );
  INV_X1 U5818 ( .A(n5474), .ZN(n5364) );
  AND4_X2 U5819 ( .A1(n2182), .A2(n2183), .A3(n2184), .A4(n2185), .ZN(n5318)
         );
  INV_X8 U5820 ( .A(n7057), .ZN(n7058) );
  AND2_X2 U5821 ( .A1(n7355), .A2(n7354), .ZN(n7364) );
  AND4_X2 U5822 ( .A1(n2266), .A2(n2268), .A3(n2267), .A4(n2269), .ZN(n866) );
  INV_X2 U5823 ( .A(n217), .ZN(n207) );
  INV_X1 U5824 ( .A(n5468), .ZN(n7362) );
  OR2_X4 U5825 ( .A1(\UUT/Mpath/N115 ), .A2(\UUT/Mpath/N119 ), .ZN(n5468) );
  NAND2_X1 U5826 ( .A1(n6908), .A2(n7022), .ZN(n7060) );
  NAND2_X1 U5827 ( .A1(n7013), .A2(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
        .ZN(n7062) );
  NAND2_X1 U5828 ( .A1(n7013), .A2(n6891), .ZN(n7061) );
  NAND2_X1 U5829 ( .A1(n7013), .A2(n6891), .ZN(n2265) );
  INV_X1 U5830 ( .A(\UUT/Mcontrol/st_logic/branchlw_stall ), .ZN(
        \UUT/Mcontrol/st_logic/N13 ) );
  INV_X1 U5831 ( .A(n6920), .ZN(\UUT/Mcontrol/st_logic/N25 ) );
  NAND2_X1 U5832 ( .A1(n7173), .A2(n7063), .ZN(n1006) );
  NOR2_X1 U5833 ( .A1(n2764), .A2(n6997), .ZN(n7063) );
  NAND2_X1 U5834 ( .A1(n7064), .A2(n7044), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1950 ) );
  NAND2_X2 U5835 ( .A1(\UUT/Mpath/N115 ), .A2(n5466), .ZN(n5525) );
  INV_X4 U5836 ( .A(\UUT/Mpath/N119 ), .ZN(n5466) );
  NAND2_X1 U5837 ( .A1(n6907), .A2(n7022), .ZN(n7069) );
  NAND2_X1 U5838 ( .A1(n6050), .A2(n7022), .ZN(n7078) );
  INV_X8 U5839 ( .A(n7065), .ZN(n7066) );
  OR2_X2 U5840 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2057 ), .A2(n7043), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N2054 ) );
  OR2_X2 U5841 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1950 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1922 ), .ZN(n7067) );
  CLKBUF_X1 U5842 ( .A(n7061), .Z(n7068) );
  CLKBUF_X1 U5843 ( .A(n7067), .Z(n7071) );
  NOR2_X2 U5844 ( .A1(n6263), .A2(\UUT/rs1_addr [1]), .ZN(n6266) );
  AND3_X4 U5845 ( .A1(n6265), .A2(n2606), .A3(n6267), .ZN(n2108) );
  AND2_X1 U5846 ( .A1(n7357), .A2(n7347), .ZN(n7072) );
  OR2_X2 U5847 ( .A1(n7073), .A2(n7074), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1957 ) );
  OR2_X1 U5848 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1921 ), .ZN(n7074) );
  CLKBUF_X1 U5849 ( .A(\UUT/Mcontrol/Operation_decoding32/N1995 ), .Z(n7075)
         );
  OR2_X1 U5850 ( .A1(n7179), .A2(n6071), .ZN(n7076) );
  BUF_X1 U5851 ( .A(\UUT/branch_rega [28]), .Z(n7077) );
  OAI222_X4 U5852 ( .A1(n5382), .A2(n99), .B1(n5383), .B2(n5334), .C1(n5384), 
        .C2(n5336), .ZN(\UUT/branch_regb [23]) );
  INV_X8 U5853 ( .A(n7079), .ZN(n7080) );
  CLKBUF_X1 U5854 ( .A(\UUT/Mcontrol/Operation_decoding32/N2054 ), .Z(n7081)
         );
  CLKBUF_X1 U5855 ( .A(n6907), .Z(n7083) );
  OR2_X1 U5856 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1956 ), .ZN(n7103) );
  OR2_X1 U5857 ( .A1(n113), .A2(n99), .ZN(n7084) );
  OR2_X2 U5858 ( .A1(n114), .A2(n101), .ZN(n7085) );
  OR2_X1 U5859 ( .A1(n5365), .A2(n102), .ZN(n7086) );
  NAND3_X1 U5860 ( .A1(n7084), .A2(n7085), .A3(n7086), .ZN(n111) );
  NAND2_X4 U5861 ( .A1(n6397), .A2(n917), .ZN(n7087) );
  NAND2_X1 U5862 ( .A1(n291), .A2(n918), .ZN(n7088) );
  NAND2_X1 U5863 ( .A1(\UUT/Mpath/the_mult/x_mult_out[29] ), .A2(n6357), .ZN(
        n7089) );
  AND3_X1 U5864 ( .A1(n7087), .A2(n7088), .A3(n7089), .ZN(n916) );
  INV_X2 U5865 ( .A(n130), .ZN(n113) );
  AND4_X2 U5866 ( .A1(n1873), .A2(n1874), .A3(n1875), .A4(n1876), .ZN(n5365)
         );
  INV_X1 U5867 ( .A(\UUT/Mpath/the_mult/x_operand2 [15]), .ZN(n7090) );
  INV_X1 U5868 ( .A(\UUT/Mcontrol/Operation_decoding32/N1945 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1946 ) );
  AND2_X1 U5869 ( .A1(n7368), .A2(n7351), .ZN(n7092) );
  CLKBUF_X1 U5870 ( .A(\UUT/Mcontrol/Operation_decoding32/N2001 ), .Z(n7093)
         );
  NOR2_X1 U5871 ( .A1(n7154), .A2(\UUT/Mcontrol/Operation_decoding32/N1999 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N2001 ) );
  INV_X1 U5872 ( .A(\UUT/Mcontrol/Operation_decoding32/N1927 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1928 ) );
  NAND2_X4 U5873 ( .A1(n1048), .A2(n1051), .ZN(n6071) );
  INV_X1 U5874 ( .A(\UUT/Mpath/the_alu/N44 ), .ZN(n7094) );
  NOR2_X1 U5875 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2023 ), .ZN(n7096) );
  NOR2_X1 U5876 ( .A1(\UUT/Mcontrol/d_instr [26]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2023 ), .ZN(n7095) );
  INV_X1 U5877 ( .A(n1056), .ZN(n7097) );
  INV_X1 U5878 ( .A(n7097), .ZN(n7098) );
  INV_X1 U5879 ( .A(\UUT/Mpath/the_alu/N72 ), .ZN(n7099) );
  NAND3_X1 U5880 ( .A1(n2764), .A2(n7102), .A3(\UUT/Mcontrol/d_instr [26]), 
        .ZN(n7101) );
  NOR2_X1 U5881 ( .A1(n7033), .A2(\UUT/Mcontrol/Operation_decoding32/N2009 ), 
        .ZN(n7102) );
  NAND2_X1 U5882 ( .A1(n7082), .A2(n7118), .ZN(n7252) );
  CLKBUF_X1 U5883 ( .A(n7037), .Z(n7105) );
  INV_X4 U5884 ( .A(\UUT/Mpath/the_alu/N71 ), .ZN(n7106) );
  OR2_X2 U5885 ( .A1(n7300), .A2(\UUT/branch_rega [26]), .ZN(n7299) );
  INV_X2 U5886 ( .A(n5498), .ZN(n5373) );
  INV_X1 U5887 ( .A(\UUT/Mpath/the_alu/N62 ), .ZN(n7107) );
  INV_X1 U5888 ( .A(n1038), .ZN(n7108) );
  NOR2_X4 U5889 ( .A1(n1058), .A2(n6071), .ZN(n1039) );
  NOR2_X2 U5890 ( .A1(n2265), .A2(n6873), .ZN(n1048) );
  AND2_X2 U5891 ( .A1(n7144), .A2(n2765), .ZN(n7109) );
  NAND2_X1 U5892 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1945 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1927 ), .ZN(n7110) );
  NAND2_X1 U5893 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1945 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1927 ), .ZN(n5927) );
  OR2_X1 U5894 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1921 ), .A2(
        \UUT/Mcontrol/d_instr [26]), .ZN(n7111) );
  INV_X4 U5895 ( .A(\UUT/Mpath/the_alu/N53 ), .ZN(n7112) );
  INV_X4 U5896 ( .A(\UUT/Mpath/the_alu/N55 ), .ZN(n7113) );
  INV_X1 U5897 ( .A(\UUT/Mpath/the_alu/N74 ), .ZN(n7114) );
  INV_X2 U5898 ( .A(n5482), .ZN(n5367) );
  NAND2_X1 U5899 ( .A1(\UUT/Mpath/the_alu/diff[29] ), .A2(n1223), .ZN(n7115)
         );
  NAND2_X1 U5900 ( .A1(\UUT/Mpath/the_alu/sum[29] ), .A2(n7213), .ZN(n7116) );
  AND2_X2 U5901 ( .A1(n7115), .A2(n7116), .ZN(n1424) );
  NAND2_X2 U5902 ( .A1(\UUT/Mcontrol/d_sampled_finstr [21]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1871 ), .ZN(n7375) );
  INV_X2 U5903 ( .A(n7375), .ZN(\UUT/rs1_addr [0]) );
  NOR2_X2 U5904 ( .A1(n7375), .A2(\UUT/rs1_addr [4]), .ZN(n6278) );
  AND2_X2 U5905 ( .A1(n6271), .A2(n7370), .ZN(n6269) );
  INV_X1 U5906 ( .A(n5916), .ZN(n7117) );
  OAI222_X4 U5907 ( .A1(n5904), .A2(n6956), .B1(n7168), .B2(n5769), .C1(n7021), 
        .C2(n5906), .ZN(n6233) );
  NOR4_X4 U5908 ( .A1(n2235), .A2(n7212), .A3(n2238), .A4(
        \UUT/Mpath/the_alu/N498 ), .ZN(n6323) );
  NAND2_X2 U5909 ( .A1(\UUT/Mpath/the_alu/N515 ), .A2(\UUT/Mpath/the_alu/N509 ), .ZN(n2235) );
  AND2_X1 U5910 ( .A1(n6397), .A2(n1205), .ZN(n7119) );
  AND2_X1 U5911 ( .A1(n291), .A2(n1206), .ZN(n7120) );
  INV_X1 U5912 ( .A(\UUT/Mpath/the_alu/N58 ), .ZN(n7122) );
  NOR2_X1 U5913 ( .A1(n5927), .A2(n7252), .ZN(n7123) );
  INV_X4 U5914 ( .A(\UUT/Mpath/the_alu/N57 ), .ZN(n1245) );
  AND3_X1 U5915 ( .A1(n7071), .A2(n7103), .A3(n6890), .ZN(n7124) );
  INV_X1 U5916 ( .A(n7071), .ZN(\UUT/Mcontrol/Operation_decoding32/N1952 ) );
  INV_X1 U5917 ( .A(\UUT/Mpath/the_alu/N54 ), .ZN(n7125) );
  NAND2_X1 U5918 ( .A1(n2765), .A2(n7126), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2071 ) );
  NOR2_X1 U5919 ( .A1(n6851), .A2(\UUT/Mcontrol/Operation_decoding32/N1921 ), 
        .ZN(n7126) );
  CLKBUF_X1 U5920 ( .A(\UUT/Mcontrol/Operation_decoding32/N2066 ), .Z(n7127)
         );
  INV_X1 U5921 ( .A(\UUT/Mpath/the_alu/N66 ), .ZN(n7128) );
  INV_X4 U5922 ( .A(\UUT/Mpath/the_alu/N51 ), .ZN(n7129) );
  AND4_X2 U5923 ( .A1(n5913), .A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
        .A3(\UUT/Mcontrol/Operation_decoding32/N1987 ), .A4(n7101), .ZN(n6032)
         );
  CLKBUF_X1 U5924 ( .A(\UUT/Mcontrol/Operation_decoding32/N2071 ), .Z(n7130)
         );
  CLKBUF_X1 U5925 ( .A(n5915), .Z(n7131) );
  NOR2_X1 U5926 ( .A1(n7104), .A2(n7110), .ZN(n5915) );
  AND2_X2 U5927 ( .A1(n1369), .A2(n1368), .ZN(n5969) );
  NOR2_X4 U5928 ( .A1(n1442), .A2(\UUT/Mpath/the_shift/N118 ), .ZN(n1229) );
  INV_X4 U5929 ( .A(\UUT/Mpath/the_alu/N65 ), .ZN(n7132) );
  INV_X2 U5930 ( .A(n7195), .ZN(n7196) );
  NAND2_X1 U5931 ( .A1(n2765), .A2(n2764), .ZN(n7133) );
  INV_X1 U5932 ( .A(\UUT/Mpath/the_alu/N60 ), .ZN(n7134) );
  INV_X4 U5933 ( .A(\UUT/Mpath/the_alu/N73 ), .ZN(n1321) );
  INV_X1 U5934 ( .A(\UUT/Mpath/the_alu/N48 ), .ZN(n7135) );
  INV_X1 U5935 ( .A(\UUT/Mpath/the_alu/N52 ), .ZN(n7136) );
  INV_X1 U5936 ( .A(\UUT/Mpath/the_alu/N64 ), .ZN(n7137) );
  INV_X4 U5937 ( .A(\UUT/Mpath/the_alu/N43 ), .ZN(n7138) );
  INV_X1 U5938 ( .A(\UUT/Mpath/the_alu/N56 ), .ZN(n7140) );
  INV_X2 U5939 ( .A(\UUT/Mpath/the_alu/N59 ), .ZN(n7141) );
  INV_X2 U5940 ( .A(\UUT/Mpath/the_alu/N47 ), .ZN(n1265) );
  NAND2_X1 U5941 ( .A1(n7142), .A2(n7143), .ZN(n7209) );
  AND2_X2 U5942 ( .A1(\UUT/Mcontrol/d_instr [0]), .A2(
        \UUT/Mcontrol/d_instr [1]), .ZN(n7143) );
  NOR2_X4 U5943 ( .A1(n947), .A2(n7095), .ZN(n5920) );
  OR2_X1 U5944 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N73 ) );
  NAND2_X1 U5945 ( .A1(n7109), .A2(n7330), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1882 ) );
  AND2_X1 U5946 ( .A1(n2763), .A2(n2764), .ZN(n7144) );
  NOR3_X1 U5947 ( .A1(n7093), .A2(n7012), .A3(n7075), .ZN(n7145) );
  NAND2_X1 U5948 ( .A1(\UUT/jar_in [20]), .A2(n6867), .ZN(n7146) );
  NAND2_X1 U5949 ( .A1(n300), .A2(\UUT/branch_rega [20]), .ZN(n7147) );
  NAND2_X1 U5950 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [20]), .A2(n301), 
        .ZN(n7148) );
  AND3_X2 U5951 ( .A1(n7146), .A2(n7147), .A3(n7148), .ZN(n350) );
  OR2_X2 U5952 ( .A1(n7237), .A2(\UUT/Mcontrol/d_sampled_finstr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2002 ) );
  OAI222_X2 U5953 ( .A1(n5393), .A2(n5432), .B1(n5431), .B2(n360), .C1(n5391), 
        .C2(n5430), .ZN(\UUT/branch_rega [20]) );
  INV_X1 U5954 ( .A(n7104), .ZN(n5916) );
  BUF_X2 U5955 ( .A(n7228), .Z(n7201) );
  CLKBUF_X1 U5956 ( .A(n5948), .Z(n7151) );
  NAND3_X1 U5957 ( .A1(n7049), .A2(n7037), .A3(n6871), .ZN(n7153) );
  NAND3_X1 U5958 ( .A1(n7059), .A2(n6870), .A3(n6871), .ZN(n7152) );
  CLKBUF_X1 U5959 ( .A(\UUT/Mpath/the_mult/x_mult_out[31] ), .Z(n7155) );
  NOR2_X1 U5960 ( .A1(\UUT/branch_rega [25]), .A2(n7050), .ZN(n7157) );
  NOR2_X1 U5961 ( .A1(n7273), .A2(n7220), .ZN(n7158) );
  AND2_X2 U5962 ( .A1(n7363), .A2(n7364), .ZN(n7372) );
  NOR2_X1 U5963 ( .A1(n7160), .A2(n7182), .ZN(n7159) );
  NAND2_X1 U5964 ( .A1(n7345), .A2(n7352), .ZN(n7160) );
  NAND2_X2 U5965 ( .A1(n7162), .A2(n7224), .ZN(n7161) );
  NOR2_X1 U5966 ( .A1(\UUT/branch_rega [5]), .A2(n7265), .ZN(n7162) );
  NAND3_X1 U5967 ( .A1(n7059), .A2(n6871), .A3(n6870), .ZN(n7163) );
  INV_X1 U5968 ( .A(n7205), .ZN(n7164) );
  INV_X2 U5969 ( .A(\UUT/Mpath/the_alu/N49 ), .ZN(n1261) );
  NAND2_X1 U5970 ( .A1(n6212), .A2(n2425), .ZN(n7338) );
  INV_X1 U5971 ( .A(n7201), .ZN(\UUT/Mcontrol/d_instr [31]) );
  CLKBUF_X1 U5972 ( .A(n7077), .Z(n7166) );
  INV_X4 U5973 ( .A(\UUT/Mpath/the_alu/N45 ), .ZN(n7167) );
  CLKBUF_X1 U5974 ( .A(n7060), .Z(n7168) );
  INV_X1 U5975 ( .A(n7103), .ZN(\UUT/Mcontrol/Operation_decoding32/N1958 ) );
  OAI222_X1 U5976 ( .A1(n5899), .A2(n7225), .B1(n7168), .B2(n5905), .C1(n7021), 
        .C2(n5902), .ZN(n6085) );
  OAI222_X1 U5977 ( .A1(n5901), .A2(n7225), .B1(n7168), .B2(n5906), .C1(n7021), 
        .C2(n5903), .ZN(n6095) );
  OAI222_X4 U5978 ( .A1(n6017), .A2(n5903), .B1(n7203), .B2(n7060), .C1(n5971), 
        .C2(n7021), .ZN(n6162) );
  OAI222_X4 U5979 ( .A1(n6017), .A2(n5905), .B1(n7221), .B2(n7168), .C1(n7021), 
        .C2(n6035), .ZN(n6171) );
  NAND3_X4 U5980 ( .A1(n6263), .A2(n6275), .A3(n6276), .ZN(n5453) );
  NAND2_X1 U5981 ( .A1(n7170), .A2(n7171), .ZN(n7172) );
  INV_X1 U5982 ( .A(\UUT/Mcontrol/Operation_decoding32/N2071 ), .ZN(n7170) );
  INV_X1 U5983 ( .A(n6976), .ZN(n7171) );
  INV_X1 U5984 ( .A(n7327), .ZN(n805) );
  NAND2_X1 U5985 ( .A1(n7044), .A2(n7004), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2047 ) );
  NOR2_X1 U5986 ( .A1(n6851), .A2(\UUT/Mcontrol/Operation_decoding32/N1989 ), 
        .ZN(n7173) );
  NAND2_X1 U5987 ( .A1(n7231), .A2(n7232), .ZN(n7174) );
  INV_X1 U5988 ( .A(n7174), .ZN(n7233) );
  OR2_X1 U5989 ( .A1(n7154), .A2(\UUT/Mcontrol/Operation_decoding32/N2047 ), 
        .ZN(n7175) );
  NAND3_X4 U5990 ( .A1(\UUT/rs1_addr [1]), .A2(n6273), .A3(n6278), .ZN(n5461)
         );
  AND2_X4 U5991 ( .A1(n6278), .A2(n6275), .ZN(n6274) );
  AND2_X4 U5992 ( .A1(n6269), .A2(n6278), .ZN(n2115) );
  AND2_X4 U5993 ( .A1(n6274), .A2(n6266), .ZN(n5458) );
  OR2_X4 U5994 ( .A1(n5475), .A2(n5466), .ZN(n7176) );
  OR2_X1 U5995 ( .A1(n5476), .A2(n5468), .ZN(n7177) );
  NAND2_X1 U5996 ( .A1(n7176), .A2(n7177), .ZN(n5474) );
  INV_X1 U5997 ( .A(n1422), .ZN(n5476) );
  OR2_X1 U5998 ( .A1(n7153), .A2(n7096), .ZN(n7179) );
  INV_X1 U5999 ( .A(n7183), .ZN(n7181) );
  NAND2_X1 U6000 ( .A1(n7369), .A2(n7181), .ZN(n7182) );
  AND4_X2 U6001 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n312) );
  NAND2_X1 U6002 ( .A1(n7187), .A2(n7333), .ZN(n7183) );
  INV_X1 U6003 ( .A(n7153), .ZN(n1050) );
  AND2_X4 U6004 ( .A1(n7154), .A2(n7184), .ZN(n1058) );
  NOR2_X1 U6005 ( .A1(n7044), .A2(\UUT/Mcontrol/Operation_decoding32/N2088 ), 
        .ZN(n7184) );
  INV_X1 U6006 ( .A(n7051), .ZN(n1059) );
  OAI222_X4 U6007 ( .A1(n5373), .A2(n99), .B1(n5374), .B2(n5334), .C1(n5375), 
        .C2(n5336), .ZN(\UUT/branch_regb [26]) );
  OAI222_X1 U6008 ( .A1(n5364), .A2(n5430), .B1(n5318), .B2(n5431), .C1(n5366), 
        .C2(n5432), .ZN(\UUT/branch_rega [29]) );
  NOR2_X1 U6009 ( .A1(n7178), .A2(\UUT/Mcontrol/Nextpc_decoding/N127 ), .ZN(
        n7277) );
  NAND2_X1 U6010 ( .A1(\UUT/Mpath/the_alu/N474 ), .A2(n2228), .ZN(n1305) );
  INV_X1 U6011 ( .A(n7301), .ZN(n7187) );
  INV_X1 U6012 ( .A(\UUT/Mpath/out_regA[9] ), .ZN(n7195) );
  INV_X4 U6013 ( .A(\UUT/Mpath/the_alu/N67 ), .ZN(n7189) );
  INV_X1 U6014 ( .A(\UUT/Mpath/the_alu/N46 ), .ZN(n7190) );
  INV_X1 U6015 ( .A(n7164), .ZN(n7191) );
  INV_X2 U6016 ( .A(\UUT/Mpath/the_alu/N63 ), .ZN(n1219) );
  INV_X1 U6017 ( .A(\UUT/Mpath/the_alu/N59 ), .ZN(n7193) );
  INV_X1 U6018 ( .A(\UUT/Mpath/the_alu/N44 ), .ZN(n7194) );
  AND4_X1 U6019 ( .A1(n2523), .A2(n2524), .A3(n2525), .A4(n2526), .ZN(n686) );
  BUF_X8 U6020 ( .A(\UUT/Mpath/out_regB[2] ), .Z(n7402) );
  INV_X1 U6021 ( .A(\UUT/Mpath/the_alu/N50 ), .ZN(n7197) );
  INV_X4 U6022 ( .A(\UUT/Mpath/the_alu/N61 ), .ZN(n7198) );
  INV_X1 U6023 ( .A(n7199), .ZN(n7200) );
  INV_X1 U6024 ( .A(n7221), .ZN(n7202) );
  INV_X1 U6025 ( .A(\UUT/Mcontrol/d_sampled_finstr [5]), .ZN(n7203) );
  OAI222_X4 U6026 ( .A1(n5364), .A2(n99), .B1(n5365), .B2(n5334), .C1(n5366), 
        .C2(n5336), .ZN(\UUT/branch_regb [29]) );
  AOI221_X4 U6027 ( .B1(n5991), .B2(n2242), .C1(
        \UUT/Mcontrol/d_sampled_finstr [5]), .C2(n2243), .A(n2244), .ZN(n325)
         );
  OR2_X1 U6028 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1900 ), .A2(
        \UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1902 ) );
  CLKBUF_X1 U6029 ( .A(n6827), .Z(n7204) );
  AOI221_X4 U6030 ( .B1(n1121), .B2(n1050), .C1(n1122), .C2(n1123), .A(n7204), 
        .ZN(n1116) );
  NAND2_X1 U6031 ( .A1(\UUT/Mpath/the_alu/diff[30] ), .A2(n1223), .ZN(n7206)
         );
  NAND2_X1 U6032 ( .A1(\UUT/Mpath/the_alu/sum[30] ), .A2(n7213), .ZN(n7207) );
  AND2_X2 U6033 ( .A1(n7206), .A2(n7207), .ZN(n1433) );
  INV_X1 U6034 ( .A(n6892), .ZN(n1051) );
  OR2_X1 U6035 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N1917 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1918 ) );
  OR2_X1 U6036 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N2081 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N2088 ) );
  OR2_X1 U6037 ( .A1(\UUT/Mcontrol/Operation_decoding32/N2081 ), .A2(n6939), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N2082 ) );
  OR2_X1 U6038 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N1984 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1985 ) );
  OR2_X1 U6039 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N1978 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1979 ) );
  OR2_X1 U6040 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N1984 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1973 ) );
  INV_X1 U6041 ( .A(n7221), .ZN(\UUT/Mcontrol/d_instr [4]) );
  OR2_X1 U6042 ( .A1(\UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1903 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1904 ) );
  OR2_X1 U6043 ( .A1(\UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1909 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1910 ) );
  AND2_X1 U6044 ( .A1(\UUT/Mcontrol/d_instr [2]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1895 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1896 ) );
  OR2_X1 U6045 ( .A1(n6939), .A2(\UUT/Mcontrol/Operation_decoding32/N1890 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1891 ) );
  AOI221_X4 U6046 ( .B1(n6001), .B2(n2242), .C1(\UUT/Mcontrol/d_instr [4]), 
        .C2(n2243), .A(n2244), .ZN(n348) );
  INV_X1 U6047 ( .A(\UUT/Mcontrol/d_instr [4]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1900 ) );
  OR2_X1 U6048 ( .A1(\UUT/Mcontrol/d_instr [4]), .A2(\UUT/Mcontrol/d_instr [5]), .ZN(\UUT/Mcontrol/Operation_decoding32/N1908 ) );
  AND2_X1 U6049 ( .A1(n7202), .A2(\UUT/Mcontrol/d_instr [5]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1894 ) );
  INV_X2 U6050 ( .A(n1216), .ZN(n7211) );
  INV_X1 U6051 ( .A(n7211), .ZN(n7212) );
  INV_X8 U6052 ( .A(n7211), .ZN(n7213) );
  INV_X1 U6053 ( .A(n1295), .ZN(n7214) );
  INV_X4 U6054 ( .A(n7214), .ZN(n7215) );
  NOR2_X1 U6055 ( .A1(n1218), .A2(n6834), .ZN(n1295) );
  INV_X4 U6056 ( .A(n1305), .ZN(n1220) );
  INV_X1 U6057 ( .A(\UUT/Mcontrol/d_sampled_finstr [3]), .ZN(n5327) );
  OAI221_X1 U6058 ( .B1(n2253), .B2(n2254), .C1(n5327), .C2(n2255), .A(n2256), 
        .ZN(\UUT/break_code[19] ) );
  AND2_X1 U6059 ( .A1(\UUT/Mpath/out_regA[2] ), .A2(n7404), .ZN(
        \UUT/Mpath/the_alu/N123 ) );
  OR2_X1 U6060 ( .A1(\UUT/Mpath/out_regA[2] ), .A2(n7404), .ZN(
        \UUT/Mpath/the_alu/N155 ) );
  OR2_X1 U6061 ( .A1(\UUT/Mcontrol/d_sampled_finstr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1902 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1903 ) );
  OR2_X1 U6062 ( .A1(\UUT/Mcontrol/d_sampled_finstr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1908 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1909 ) );
  AND2_X1 U6063 ( .A1(\UUT/Mcontrol/d_sampled_finstr [3]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1894 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1895 ) );
  INV_X4 U6064 ( .A(\UUT/branch_rega [10]), .ZN(n7342) );
  INV_X1 U6065 ( .A(\UUT/Mcontrol/d_instr [29]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1877 ) );
  AND2_X2 U6066 ( .A1(n1366), .A2(n1367), .ZN(n5980) );
  OR2_X1 U6067 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1877 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1916 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1917 ) );
  OR2_X1 U6068 ( .A1(\UUT/Mcontrol/d_instr [29]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N2008 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2009 ) );
  OR2_X1 U6069 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1889 ), .A2(n7216), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1890 ) );
  AND2_X2 U6070 ( .A1(n1292), .A2(n1293), .ZN(n6111) );
  AND4_X2 U6071 ( .A1(n2130), .A2(n2131), .A3(n2132), .A4(n2133), .ZN(n5322)
         );
  INV_X2 U6072 ( .A(n5506), .ZN(n5376) );
  NOR2_X4 U6073 ( .A1(n5877), .A2(\UUT/rs2_addr [4]), .ZN(n5895) );
  INV_X2 U6074 ( .A(\UUT/rs2_addr [0]), .ZN(n5877) );
  OAI222_X4 U6075 ( .A1(n5402), .A2(n5432), .B1(n5431), .B2(n411), .C1(n5400), 
        .C2(n5430), .ZN(\UUT/branch_rega [18]) );
  AND2_X4 U6076 ( .A1(n6269), .A2(n6270), .ZN(n5446) );
  INV_X32 U6077 ( .A(\UUT/Mcontrol/Nextpc_decoding/N159 ), .ZN(n7218) );
  INV_X4 U6078 ( .A(\UUT/Mpath/the_shift/N117 ), .ZN(
        \UUT/Mpath/the_shift/N118 ) );
  AND2_X2 U6079 ( .A1(n6282), .A2(\UUT/Mpath/the_shift/N107 ), .ZN(n1228) );
  AOI222_X1 U6080 ( .A1(\UUT/Mpath/the_shift/sh_rol [31]), .A2(n1226), .B1(
        \UUT/Mpath/the_shift/sh_ror [31]), .B2(n6342), .C1(
        \UUT/Mpath/the_shift/sh_sll [31]), .C2(n1228), .ZN(n1293) );
  NOR2_X4 U6081 ( .A1(n1441), .A2(\UUT/Mpath/the_shift/N107 ), .ZN(n1226) );
  INV_X2 U6082 ( .A(n7217), .ZN(\UUT/Mcontrol/d_instr [5]) );
  INV_X1 U6083 ( .A(n7304), .ZN(n7220) );
  OR2_X1 U6084 ( .A1(\UUT/branch_rega [11]), .A2(n7250), .ZN(n7223) );
  OR2_X2 U6085 ( .A1(\UUT/branch_rega [30]), .A2(\UUT/branch_rega [31]), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N127 ) );
  NAND3_X4 U6086 ( .A1(n2229), .A2(n2230), .A3(\UUT/Mpath/the_alu/N480 ), .ZN(
        n1301) );
  INV_X4 U6087 ( .A(n1301), .ZN(n1221) );
  NOR2_X1 U6088 ( .A1(\UUT/branch_rega [2]), .A2(n7239), .ZN(n7224) );
  CLKBUF_X1 U6089 ( .A(n6956), .Z(n7225) );
  INV_X1 U6090 ( .A(n6855), .ZN(n7226) );
  INV_X1 U6091 ( .A(n6855), .ZN(n7227) );
  NAND2_X1 U6092 ( .A1(n6995), .A2(n6203), .ZN(n7229) );
  NAND2_X1 U6093 ( .A1(\UUT/Mcontrol/d_sampled_finstr [3]), .A2(n6134), .ZN(
        n7230) );
  AND2_X2 U6094 ( .A1(n7229), .A2(n7230), .ZN(n6202) );
  NAND2_X1 U6095 ( .A1(n6201), .A2(n2425), .ZN(n7231) );
  NAND2_X1 U6096 ( .A1(n2426), .A2(\UUT/Mcontrol/d_sampled_finstr [3]), .ZN(
        n7232) );
  INV_X1 U6097 ( .A(n5464), .ZN(n7234) );
  NOR2_X1 U6098 ( .A1(n7303), .A2(n6254), .ZN(n7235) );
  NOR2_X1 U6099 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N242 ), .A2(n6255), .ZN(
        n7236) );
  OR2_X1 U6100 ( .A1(n7235), .A2(n7236), .ZN(n6251) );
  INV_X1 U6101 ( .A(n5464), .ZN(n5358) );
  INV_X1 U6102 ( .A(\UUT/Mcontrol/Nextpc_decoding/N241 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N242 ) );
  CLKBUF_X1 U6103 ( .A(\UUT/branch_rega [30]), .Z(n7324) );
  NOR2_X2 U6104 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N25 ), .A2(n6247), .ZN(
        n6248) );
  AND2_X2 U6105 ( .A1(n7328), .A2(n7329), .ZN(n6213) );
  OR2_X1 U6106 ( .A1(n7240), .A2(\UUT/branch_rega [1]), .ZN(n7239) );
  INV_X1 U6107 ( .A(\UUT/branch_rega [0]), .ZN(n7240) );
  INV_X1 U6108 ( .A(n7259), .ZN(n7260) );
  OR2_X1 U6109 ( .A1(\UUT/branch_rega [26]), .A2(\UUT/branch_rega [25]), .ZN(
        n7259) );
  OAI222_X4 U6110 ( .A1(n5363), .A2(n5432), .B1(n5431), .B2(n816), .C1(n5361), 
        .C2(n5430), .ZN(\UUT/branch_rega [2]) );
  NAND3_X4 U6111 ( .A1(\UUT/rs2_addr [1]), .A2(n6933), .A3(n5891), .ZN(n5648)
         );
  AND2_X2 U6112 ( .A1(n5895), .A2(n5892), .ZN(n5891) );
  INV_X4 U6113 ( .A(\UUT/branch_rega [9]), .ZN(n7292) );
  OR2_X2 U6114 ( .A1(\UUT/branch_rega [9]), .A2(n7263), .ZN(n7262) );
  OR2_X1 U6115 ( .A1(n7280), .A2(n7242), .ZN(n7241) );
  INV_X1 U6116 ( .A(n7278), .ZN(n7242) );
  INV_X1 U6117 ( .A(n7241), .ZN(n7243) );
  NAND2_X2 U6118 ( .A1(n7342), .A2(n7243), .ZN(n7244) );
  NAND2_X1 U6119 ( .A1(n7305), .A2(n7248), .ZN(n7245) );
  NAND2_X1 U6120 ( .A1(n7245), .A2(n7246), .ZN(n6253) );
  OR2_X1 U6121 ( .A1(n7247), .A2(\UUT/Mcontrol/Nextpc_decoding/N159 ), .ZN(
        n7246) );
  INV_X1 U6122 ( .A(\UUT/Mcontrol/Nextpc_decoding/N248 ), .ZN(n7247) );
  AND2_X1 U6123 ( .A1(n7269), .A2(\UUT/Mcontrol/Nextpc_decoding/N248 ), .ZN(
        n7248) );
  INV_X1 U6124 ( .A(n7271), .ZN(n7249) );
  NAND2_X1 U6125 ( .A1(n7311), .A2(n7249), .ZN(n7250) );
  NOR4_X4 U6126 ( .A1(n5922), .A2(n5899), .A3(n5923), .A4(n5924), .ZN(
        \UUT/Mcontrol/st_logic/N104 ) );
  NAND3_X4 U6127 ( .A1(n5926), .A2(n7251), .A3(n6243), .ZN(
        \UUT/Mcontrol/d_jump_type[3] ) );
  NAND2_X2 U6128 ( .A1(n1039), .A2(n1050), .ZN(n947) );
  OAI221_X4 U6129 ( .B1(n2253), .B2(n2257), .C1(n7210), .C2(n2255), .A(n2256), 
        .ZN(\UUT/break_code[18] ) );
  OR2_X1 U6130 ( .A1(\UUT/Mpath/out_regA[3] ), .A2(n7401), .ZN(
        \UUT/Mpath/the_alu/N154 ) );
  AND2_X1 U6131 ( .A1(\UUT/Mpath/out_regA[3] ), .A2(n7401), .ZN(
        \UUT/Mpath/the_alu/N122 ) );
  INV_X4 U6132 ( .A(\UUT/branch_rega [23]), .ZN(n7291) );
  INV_X4 U6133 ( .A(\UUT/branch_rega [23]), .ZN(n7346) );
  NOR2_X2 U6134 ( .A1(\UUT/branch_rega [24]), .A2(\UUT/branch_rega [23]), .ZN(
        n7275) );
  INV_X1 U6135 ( .A(n5923), .ZN(n7251) );
  INV_X1 U6136 ( .A(n7124), .ZN(n5923) );
  AND2_X2 U6137 ( .A1(n7373), .A2(n7374), .ZN(n7294) );
  AND2_X2 U6138 ( .A1(n7365), .A2(n7366), .ZN(n7374) );
  INV_X4 U6139 ( .A(\UUT/branch_rega [15]), .ZN(n7371) );
  INV_X1 U6140 ( .A(\UUT/Mcontrol/Operation_decoding32/N1933 ), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1934 ) );
  INV_X1 U6141 ( .A(n7118), .ZN(\UUT/Mcontrol/Operation_decoding32/N1940 ) );
  AOI211_X4 U6142 ( .C1(n5916), .C2(n5917), .A(n7046), .B(n5934), .ZN(n6133)
         );
  INV_X4 U6143 ( .A(\UUT/branch_rega [6]), .ZN(n7331) );
  INV_X4 U6144 ( .A(n7262), .ZN(n7264) );
  INV_X4 U6145 ( .A(\UUT/branch_rega [16]), .ZN(n7363) );
  AND3_X2 U6146 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1951 ), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1957 ), .A3(n6135), .ZN(n7253) );
  INV_X1 U6147 ( .A(\UUT/branch_rega [5]), .ZN(n7349) );
  INV_X1 U6148 ( .A(\UUT/branch_rega [5]), .ZN(n7345) );
  OAI222_X4 U6149 ( .A1(n5348), .A2(n5432), .B1(n5431), .B2(n741), .C1(n5346), 
        .C2(n5430), .ZN(\UUT/branch_rega [5]) );
  NAND2_X1 U6150 ( .A1(\UUT/jar_in [21]), .A2(n6867), .ZN(n7255) );
  NAND2_X1 U6151 ( .A1(n300), .A2(\UUT/branch_rega [21]), .ZN(n7256) );
  NAND2_X1 U6152 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [21]), .A2(n301), 
        .ZN(n7257) );
  AND3_X2 U6153 ( .A1(n7255), .A2(n7256), .A3(n7257), .ZN(n327) );
  INV_X4 U6154 ( .A(\UUT/branch_rega [2]), .ZN(n7333) );
  INV_X4 U6155 ( .A(\UUT/branch_rega [2]), .ZN(n7293) );
  OR2_X1 U6156 ( .A1(n7051), .A2(n6030), .ZN(n7258) );
  NAND2_X1 U6157 ( .A1(n7258), .A2(n6031), .ZN(n5960) );
  NOR2_X2 U6158 ( .A1(\UUT/branch_rega [27]), .A2(
        \UUT/Mcontrol/Nextpc_decoding/N194 ), .ZN(n7261) );
  INV_X1 U6159 ( .A(n7296), .ZN(n7263) );
  INV_X1 U6160 ( .A(n7295), .ZN(n7265) );
  INV_X1 U6161 ( .A(\UUT/branch_rega [17]), .ZN(n7354) );
  INV_X1 U6162 ( .A(n7334), .ZN(n7267) );
  OR2_X1 U6163 ( .A1(\UUT/branch_rega [1]), .A2(\UUT/branch_rega [0]), .ZN(
        n7268) );
  INV_X32 U6164 ( .A(n7268), .ZN(n7269) );
  INV_X1 U6165 ( .A(n7291), .ZN(n7270) );
  OR2_X1 U6166 ( .A1(n7272), .A2(\UUT/branch_rega [14]), .ZN(n7271) );
  INV_X1 U6167 ( .A(n7320), .ZN(n7272) );
  OR2_X1 U6168 ( .A1(n7274), .A2(\UUT/branch_rega [10]), .ZN(n7273) );
  INV_X1 U6169 ( .A(n7292), .ZN(n7274) );
  OAI222_X4 U6170 ( .A1(n5427), .A2(n5430), .B1(n5324), .B2(n5431), .C1(n5429), 
        .C2(n5432), .ZN(\UUT/branch_rega [0]) );
  NOR2_X1 U6171 ( .A1(\UUT/branch_rega [28]), .A2(\UUT/branch_rega [27]), .ZN(
        n7276) );
  AND2_X1 U6172 ( .A1(n7279), .A2(n7306), .ZN(n7278) );
  INV_X1 U6173 ( .A(\UUT/branch_rega [6]), .ZN(n7279) );
  OR2_X1 U6174 ( .A1(n7281), .A2(\UUT/branch_rega [9]), .ZN(n7280) );
  INV_X1 U6175 ( .A(n7282), .ZN(n7281) );
  AND2_X2 U6176 ( .A1(n7293), .A2(n7294), .ZN(n7305) );
  INV_X1 U6177 ( .A(\UUT/branch_rega [18]), .ZN(n7353) );
  AND4_X2 U6178 ( .A1(n2344), .A2(n2345), .A3(n2346), .A4(n2347), .ZN(n411) );
  OAI221_X1 U6179 ( .B1(n507), .B2(n296), .C1(n297), .C2(n2666), .A(n509), 
        .ZN(n3262) );
  NAND2_X1 U6180 ( .A1(n7314), .A2(n7315), .ZN(n7283) );
  NAND2_X1 U6181 ( .A1(n298), .A2(n7284), .ZN(n2942) );
  INV_X1 U6182 ( .A(n7283), .ZN(n7284) );
  OR2_X1 U6183 ( .A1(n7313), .A2(\UUT/Mcontrol/Operation_decoding32/N1901 ), 
        .ZN(n7285) );
  NAND2_X1 U6184 ( .A1(n7285), .A2(n2264), .ZN(\UUT/break_code[0] ) );
  AND3_X2 U6185 ( .A1(n7316), .A2(n7317), .A3(n7318), .ZN(n298) );
  INV_X1 U6186 ( .A(\UUT/Mcontrol/d_instr [0]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1901 ) );
  INV_X4 U6187 ( .A(\UUT/branch_rega [19]), .ZN(n7343) );
  OAI221_X1 U6188 ( .B1(n325), .B2(n296), .C1(n297), .C2(n2645), .A(n327), 
        .ZN(n2982) );
  NAND2_X1 U6189 ( .A1(n92), .A2(n93), .ZN(n7286) );
  NAND2_X4 U6190 ( .A1(\UUT/Mpath/the_mult/x_operand2 [30]), .A2(n6340), .ZN(
        n7287) );
  AND2_X1 U6191 ( .A1(n7286), .A2(n7287), .ZN(n91) );
  NAND2_X4 U6192 ( .A1(n6397), .A2(n943), .ZN(n7288) );
  NAND2_X1 U6193 ( .A1(n291), .A2(n944), .ZN(n7289) );
  NAND2_X1 U6194 ( .A1(\UUT/Mpath/the_mult/x_mult_out[30] ), .A2(n6357), .ZN(
        n7290) );
  INV_X1 U6195 ( .A(\UUT/branch_rega [20]), .ZN(n7334) );
  AND2_X1 U6196 ( .A1(n7358), .A2(n7348), .ZN(n7295) );
  AND2_X1 U6197 ( .A1(n7297), .A2(n7379), .ZN(n7296) );
  INV_X1 U6198 ( .A(\UUT/branch_rega [6]), .ZN(n7297) );
  CLKBUF_X1 U6199 ( .A(\UUT/branch_rega [31]), .Z(n7303) );
  AND4_X2 U6200 ( .A1(n2208), .A2(n2209), .A3(n2210), .A4(n2211), .ZN(n5316)
         );
  OAI221_X1 U6201 ( .B1(n86), .B2(n81), .C1(n87), .C2(n6340), .A(n88), .ZN(
        n2869) );
  AND3_X4 U6202 ( .A1(n6275), .A2(n6267), .A3(n6265), .ZN(n5459) );
  AND2_X2 U6203 ( .A1(n6266), .A2(n7375), .ZN(n6265) );
  OAI222_X4 U6204 ( .A1(n5420), .A2(n5432), .B1(n5431), .B2(n568), .C1(n5418), 
        .C2(n5430), .ZN(\UUT/branch_rega [12]) );
  INV_X2 U6205 ( .A(n6221), .ZN(n5418) );
  INV_X1 U6206 ( .A(n7321), .ZN(n7300) );
  OR2_X1 U6207 ( .A1(\UUT/branch_rega [1]), .A2(\UUT/branch_rega [0]), .ZN(
        n7301) );
  OAI222_X1 U6208 ( .A1(n7359), .A2(n5430), .B1(n5316), .B2(n5431), .C1(n5357), 
        .C2(n5432), .ZN(\UUT/branch_rega [31]) );
  OR2_X1 U6209 ( .A1(n7302), .A2(n7303), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N27 ) );
  OAI221_X1 U6210 ( .B1(n833), .B2(n296), .C1(n297), .C2(n2703), .A(n836), 
        .ZN(n3780) );
  OAI222_X4 U6211 ( .A1(n5339), .A2(n5432), .B1(n5431), .B2(n662), .C1(n5337), 
        .C2(n5430), .ZN(\UUT/branch_rega [8]) );
  OAI222_X4 U6212 ( .A1(n5342), .A2(n5432), .B1(n5431), .B2(n686), .C1(n5340), 
        .C2(n5430), .ZN(\UUT/branch_rega [7]) );
  OAI221_X1 U6213 ( .B1(n422), .B2(n296), .C1(n297), .C2(n2657), .A(n425), 
        .ZN(n3142) );
  OAI221_X1 U6214 ( .B1(n398), .B2(n296), .C1(n297), .C2(n2654), .A(n401), 
        .ZN(n3102) );
  INV_X1 U6215 ( .A(n7322), .ZN(n7307) );
  NOR2_X1 U6216 ( .A1(\UUT/branch_rega [13]), .A2(n7307), .ZN(n7308) );
  OR2_X1 U6217 ( .A1(\UUT/branch_rega [19]), .A2(\UUT/branch_rega [20]), .ZN(
        n7309) );
  AND2_X1 U6218 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N236 ), .A2(n7303), .ZN(
        n7310) );
  NOR2_X1 U6219 ( .A1(n7310), .A2(n6256), .ZN(n6255) );
  INV_X1 U6220 ( .A(\UUT/Mcontrol/Nextpc_decoding/N235 ), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/N236 ) );
  OAI22_X1 U6221 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N27 ), .A2(n6249), .B1(
        n6250), .B2(\UUT/Mcontrol/Nextpc_decoding/N254 ), .ZN(n6246) );
  OAI221_X1 U6222 ( .B1(n371), .B2(n296), .C1(n297), .C2(n2651), .A(n374), 
        .ZN(n3062) );
  NOR2_X4 U6223 ( .A1(n2231), .A2(\UUT/Mpath/the_alu/N474 ), .ZN(n1218) );
  OAI222_X4 U6224 ( .A1(n5417), .A2(n5432), .B1(n5431), .B2(n543), .C1(n5415), 
        .C2(n5430), .ZN(\UUT/branch_rega [13]) );
  NAND3_X2 U6225 ( .A1(n6267), .A2(n7375), .A3(n6269), .ZN(n2112) );
  AND2_X1 U6226 ( .A1(\UUT/Mpath/out_regA[4] ), .A2(n7400), .ZN(
        \UUT/Mpath/the_alu/N121 ) );
  OR2_X1 U6227 ( .A1(\UUT/Mpath/out_regA[4] ), .A2(n7400), .ZN(
        \UUT/Mpath/the_alu/N153 ) );
  AOI22_X1 U6228 ( .A1(n1056), .A2(n5959), .B1(n5900), .B2(n7068), .ZN(n7313)
         );
  OR2_X1 U6229 ( .A1(n294), .A2(n296), .ZN(n7314) );
  OR2_X1 U6230 ( .A1(n297), .A2(n2642), .ZN(n7315) );
  NAND2_X1 U6231 ( .A1(\UUT/jar_in [22]), .A2(n6867), .ZN(n7316) );
  NAND2_X1 U6232 ( .A1(n300), .A2(\UUT/branch_rega [22]), .ZN(n7317) );
  NAND2_X1 U6233 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [22]), .A2(n6930), 
        .ZN(n7318) );
  AOI22_X1 U6234 ( .A1(n5959), .A2(n1056), .B1(n5900), .B2(n7068), .ZN(n2252)
         );
  INV_X1 U6235 ( .A(\UUT/branch_rega [25]), .ZN(n7321) );
  NAND2_X1 U6236 ( .A1(\UUT/Mcontrol/Nextpc_decoding/Bta [23]), .A2(n6930), 
        .ZN(n7319) );
  INV_X1 U6237 ( .A(\UUT/branch_rega [12]), .ZN(n7351) );
  AND2_X1 U6238 ( .A1(n7323), .A2(n7335), .ZN(n7322) );
  INV_X1 U6239 ( .A(\UUT/branch_rega [14]), .ZN(n7323) );
  NAND2_X1 U6240 ( .A1(n7336), .A2(n7337), .ZN(n7325) );
  NAND2_X1 U6241 ( .A1(n7319), .A2(n7149), .ZN(n4159) );
  INV_X1 U6242 ( .A(n7325), .ZN(n7326) );
  CLKBUF_X1 U6243 ( .A(n7238), .Z(n7327) );
  NAND2_X1 U6244 ( .A1(n6214), .A2(n6849), .ZN(n7328) );
  NAND2_X1 U6245 ( .A1(\UUT/Mcontrol/d_instr [2]), .A2(n6134), .ZN(n7329) );
  INV_X2 U6246 ( .A(n7210), .ZN(\UUT/Mcontrol/d_instr [2]) );
  INV_X1 U6247 ( .A(\UUT/branch_rega [15]), .ZN(n7335) );
  NOR2_X1 U6248 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1889 ), .A2(n7216), 
        .ZN(n7330) );
  OAI221_X1 U6249 ( .B1(n348), .B2(n296), .C1(n297), .C2(n2648), .A(n350), 
        .ZN(n3022) );
  OAI221_X1 U6250 ( .B1(n446), .B2(n296), .C1(n297), .C2(n2660), .A(n449), 
        .ZN(n3182) );
  BUF_X8 U6251 ( .A(\UUT/Mpath/out_regB[3] ), .Z(n7401) );
  NOR2_X2 U6252 ( .A1(n6275), .A2(\UUT/rs1_addr [2]), .ZN(n6271) );
  NAND2_X4 U6253 ( .A1(n6276), .A2(n6271), .ZN(n5462) );
  INV_X2 U6254 ( .A(\UUT/rs1_addr [2]), .ZN(n6263) );
  NAND3_X4 U6255 ( .A1(n6263), .A2(n7370), .A3(n6274), .ZN(n2113) );
  OR2_X1 U6256 ( .A1(\UUT/Mcontrol/d_jump_type[3] ), .A2(
        \UUT/Mcontrol/st_logic/N104 ), .ZN(\UUT/Mcontrol/st_logic/N79 ) );
  INV_X8 U6257 ( .A(n556), .ZN(n297) );
  NAND2_X4 U6258 ( .A1(\UUT/Mcontrol/N22 ), .A2(n1013), .ZN(n556) );
  AND2_X1 U6259 ( .A1(\UUT/Mpath/out_regA[23] ), .A2(\UUT/Mpath/out_regB[23] ), 
        .ZN(\UUT/Mpath/the_alu/N102 ) );
  OR2_X1 U6260 ( .A1(\UUT/Mpath/out_regA[23] ), .A2(\UUT/Mpath/out_regB[23] ), 
        .ZN(\UUT/Mpath/the_alu/N134 ) );
  AND2_X1 U6261 ( .A1(\UUT/Mpath/out_regA[22] ), .A2(\UUT/Mpath/out_regB[22] ), 
        .ZN(\UUT/Mpath/the_alu/N103 ) );
  OR2_X1 U6262 ( .A1(\UUT/Mpath/out_regA[22] ), .A2(\UUT/Mpath/out_regB[22] ), 
        .ZN(\UUT/Mpath/the_alu/N135 ) );
  OR2_X1 U6263 ( .A1(n84), .A2(n296), .ZN(n7336) );
  OR2_X1 U6264 ( .A1(n297), .A2(n2710), .ZN(n7337) );
  NAND2_X1 U6265 ( .A1(n2426), .A2(\UUT/Mcontrol/d_sampled_finstr [2]), .ZN(
        n7339) );
  AND2_X1 U6266 ( .A1(n300), .A2(\UUT/branch_rega [23]), .ZN(n7340) );
  AND2_X2 U6267 ( .A1(n6189), .A2(n1132), .ZN(n2425) );
  OAI222_X4 U6268 ( .A1(n5384), .A2(n5432), .B1(n5431), .B2(n866), .C1(n5382), 
        .C2(n5430), .ZN(\UUT/branch_rega [23]) );
  INV_X4 U6269 ( .A(\UUT/branch_rega [11]), .ZN(n7368) );
  INV_X4 U6270 ( .A(\UUT/branch_rega [11]), .ZN(n7357) );
  AND4_X2 U6271 ( .A1(n7123), .A2(n7024), .A3(n7253), .A4(n7008), .ZN(n7341)
         );
  OAI222_X4 U6272 ( .A1(n5358), .A2(n99), .B1(n5359), .B2(n5334), .C1(n5360), 
        .C2(n5336), .ZN(\UUT/branch_regb [30]) );
  OAI222_X1 U6273 ( .A1(n7234), .A2(n5430), .B1(n5317), .B2(n5431), .C1(n5360), 
        .C2(n5432), .ZN(\UUT/branch_rega [30]) );
  AND2_X1 U6274 ( .A1(n7167), .A2(n7190), .ZN(\UUT/Mpath/the_alu/N106 ) );
  OR2_X1 U6275 ( .A1(n7167), .A2(n7190), .ZN(\UUT/Mpath/the_alu/N138 ) );
  OAI222_X1 U6276 ( .A1(n6017), .A2(n5776), .B1(n7078), .B2(n5330), .C1(n7022), 
        .C2(n7210), .ZN(n6214) );
  OAI21_X4 U6277 ( .B1(\UUT/Mcontrol/Nextpc_decoding/condition ), .B2(n2588), 
        .A(n2609), .ZN(n984) );
  OAI222_X4 U6278 ( .A1(n5387), .A2(n5432), .B1(n5431), .B2(n312), .C1(n5385), 
        .C2(n5430), .ZN(\UUT/branch_rega [22]) );
  INV_X1 U6279 ( .A(\UUT/branch_rega [3]), .ZN(n7358) );
  INV_X1 U6280 ( .A(\UUT/branch_rega [3]), .ZN(n7373) );
  INV_X1 U6281 ( .A(\UUT/branch_rega [3]), .ZN(n7369) );
  OAI222_X4 U6282 ( .A1(n5354), .A2(n5432), .B1(n5431), .B2(n791), .C1(n5352), 
        .C2(n5430), .ZN(\UUT/branch_rega [3]) );
  INV_X4 U6283 ( .A(\UUT/rs1_addr [4]), .ZN(n6267) );
  AND2_X2 U6284 ( .A1(n6262), .A2(n6263), .ZN(n6258) );
  AND2_X1 U6285 ( .A1(\UUT/Mpath/out_regA[21] ), .A2(\UUT/Mpath/out_regB[21] ), 
        .ZN(\UUT/Mpath/the_alu/N104 ) );
  OR2_X1 U6286 ( .A1(\UUT/Mpath/out_regA[21] ), .A2(\UUT/Mpath/out_regB[21] ), 
        .ZN(\UUT/Mpath/the_alu/N136 ) );
  OR2_X4 U6287 ( .A1(n7209), .A2(\UUT/Mcontrol/Operation_decoding32/N1882 ), 
        .ZN(\UUT/Mcontrol/Operation_decoding32/N1871 ) );
  NAND2_X4 U6288 ( .A1(\UUT/byp_controlA[2] ), .A2(\UUT/Mcontrol/st_logic/N47 ), .ZN(n5430) );
  OR2_X1 U6289 ( .A1(\UUT/rs1_addr [3]), .A2(\UUT/rs1_addr [4]), .ZN(
        \UUT/regfile/N260 ) );
  AND3_X4 U6290 ( .A1(n6270), .A2(\UUT/rs1_addr [3]), .A3(n6266), .ZN(n5451)
         );
  AND2_X1 U6291 ( .A1(n7112), .A2(n7125), .ZN(\UUT/Mpath/the_alu/N110 ) );
  OR2_X1 U6292 ( .A1(n7112), .A2(n7125), .ZN(\UUT/Mpath/the_alu/N142 ) );
  AND2_X4 U6293 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1871 ), .A2(
        \UUT/Mcontrol/d_sampled_finstr [25]), .ZN(\UUT/rs1_addr [4]) );
  NAND2_X2 U6294 ( .A1(\UUT/Mcontrol/Operation_decoding32/N1871 ), .A2(n5768), 
        .ZN(\UUT/rs1_addr [2]) );
  NAND2_X4 U6295 ( .A1(\UUT/byp_controlA[2] ), .A2(\UUT/byp_controlA[0] ), 
        .ZN(n5432) );
  NAND2_X2 U6296 ( .A1(\UUT/Mcontrol/d_sampled_finstr [22]), .A2(
        \UUT/Mcontrol/Operation_decoding32/N1871 ), .ZN(n7370) );
  INV_X1 U6297 ( .A(\UUT/Mcontrol/Operation_decoding32/N1871 ), .ZN(n6279) );
  INV_X8 U6298 ( .A(n940), .ZN(n5431) );
  OR2_X1 U6299 ( .A1(\UUT/rs1_addr [2]), .A2(\UUT/regfile/N260 ), .ZN(
        \UUT/regfile/N261 ) );
  OAI22_X2 U6300 ( .A1(\UUT/Mcontrol/Nextpc_decoding/N22 ), .A2(n6244), .B1(
        \UUT/Mcontrol/Nextpc_decoding/N266 ), .B2(n6245), .ZN(
        \UUT/Mcontrol/Nextpc_decoding/condition ) );
  AND2_X1 U6301 ( .A1(\UUT/Mpath/out_regA[18] ), .A2(n7135), .ZN(
        \UUT/Mpath/the_alu/N107 ) );
  OR2_X1 U6302 ( .A1(\UUT/Mpath/out_regA[18] ), .A2(n7135), .ZN(
        \UUT/Mpath/the_alu/N139 ) );
  OR2_X1 U6303 ( .A1(\UUT/Mcontrol/d_sampled_finstr [31]), .A2(
        \UUT/Mcontrol/d_sampled_finstr [30]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2056 ) );
  OR2_X1 U6304 ( .A1(n7205), .A2(\UUT/Mcontrol/d_instr [31]), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N2008 ) );
  OR2_X1 U6305 ( .A1(n7205), .A2(n7201), .ZN(
        \UUT/Mcontrol/Operation_decoding32/N1916 ) );
  NAND2_X4 U6306 ( .A1(n6276), .A2(n6273), .ZN(n5460) );
  NAND3_X4 U6307 ( .A1(\UUT/rs1_addr [1]), .A2(n6263), .A3(n6274), .ZN(n5454)
         );
  NOR2_X1 U6308 ( .A1(n2587), .A2(n2588), .ZN(n7380) );
  NOR2_X2 U6309 ( .A1(\UUT/Mcontrol/Nextpc_decoding/condition ), .A2(n7381), 
        .ZN(n983) );
  INV_X1 U6310 ( .A(n7380), .ZN(n7381) );
  AND2_X1 U6311 ( .A1(\UUT/Mpath/out_regA[17] ), .A2(n7197), .ZN(
        \UUT/Mpath/the_alu/N108 ) );
  OR2_X1 U6312 ( .A1(\UUT/Mpath/out_regA[17] ), .A2(n7197), .ZN(
        \UUT/Mpath/the_alu/N140 ) );
  AND2_X1 U6313 ( .A1(\UUT/Mpath/out_regA[13] ), .A2(n7122), .ZN(
        \UUT/Mpath/the_alu/N112 ) );
  OR2_X1 U6314 ( .A1(n1245), .A2(n7122), .ZN(\UUT/Mpath/the_alu/N144 ) );
  AND2_X1 U6315 ( .A1(\UUT/Mpath/out_regA[7] ), .A2(\UUT/Mpath/out_regB[7] ), 
        .ZN(\UUT/Mpath/the_alu/N118 ) );
  OR2_X1 U6316 ( .A1(\UUT/Mpath/out_regA[7] ), .A2(\UUT/Mpath/out_regB[7] ), 
        .ZN(\UUT/Mpath/the_alu/N150 ) );
  AND2_X1 U6317 ( .A1(n7198), .A2(n7107), .ZN(\UUT/Mpath/the_alu/N114 ) );
  OR2_X1 U6318 ( .A1(n7198), .A2(n7107), .ZN(\UUT/Mpath/the_alu/N146 ) );
  AND2_X1 U6319 ( .A1(n7138), .A2(n7194), .ZN(\UUT/Mpath/the_alu/N105 ) );
  OR2_X1 U6320 ( .A1(n7138), .A2(n7194), .ZN(\UUT/Mpath/the_alu/N137 ) );
  AND2_X1 U6321 ( .A1(n7129), .A2(n7136), .ZN(\UUT/Mpath/the_alu/N109 ) );
  OR2_X1 U6322 ( .A1(n7129), .A2(n7136), .ZN(\UUT/Mpath/the_alu/N141 ) );
  AND2_X1 U6323 ( .A1(n7132), .A2(n7128), .ZN(\UUT/Mpath/the_alu/N116 ) );
  OR2_X1 U6324 ( .A1(n7132), .A2(n7128), .ZN(\UUT/Mpath/the_alu/N148 ) );
  AND2_X1 U6325 ( .A1(n7193), .A2(n7134), .ZN(\UUT/Mpath/the_alu/N113 ) );
  OR2_X1 U6326 ( .A1(n7193), .A2(n7134), .ZN(\UUT/Mpath/the_alu/N145 ) );
  AND2_X1 U6327 ( .A1(n7106), .A2(n7099), .ZN(\UUT/Mpath/the_alu/N119 ) );
  OR2_X1 U6328 ( .A1(n7106), .A2(n7099), .ZN(\UUT/Mpath/the_alu/N151 ) );
  AND2_X1 U6329 ( .A1(n7113), .A2(n7140), .ZN(\UUT/Mpath/the_alu/N111 ) );
  OR2_X1 U6330 ( .A1(n7113), .A2(n7140), .ZN(\UUT/Mpath/the_alu/N143 ) );
  AND2_X1 U6331 ( .A1(n7189), .A2(\UUT/Mpath/out_regB[8] ), .ZN(
        \UUT/Mpath/the_alu/N117 ) );
  OR2_X1 U6332 ( .A1(n7189), .A2(\UUT/Mpath/out_regB[8] ), .ZN(
        \UUT/Mpath/the_alu/N149 ) );
  INV_X1 U6333 ( .A(n7303), .ZN(\UUT/Mcontrol/Nextpc_decoding/N159 ) );
  AND2_X1 U6334 ( .A1(\UUT/Mpath/out_regA[10] ), .A2(n7137), .ZN(
        \UUT/Mpath/the_alu/N115 ) );
  OR2_X1 U6335 ( .A1(\UUT/Mpath/out_regA[10] ), .A2(n7137), .ZN(
        \UUT/Mpath/the_alu/N147 ) );
  AND2_X1 U6336 ( .A1(\UUT/Mpath/out_regA[5] ), .A2(n7114), .ZN(
        \UUT/Mpath/the_alu/N120 ) );
  OR2_X1 U6337 ( .A1(\UUT/Mpath/out_regA[5] ), .A2(n7114), .ZN(
        \UUT/Mpath/the_alu/N152 ) );
  NOR2_X4 U6338 ( .A1(n7213), .A2(n2239), .ZN(n1223) );
  CLKBUF_X1 U6339 ( .A(n122), .Z(n7382) );
  CLKBUF_X1 U6340 ( .A(n122), .Z(n7383) );
  CLKBUF_X1 U6341 ( .A(n122), .Z(n7384) );
  CLKBUF_X1 U6342 ( .A(n122), .Z(n7385) );
  CLKBUF_X1 U6343 ( .A(n122), .Z(n7386) );
  CLKBUF_X1 U6344 ( .A(n122), .Z(n7387) );
  CLKBUF_X1 U6345 ( .A(n122), .Z(n7388) );
  CLKBUF_X1 U6346 ( .A(n122), .Z(n7389) );
  CLKBUF_X1 U6347 ( .A(n122), .Z(n7390) );
  CLKBUF_X1 U6348 ( .A(n122), .Z(n7391) );
  CLKBUF_X1 U6349 ( .A(n122), .Z(n7392) );
  CLKBUF_X1 U6350 ( .A(n122), .Z(n7393) );
  CLKBUF_X1 U6351 ( .A(n122), .Z(n7394) );
  CLKBUF_X1 U6352 ( .A(n122), .Z(n7395) );
  CLKBUF_X1 U6353 ( .A(n122), .Z(n7396) );
  CLKBUF_X1 U6354 ( .A(n122), .Z(n7397) );
  CLKBUF_X1 U6355 ( .A(n122), .Z(n7398) );
  CLKBUF_X3 U6356 ( .A(\UUT/Mpath/out_regB[4] ), .Z(n7399) );
  CLKBUF_X3 U6357 ( .A(\UUT/Mpath/out_regB[4] ), .Z(n7400) );
  CLKBUF_X1 U6358 ( .A(\UUT/Mpath/out_regB[2] ), .Z(n7403) );
  CLKBUF_X1 U6359 ( .A(\UUT/Mpath/out_regB[2] ), .Z(n7404) );
  CLKBUF_X3 U6360 ( .A(\UUT/Mpath/out_regB[1] ), .Z(n7405) );
  CLKBUF_X3 U6361 ( .A(\UUT/Mpath/out_regB[1] ), .Z(n7406) );
  CLKBUF_X3 U6362 ( .A(\UUT/Mpath/out_regB[0] ), .Z(n7407) );
  CLKBUF_X3 U6363 ( .A(\UUT/Mpath/out_regB[0] ), .Z(n7408) );
  XNOR2_X1 U6364 ( .A(\UUT/Mcontrol/x_rd[0] ), .B(\UUT/rs2_addr [0]), .ZN(
        n7411) );
  XNOR2_X1 U6365 ( .A(\UUT/Mcontrol/x_rd[2] ), .B(\UUT/rs2_addr [2]), .ZN(
        n7410) );
  XNOR2_X1 U6366 ( .A(\UUT/Mcontrol/x_rd[1] ), .B(\UUT/rs2_addr [1]), .ZN(
        n7409) );
  NAND3_X1 U6367 ( .A1(n7411), .A2(n7410), .A3(n7409), .ZN(n7414) );
  XOR2_X1 U6368 ( .A(\UUT/Mcontrol/x_rd[3] ), .B(\UUT/rs2_addr [3]), .Z(n7413)
         );
  XOR2_X1 U6369 ( .A(\UUT/Mcontrol/x_rd[4] ), .B(\UUT/rs2_addr [4]), .Z(n7412)
         );
  NOR3_X1 U6370 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(
        \UUT/Mcontrol/bp_logicB/N2 ) );
  XNOR2_X1 U6371 ( .A(\UUT/Mcontrol/m_sampled_xrd[0] ), .B(\UUT/rs2_addr [0]), 
        .ZN(n7417) );
  XNOR2_X1 U6372 ( .A(\UUT/Mcontrol/m_sampled_xrd[2] ), .B(\UUT/rs2_addr [2]), 
        .ZN(n7416) );
  XNOR2_X1 U6373 ( .A(\UUT/Mcontrol/m_sampled_xrd[1] ), .B(\UUT/rs2_addr [1]), 
        .ZN(n7415) );
  NAND3_X1 U6374 ( .A1(n7417), .A2(n7416), .A3(n7415), .ZN(n7420) );
  XOR2_X1 U6375 ( .A(\UUT/Mcontrol/m_sampled_xrd[3] ), .B(\UUT/rs2_addr [3]), 
        .Z(n7419) );
  XOR2_X1 U6376 ( .A(\UUT/Mcontrol/m_sampled_xrd[4] ), .B(\UUT/rs2_addr [4]), 
        .Z(n7418) );
  NOR3_X1 U6377 ( .A1(n7420), .A2(n7419), .A3(n7418), .ZN(
        \UUT/Mcontrol/bp_logicB/N3 ) );
  XNOR2_X1 U6378 ( .A(\UUT/Mcontrol/x_rd[0] ), .B(\UUT/rs1_addr [0]), .ZN(
        n7423) );
  XNOR2_X1 U6379 ( .A(\UUT/Mcontrol/x_rd[2] ), .B(\UUT/rs1_addr [2]), .ZN(
        n7422) );
  XNOR2_X1 U6380 ( .A(\UUT/Mcontrol/x_rd[1] ), .B(\UUT/rs1_addr [1]), .ZN(
        n7421) );
  NAND3_X1 U6381 ( .A1(n7423), .A2(n7422), .A3(n7421), .ZN(n7426) );
  XOR2_X1 U6382 ( .A(\UUT/Mcontrol/x_rd[3] ), .B(\UUT/rs1_addr [3]), .Z(n7425)
         );
  XOR2_X1 U6383 ( .A(\UUT/Mcontrol/x_rd[4] ), .B(\UUT/rs1_addr [4]), .Z(n7424)
         );
  NOR3_X1 U6384 ( .A1(n7426), .A2(n7425), .A3(n7424), .ZN(
        \UUT/Mcontrol/bp_logicA/N2 ) );
  XNOR2_X1 U6385 ( .A(\UUT/Mcontrol/m_sampled_xrd[0] ), .B(\UUT/rs1_addr [0]), 
        .ZN(n7429) );
  XNOR2_X1 U6386 ( .A(\UUT/Mcontrol/m_sampled_xrd[2] ), .B(\UUT/rs1_addr [2]), 
        .ZN(n7428) );
  XNOR2_X1 U6387 ( .A(\UUT/Mcontrol/m_sampled_xrd[1] ), .B(\UUT/rs1_addr [1]), 
        .ZN(n7427) );
  NAND3_X1 U6388 ( .A1(n7429), .A2(n7428), .A3(n7427), .ZN(n7432) );
  XOR2_X1 U6389 ( .A(\UUT/Mcontrol/m_sampled_xrd[3] ), .B(\UUT/rs1_addr [3]), 
        .Z(n7431) );
  XOR2_X1 U6390 ( .A(\UUT/Mcontrol/m_sampled_xrd[4] ), .B(\UUT/rs1_addr [4]), 
        .Z(n7430) );
  NOR3_X1 U6391 ( .A1(n7432), .A2(n7431), .A3(n7430), .ZN(
        \UUT/Mcontrol/bp_logicA/N3 ) );
endmodule

