##
## LEF for PtnCells ;
## created by Encounter v09.10-p004_1 on Mon Mar  3 19:07:24 2014
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO up_island
  CLASS BLOCK ;
  SIZE 184.6000 BY 184.4600 ;
  FOREIGN up_island 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.0600 184.3900 76.1300 184.4600 ;
    END
  END CLK
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.0100 184.3900 77.0800 184.4600 ;
    END
  END reset
  PIN BUS_NREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.9600 184.3900 78.0300 184.4600 ;
    END
  END BUS_NREADY
  PIN BUS_BUSY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.5100 0.0000 29.5800 0.0700 ;
    END
  END BUS_BUSY
  PIN BUS_MR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.3100 0.0000 33.3800 0.0700 ;
    END
  END BUS_MR
  PIN BUS_MW
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.4100 0.0000 31.4800 0.0700 ;
    END
  END BUS_MW
  PIN BUS_ADDR_OUTBUS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.1100 0.0000 94.1800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[31]
  PIN BUS_ADDR_OUTBUS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.2100 0.0000 92.2800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[30]
  PIN BUS_ADDR_OUTBUS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.3100 0.0000 90.3800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[29]
  PIN BUS_ADDR_OUTBUS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.4100 0.0000 88.4800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[28]
  PIN BUS_ADDR_OUTBUS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.5100 0.0000 86.5800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[27]
  PIN BUS_ADDR_OUTBUS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.6100 0.0000 84.6800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[26]
  PIN BUS_ADDR_OUTBUS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.7100 0.0000 82.7800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[25]
  PIN BUS_ADDR_OUTBUS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.8100 0.0000 80.8800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[24]
  PIN BUS_ADDR_OUTBUS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.9100 0.0000 78.9800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[23]
  PIN BUS_ADDR_OUTBUS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.0100 0.0000 77.0800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[22]
  PIN BUS_ADDR_OUTBUS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.1100 0.0000 75.1800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[21]
  PIN BUS_ADDR_OUTBUS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.2100 0.0000 73.2800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[20]
  PIN BUS_ADDR_OUTBUS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.3100 0.0000 71.3800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[19]
  PIN BUS_ADDR_OUTBUS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.4100 0.0000 69.4800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[18]
  PIN BUS_ADDR_OUTBUS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.5100 0.0000 67.5800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[17]
  PIN BUS_ADDR_OUTBUS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.6100 0.0000 65.6800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[16]
  PIN BUS_ADDR_OUTBUS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.7100 0.0000 63.7800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[15]
  PIN BUS_ADDR_OUTBUS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.8100 0.0000 61.8800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[14]
  PIN BUS_ADDR_OUTBUS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.9100 0.0000 59.9800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[13]
  PIN BUS_ADDR_OUTBUS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.0100 0.0000 58.0800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[12]
  PIN BUS_ADDR_OUTBUS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.1100 0.0000 56.1800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[11]
  PIN BUS_ADDR_OUTBUS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.2100 0.0000 54.2800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[10]
  PIN BUS_ADDR_OUTBUS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.3100 0.0000 52.3800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[9]
  PIN BUS_ADDR_OUTBUS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.4100 0.0000 50.4800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[8]
  PIN BUS_ADDR_OUTBUS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.5100 0.0000 48.5800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[7]
  PIN BUS_ADDR_OUTBUS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.6100 0.0000 46.6800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[6]
  PIN BUS_ADDR_OUTBUS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.7100 0.0000 44.7800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[5]
  PIN BUS_ADDR_OUTBUS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.8100 0.0000 42.8800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[4]
  PIN BUS_ADDR_OUTBUS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.9100 0.0000 40.9800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[3]
  PIN BUS_ADDR_OUTBUS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.0100 0.0000 39.0800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[2]
  PIN BUS_ADDR_OUTBUS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.1100 0.0000 37.1800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[1]
  PIN BUS_ADDR_OUTBUS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.2100 0.0000 35.2800 0.0700 ;
    END
  END BUS_ADDR_OUTBUS[0]
  PIN BUS_DATA_INBUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.3600 184.3900 108.4300 184.4600 ;
    END
  END BUS_DATA_INBUS[31]
  PIN BUS_DATA_INBUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.4100 184.3900 107.4800 184.4600 ;
    END
  END BUS_DATA_INBUS[30]
  PIN BUS_DATA_INBUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.4600 184.3900 106.5300 184.4600 ;
    END
  END BUS_DATA_INBUS[29]
  PIN BUS_DATA_INBUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.5100 184.3900 105.5800 184.4600 ;
    END
  END BUS_DATA_INBUS[28]
  PIN BUS_DATA_INBUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.5600 184.3900 104.6300 184.4600 ;
    END
  END BUS_DATA_INBUS[27]
  PIN BUS_DATA_INBUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.6100 184.3900 103.6800 184.4600 ;
    END
  END BUS_DATA_INBUS[26]
  PIN BUS_DATA_INBUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.6600 184.3900 102.7300 184.4600 ;
    END
  END BUS_DATA_INBUS[25]
  PIN BUS_DATA_INBUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.7100 184.3900 101.7800 184.4600 ;
    END
  END BUS_DATA_INBUS[24]
  PIN BUS_DATA_INBUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.7600 184.3900 100.8300 184.4600 ;
    END
  END BUS_DATA_INBUS[23]
  PIN BUS_DATA_INBUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.8100 184.3900 99.8800 184.4600 ;
    END
  END BUS_DATA_INBUS[22]
  PIN BUS_DATA_INBUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.8600 184.3900 98.9300 184.4600 ;
    END
  END BUS_DATA_INBUS[21]
  PIN BUS_DATA_INBUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.9100 184.3900 97.9800 184.4600 ;
    END
  END BUS_DATA_INBUS[20]
  PIN BUS_DATA_INBUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.9600 184.3900 97.0300 184.4600 ;
    END
  END BUS_DATA_INBUS[19]
  PIN BUS_DATA_INBUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.0100 184.3900 96.0800 184.4600 ;
    END
  END BUS_DATA_INBUS[18]
  PIN BUS_DATA_INBUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.0600 184.3900 95.1300 184.4600 ;
    END
  END BUS_DATA_INBUS[17]
  PIN BUS_DATA_INBUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.1100 184.3900 94.1800 184.4600 ;
    END
  END BUS_DATA_INBUS[16]
  PIN BUS_DATA_INBUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.1600 184.3900 93.2300 184.4600 ;
    END
  END BUS_DATA_INBUS[15]
  PIN BUS_DATA_INBUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.2100 184.3900 92.2800 184.4600 ;
    END
  END BUS_DATA_INBUS[14]
  PIN BUS_DATA_INBUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.2600 184.3900 91.3300 184.4600 ;
    END
  END BUS_DATA_INBUS[13]
  PIN BUS_DATA_INBUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.3100 184.3900 90.3800 184.4600 ;
    END
  END BUS_DATA_INBUS[12]
  PIN BUS_DATA_INBUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.3600 184.3900 89.4300 184.4600 ;
    END
  END BUS_DATA_INBUS[11]
  PIN BUS_DATA_INBUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.4100 184.3900 88.4800 184.4600 ;
    END
  END BUS_DATA_INBUS[10]
  PIN BUS_DATA_INBUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.4600 184.3900 87.5300 184.4600 ;
    END
  END BUS_DATA_INBUS[9]
  PIN BUS_DATA_INBUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.5100 184.3900 86.5800 184.4600 ;
    END
  END BUS_DATA_INBUS[8]
  PIN BUS_DATA_INBUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.5600 184.3900 85.6300 184.4600 ;
    END
  END BUS_DATA_INBUS[7]
  PIN BUS_DATA_INBUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.6100 184.3900 84.6800 184.4600 ;
    END
  END BUS_DATA_INBUS[6]
  PIN BUS_DATA_INBUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.6600 184.3900 83.7300 184.4600 ;
    END
  END BUS_DATA_INBUS[5]
  PIN BUS_DATA_INBUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.7100 184.3900 82.7800 184.4600 ;
    END
  END BUS_DATA_INBUS[4]
  PIN BUS_DATA_INBUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.7600 184.3900 81.8300 184.4600 ;
    END
  END BUS_DATA_INBUS[3]
  PIN BUS_DATA_INBUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.8100 184.3900 80.8800 184.4600 ;
    END
  END BUS_DATA_INBUS[2]
  PIN BUS_DATA_INBUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.8600 184.3900 79.9300 184.4600 ;
    END
  END BUS_DATA_INBUS[1]
  PIN BUS_DATA_INBUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.9100 184.3900 78.9800 184.4600 ;
    END
  END BUS_DATA_INBUS[0]
  PIN BUS_DATA_OUTBUS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 154.9100 0.0000 154.9800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[31]
  PIN BUS_DATA_OUTBUS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 153.0100 0.0000 153.0800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[30]
  PIN BUS_DATA_OUTBUS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 151.1100 0.0000 151.1800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[29]
  PIN BUS_DATA_OUTBUS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.2100 0.0000 149.2800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[28]
  PIN BUS_DATA_OUTBUS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 147.3100 0.0000 147.3800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[27]
  PIN BUS_DATA_OUTBUS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.4100 0.0000 145.4800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[26]
  PIN BUS_DATA_OUTBUS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 143.5100 0.0000 143.5800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[25]
  PIN BUS_DATA_OUTBUS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.6100 0.0000 141.6800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[24]
  PIN BUS_DATA_OUTBUS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.7100 0.0000 139.7800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[23]
  PIN BUS_DATA_OUTBUS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 137.8100 0.0000 137.8800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[22]
  PIN BUS_DATA_OUTBUS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 135.9100 0.0000 135.9800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[21]
  PIN BUS_DATA_OUTBUS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 134.0100 0.0000 134.0800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[20]
  PIN BUS_DATA_OUTBUS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.1100 0.0000 132.1800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[19]
  PIN BUS_DATA_OUTBUS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.2100 0.0000 130.2800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[18]
  PIN BUS_DATA_OUTBUS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 128.3100 0.0000 128.3800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[17]
  PIN BUS_DATA_OUTBUS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.4100 0.0000 126.4800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[16]
  PIN BUS_DATA_OUTBUS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 124.5100 0.0000 124.5800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[15]
  PIN BUS_DATA_OUTBUS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.6100 0.0000 122.6800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[14]
  PIN BUS_DATA_OUTBUS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.7100 0.0000 120.7800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[13]
  PIN BUS_DATA_OUTBUS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.8100 0.0000 118.8800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[12]
  PIN BUS_DATA_OUTBUS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.9100 0.0000 116.9800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[11]
  PIN BUS_DATA_OUTBUS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.0100 0.0000 115.0800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[10]
  PIN BUS_DATA_OUTBUS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.1100 0.0000 113.1800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[9]
  PIN BUS_DATA_OUTBUS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.2100 0.0000 111.2800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[8]
  PIN BUS_DATA_OUTBUS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.3100 0.0000 109.3800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[7]
  PIN BUS_DATA_OUTBUS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.4100 0.0000 107.4800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[6]
  PIN BUS_DATA_OUTBUS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.5100 0.0000 105.5800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[5]
  PIN BUS_DATA_OUTBUS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.6100 0.0000 103.6800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[4]
  PIN BUS_DATA_OUTBUS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.7100 0.0000 101.7800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[3]
  PIN BUS_DATA_OUTBUS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.8100 0.0000 99.8800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[2]
  PIN BUS_DATA_OUTBUS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.9100 0.0000 97.9800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[1]
  PIN BUS_DATA_OUTBUS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.0100 0.0000 96.0800 0.0700 ;
    END
  END BUS_DATA_OUTBUS[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal10 ;
        RECT 2.3800 0.0000 3.1800 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.3800 183.6600 3.1800 184.4600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 181.5000 0.0000 182.3000 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 181.5000 183.6600 182.3000 184.4600 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal10 ;
        RECT 0.7800 0.0000 1.5800 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 0.7800 183.6600 1.5800 184.4600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 183.1000 0.0000 183.9000 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 183.1000 183.6600 183.9000 184.4600 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal2 ;
      RECT 108.5000 184.3200 184.6000 184.4600 ;
      RECT 107.5500 184.3200 108.2900 184.4600 ;
      RECT 106.6000 184.3200 107.3400 184.4600 ;
      RECT 105.6500 184.3200 106.3900 184.4600 ;
      RECT 104.7000 184.3200 105.4400 184.4600 ;
      RECT 103.7500 184.3200 104.4900 184.4600 ;
      RECT 102.8000 184.3200 103.5400 184.4600 ;
      RECT 101.8500 184.3200 102.5900 184.4600 ;
      RECT 100.9000 184.3200 101.6400 184.4600 ;
      RECT 99.9500 184.3200 100.6900 184.4600 ;
      RECT 99.0000 184.3200 99.7400 184.4600 ;
      RECT 98.0500 184.3200 98.7900 184.4600 ;
      RECT 97.1000 184.3200 97.8400 184.4600 ;
      RECT 96.1500 184.3200 96.8900 184.4600 ;
      RECT 95.2000 184.3200 95.9400 184.4600 ;
      RECT 94.2500 184.3200 94.9900 184.4600 ;
      RECT 93.3000 184.3200 94.0400 184.4600 ;
      RECT 92.3500 184.3200 93.0900 184.4600 ;
      RECT 91.4000 184.3200 92.1400 184.4600 ;
      RECT 90.4500 184.3200 91.1900 184.4600 ;
      RECT 89.5000 184.3200 90.2400 184.4600 ;
      RECT 88.5500 184.3200 89.2900 184.4600 ;
      RECT 87.6000 184.3200 88.3400 184.4600 ;
      RECT 86.6500 184.3200 87.3900 184.4600 ;
      RECT 85.7000 184.3200 86.4400 184.4600 ;
      RECT 84.7500 184.3200 85.4900 184.4600 ;
      RECT 83.8000 184.3200 84.5400 184.4600 ;
      RECT 82.8500 184.3200 83.5900 184.4600 ;
      RECT 81.9000 184.3200 82.6400 184.4600 ;
      RECT 80.9500 184.3200 81.6900 184.4600 ;
      RECT 80.0000 184.3200 80.7400 184.4600 ;
      RECT 79.0500 184.3200 79.7900 184.4600 ;
      RECT 78.1000 184.3200 78.8400 184.4600 ;
      RECT 77.1500 184.3200 77.8900 184.4600 ;
      RECT 76.2000 184.3200 76.9400 184.4600 ;
      RECT 0.0000 184.3200 75.9900 184.4600 ;
      RECT 0.0000 0.1400 184.6000 184.3200 ;
      RECT 155.0500 0.0000 184.6000 0.1400 ;
      RECT 153.1500 0.0000 154.8400 0.1400 ;
      RECT 151.2500 0.0000 152.9400 0.1400 ;
      RECT 149.3500 0.0000 151.0400 0.1400 ;
      RECT 147.4500 0.0000 149.1400 0.1400 ;
      RECT 145.5500 0.0000 147.2400 0.1400 ;
      RECT 143.6500 0.0000 145.3400 0.1400 ;
      RECT 141.7500 0.0000 143.4400 0.1400 ;
      RECT 139.8500 0.0000 141.5400 0.1400 ;
      RECT 137.9500 0.0000 139.6400 0.1400 ;
      RECT 136.0500 0.0000 137.7400 0.1400 ;
      RECT 134.1500 0.0000 135.8400 0.1400 ;
      RECT 132.2500 0.0000 133.9400 0.1400 ;
      RECT 130.3500 0.0000 132.0400 0.1400 ;
      RECT 128.4500 0.0000 130.1400 0.1400 ;
      RECT 126.5500 0.0000 128.2400 0.1400 ;
      RECT 124.6500 0.0000 126.3400 0.1400 ;
      RECT 122.7500 0.0000 124.4400 0.1400 ;
      RECT 120.8500 0.0000 122.5400 0.1400 ;
      RECT 118.9500 0.0000 120.6400 0.1400 ;
      RECT 117.0500 0.0000 118.7400 0.1400 ;
      RECT 115.1500 0.0000 116.8400 0.1400 ;
      RECT 113.2500 0.0000 114.9400 0.1400 ;
      RECT 111.3500 0.0000 113.0400 0.1400 ;
      RECT 109.4500 0.0000 111.1400 0.1400 ;
      RECT 107.5500 0.0000 109.2400 0.1400 ;
      RECT 105.6500 0.0000 107.3400 0.1400 ;
      RECT 103.7500 0.0000 105.4400 0.1400 ;
      RECT 101.8500 0.0000 103.5400 0.1400 ;
      RECT 99.9500 0.0000 101.6400 0.1400 ;
      RECT 98.0500 0.0000 99.7400 0.1400 ;
      RECT 96.1500 0.0000 97.8400 0.1400 ;
      RECT 94.2500 0.0000 95.9400 0.1400 ;
      RECT 92.3500 0.0000 94.0400 0.1400 ;
      RECT 90.4500 0.0000 92.1400 0.1400 ;
      RECT 88.5500 0.0000 90.2400 0.1400 ;
      RECT 86.6500 0.0000 88.3400 0.1400 ;
      RECT 84.7500 0.0000 86.4400 0.1400 ;
      RECT 82.8500 0.0000 84.5400 0.1400 ;
      RECT 80.9500 0.0000 82.6400 0.1400 ;
      RECT 79.0500 0.0000 80.7400 0.1400 ;
      RECT 77.1500 0.0000 78.8400 0.1400 ;
      RECT 75.2500 0.0000 76.9400 0.1400 ;
      RECT 73.3500 0.0000 75.0400 0.1400 ;
      RECT 71.4500 0.0000 73.1400 0.1400 ;
      RECT 69.5500 0.0000 71.2400 0.1400 ;
      RECT 67.6500 0.0000 69.3400 0.1400 ;
      RECT 65.7500 0.0000 67.4400 0.1400 ;
      RECT 63.8500 0.0000 65.5400 0.1400 ;
      RECT 61.9500 0.0000 63.6400 0.1400 ;
      RECT 60.0500 0.0000 61.7400 0.1400 ;
      RECT 58.1500 0.0000 59.8400 0.1400 ;
      RECT 56.2500 0.0000 57.9400 0.1400 ;
      RECT 54.3500 0.0000 56.0400 0.1400 ;
      RECT 52.4500 0.0000 54.1400 0.1400 ;
      RECT 50.5500 0.0000 52.2400 0.1400 ;
      RECT 48.6500 0.0000 50.3400 0.1400 ;
      RECT 46.7500 0.0000 48.4400 0.1400 ;
      RECT 44.8500 0.0000 46.5400 0.1400 ;
      RECT 42.9500 0.0000 44.6400 0.1400 ;
      RECT 41.0500 0.0000 42.7400 0.1400 ;
      RECT 39.1500 0.0000 40.8400 0.1400 ;
      RECT 37.2500 0.0000 38.9400 0.1400 ;
      RECT 35.3500 0.0000 37.0400 0.1400 ;
      RECT 33.4500 0.0000 35.1400 0.1400 ;
      RECT 31.5500 0.0000 33.2400 0.1400 ;
      RECT 29.6500 0.0000 31.3400 0.1400 ;
      RECT 0.0000 0.0000 29.4400 0.1400 ;
    LAYER metal3 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal4 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal5 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal6 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal7 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal8 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal9 ;
      RECT 0.0000 0.0000 184.6000 184.4600 ;
    LAYER metal10 ;
      RECT 3.9800 182.8600 180.7000 184.4600 ;
      RECT 0.0000 1.6000 184.6000 182.8600 ;
      RECT 3.9800 0.0000 180.7000 1.6000 ;
  END
END up_island

END LIBRARY
