
module Xi_core_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n67, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n91,
         n92, n93, n94, n95, n96;

  NOR2_X4 U26 ( .A1(n27), .A2(n26), .ZN(n25) );
  XNOR2_X2 U28 ( .A(n76), .B(A[20]), .ZN(n27) );
  NAND2_X4 U29 ( .A1(n32), .A2(n29), .ZN(n28) );
  NOR2_X4 U30 ( .A1(n31), .A2(n30), .ZN(n29) );
  XNOR2_X2 U34 ( .A(n79), .B(A[17]), .ZN(n33) );
  NAND2_X4 U38 ( .A1(n40), .A2(n37), .ZN(n36) );
  XNOR2_X2 U43 ( .A(n83), .B(A[13]), .ZN(n41) );
  NAND2_X4 U53 ( .A1(n55), .A2(n52), .ZN(n51) );
  NAND2_X4 U60 ( .A1(n62), .A2(n59), .ZN(n58) );
  XNOR2_X2 U65 ( .A(n95), .B(A[1]), .ZN(n63) );
  XNOR2_X1 U102 ( .A(n92), .B(A[4]), .ZN(n57) );
  BUF_X2 U103 ( .A(n1), .Z(NE) );
  XNOR2_X2 U104 ( .A(n77), .B(A[19]), .ZN(n30) );
  XOR2_X1 U105 ( .A(B[31]), .B(A[31]), .Z(n10) );
  XOR2_X1 U106 ( .A(B[30]), .B(A[30]), .Z(n11) );
  INV_X1 U107 ( .A(B[22]), .ZN(n74) );
  NOR2_X1 U108 ( .A1(n46), .A2(n45), .ZN(n44) );
  NOR2_X1 U109 ( .A1(n14), .A2(n13), .ZN(n12) );
  NAND2_X1 U110 ( .A1(n3), .A2(n7), .ZN(n6) );
  NOR2_X1 U111 ( .A1(n24), .A2(n23), .ZN(n22) );
  XNOR2_X1 U112 ( .A(n70), .B(A[26]), .ZN(n17) );
  XNOR2_X1 U113 ( .A(n75), .B(A[21]), .ZN(n26) );
  NOR2_X2 U114 ( .A1(n28), .A2(n21), .ZN(n3) );
  NAND2_X1 U115 ( .A1(n25), .A2(n22), .ZN(n21) );
  NAND2_X1 U116 ( .A1(n47), .A2(n44), .ZN(n43) );
  CLKBUF_X1 U117 ( .A(n5), .Z(EQ) );
  XNOR2_X1 U118 ( .A(n71), .B(A[25]), .ZN(n19) );
  XOR2_X1 U119 ( .A(B[10]), .B(A[10]), .Z(n46) );
  NOR2_X2 U120 ( .A1(n4), .A2(n8), .ZN(n7) );
  INV_X1 U121 ( .A(B[27]), .ZN(n69) );
  XOR2_X1 U122 ( .A(B[28]), .B(A[28]), .Z(n14) );
  XOR2_X1 U123 ( .A(B[6]), .B(A[6]), .Z(n54) );
  NAND2_X1 U124 ( .A1(n18), .A2(n15), .ZN(n4) );
  NOR2_X1 U125 ( .A1(n17), .A2(n16), .ZN(n15) );
  XNOR2_X1 U126 ( .A(n74), .B(A[22]), .ZN(n24) );
  XNOR2_X1 U127 ( .A(n69), .B(A[27]), .ZN(n16) );
  NOR2_X2 U128 ( .A1(n64), .A2(n63), .ZN(n62) );
  XNOR2_X1 U129 ( .A(n96), .B(A[0]), .ZN(n64) );
  INV_X1 U130 ( .A(B[0]), .ZN(n96) );
  NOR2_X2 U131 ( .A1(n49), .A2(n48), .ZN(n47) );
  XNOR2_X1 U132 ( .A(n88), .B(A[8]), .ZN(n49) );
  INV_X1 U133 ( .A(B[8]), .ZN(n88) );
  INV_X1 U134 ( .A(B[1]), .ZN(n95) );
  INV_X1 U135 ( .A(B[2]), .ZN(n94) );
  INV_X1 U136 ( .A(n5), .ZN(n1) );
  NOR2_X2 U137 ( .A1(n2), .A2(n6), .ZN(n5) );
  NOR2_X2 U138 ( .A1(n39), .A2(n38), .ZN(n37) );
  XNOR2_X1 U139 ( .A(n82), .B(A[14]), .ZN(n39) );
  INV_X1 U140 ( .A(B[14]), .ZN(n82) );
  INV_X1 U141 ( .A(B[20]), .ZN(n76) );
  INV_X1 U142 ( .A(B[21]), .ZN(n75) );
  NOR2_X2 U143 ( .A1(n43), .A2(n36), .ZN(n35) );
  INV_X1 U144 ( .A(B[13]), .ZN(n83) );
  INV_X1 U145 ( .A(B[16]), .ZN(n80) );
  XNOR2_X1 U146 ( .A(n80), .B(A[16]), .ZN(n34) );
  INV_X1 U147 ( .A(B[4]), .ZN(n92) );
  INV_X1 U148 ( .A(B[19]), .ZN(n77) );
  INV_X1 U149 ( .A(B[24]), .ZN(n72) );
  XNOR2_X1 U150 ( .A(n72), .B(A[24]), .ZN(n20) );
  XNOR2_X1 U151 ( .A(n78), .B(A[18]), .ZN(n31) );
  INV_X1 U152 ( .A(B[18]), .ZN(n78) );
  INV_X4 U153 ( .A(B[26]), .ZN(n70) );
  NOR2_X2 U154 ( .A1(n42), .A2(n41), .ZN(n40) );
  XNOR2_X1 U155 ( .A(n84), .B(A[12]), .ZN(n42) );
  INV_X1 U156 ( .A(B[12]), .ZN(n84) );
  NOR2_X2 U157 ( .A1(n34), .A2(n33), .ZN(n32) );
  INV_X1 U158 ( .A(B[17]), .ZN(n79) );
  NOR2_X2 U159 ( .A1(n20), .A2(n19), .ZN(n18) );
  INV_X1 U160 ( .A(B[25]), .ZN(n71) );
  INV_X1 U161 ( .A(B[7]), .ZN(n89) );
  INV_X1 U162 ( .A(B[9]), .ZN(n87) );
  NAND2_X1 U163 ( .A1(n12), .A2(n9), .ZN(n8) );
  NOR2_X1 U164 ( .A1(n11), .A2(n10), .ZN(n9) );
  XNOR2_X1 U165 ( .A(n67), .B(A[29]), .ZN(n13) );
  INV_X1 U166 ( .A(B[29]), .ZN(n67) );
  NOR2_X2 U167 ( .A1(n58), .A2(n51), .ZN(n50) );
  INV_X1 U168 ( .A(B[15]), .ZN(n81) );
  NAND2_X1 U169 ( .A1(n50), .A2(n35), .ZN(n2) );
  INV_X1 U170 ( .A(B[23]), .ZN(n73) );
  NOR2_X2 U171 ( .A1(n61), .A2(n60), .ZN(n59) );
  XNOR2_X1 U172 ( .A(n94), .B(A[2]), .ZN(n61) );
  INV_X1 U173 ( .A(B[3]), .ZN(n93) );
  XNOR2_X1 U174 ( .A(n93), .B(A[3]), .ZN(n60) );
  XNOR2_X1 U175 ( .A(n85), .B(A[11]), .ZN(n45) );
  INV_X1 U176 ( .A(B[11]), .ZN(n85) );
  NOR2_X2 U177 ( .A1(n54), .A2(n53), .ZN(n52) );
  XNOR2_X1 U178 ( .A(n89), .B(A[7]), .ZN(n53) );
  XNOR2_X1 U179 ( .A(n87), .B(A[9]), .ZN(n48) );
  NOR2_X2 U180 ( .A1(n57), .A2(n56), .ZN(n55) );
  XNOR2_X1 U181 ( .A(n91), .B(A[5]), .ZN(n56) );
  INV_X1 U182 ( .A(B[5]), .ZN(n91) );
  XNOR2_X1 U183 ( .A(n73), .B(A[23]), .ZN(n23) );
  XNOR2_X1 U184 ( .A(n81), .B(A[15]), .ZN(n38) );
endmodule


module Xi_core_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  AOI21_X4 U7 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  OAI21_X4 U9 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  NOR2_X4 U10 ( .A1(n151), .A2(B[31]), .ZN(n14) );
  NAND2_X4 U11 ( .A1(n151), .A2(B[31]), .ZN(n15) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U28 ( .A1(n34), .A2(n32), .ZN(n30) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  OAI21_X4 U35 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NAND2_X4 U50 ( .A1(n58), .A2(n52), .ZN(n50) );
  AOI21_X4 U51 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NOR2_X4 U52 ( .A1(n56), .A2(n54), .ZN(n52) );
  OAI21_X4 U53 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  NOR2_X4 U108 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  NAND2_X4 U109 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  NOR2_X4 U118 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X4 U119 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NAND2_X4 U120 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  INV_X1 U157 ( .A(A[14]), .ZN(n134) );
  AOI21_X2 U158 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  INV_X4 U159 ( .A(A[24]), .ZN(n144) );
  OAI21_X1 U160 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NAND2_X1 U161 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  AOI21_X2 U162 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  INV_X2 U163 ( .A(A[18]), .ZN(n138) );
  INV_X1 U164 ( .A(A[26]), .ZN(n146) );
  INV_X1 U165 ( .A(A[12]), .ZN(n132) );
  INV_X2 U166 ( .A(A[28]), .ZN(n148) );
  OAI21_X1 U167 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  INV_X4 U168 ( .A(A[4]), .ZN(n124) );
  OAI21_X1 U169 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X2 U170 ( .A1(n28), .A2(n26), .ZN(n24) );
  INV_X4 U171 ( .A(A[27]), .ZN(n147) );
  OAI21_X1 U172 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X1 U173 ( .A1(n22), .A2(n20), .ZN(n18) );
  INV_X4 U174 ( .A(A[29]), .ZN(n149) );
  INV_X2 U175 ( .A(A[3]), .ZN(n123) );
  INV_X1 U176 ( .A(A[23]), .ZN(n143) );
  INV_X4 U177 ( .A(A[1]), .ZN(n121) );
  INV_X4 U178 ( .A(A[0]), .ZN(n120) );
  INV_X4 U179 ( .A(A[25]), .ZN(n145) );
  INV_X4 U180 ( .A(A[2]), .ZN(n122) );
  INV_X4 U181 ( .A(A[30]), .ZN(n150) );
  INV_X4 U182 ( .A(A[22]), .ZN(n142) );
  INV_X1 U183 ( .A(A[7]), .ZN(n127) );
  INV_X1 U184 ( .A(A[10]), .ZN(n130) );
  INV_X1 U185 ( .A(A[6]), .ZN(n126) );
  INV_X2 U186 ( .A(A[13]), .ZN(n133) );
  INV_X1 U187 ( .A(A[8]), .ZN(n128) );
  INV_X1 U188 ( .A(A[19]), .ZN(n139) );
  INV_X4 U189 ( .A(A[21]), .ZN(n141) );
  INV_X4 U190 ( .A(A[31]), .ZN(n151) );
  INV_X2 U191 ( .A(A[17]), .ZN(n137) );
  INV_X1 U192 ( .A(A[5]), .ZN(n125) );
  INV_X1 U193 ( .A(A[11]), .ZN(n131) );
  NAND2_X1 U194 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X1 U195 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  NAND2_X1 U196 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X1 U197 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X1 U198 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X1 U199 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NAND2_X1 U200 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X1 U201 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  NAND2_X1 U202 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X1 U203 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NOR2_X1 U204 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X1 U205 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  NAND2_X1 U206 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X1 U207 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  INV_X2 U208 ( .A(A[9]), .ZN(n129) );
  NAND2_X1 U209 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  NOR2_X1 U210 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X1 U211 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X1 U212 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  NAND2_X1 U213 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X1 U214 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  NAND2_X1 U215 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X1 U216 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NOR2_X1 U217 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NAND2_X1 U218 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X1 U219 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X1 U220 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  NAND2_X1 U221 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X1 U222 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NOR2_X1 U223 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  NAND2_X1 U224 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  NOR2_X1 U225 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X1 U226 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  INV_X2 U227 ( .A(A[16]), .ZN(n136) );
  INV_X4 U228 ( .A(A[15]), .ZN(n135) );
  INV_X4 U229 ( .A(A[20]), .ZN(n140) );
endmodule


module Xi_core_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  NAND2_X4 U2 ( .A1(n3), .A2(n8), .ZN(n6) );
  AOI21_X4 U3 ( .B1(n2), .B2(n8), .A(n9), .ZN(n7) );
  NOR2_X4 U4 ( .A1(n5), .A2(n10), .ZN(n8) );
  OAI21_X4 U5 ( .B1(n4), .B2(n10), .A(n11), .ZN(n9) );
  NAND2_X4 U6 ( .A1(n18), .A2(n12), .ZN(n10) );
  NOR2_X4 U8 ( .A1(n16), .A2(n14), .ZN(n12) );
  NOR2_X4 U12 ( .A1(n150), .A2(B[30]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n150), .A2(B[30]), .ZN(n17) );
  NOR2_X4 U14 ( .A1(n22), .A2(n20), .ZN(n18) );
  OAI21_X4 U15 ( .B1(n20), .B2(n23), .A(n21), .ZN(n19) );
  NOR2_X4 U16 ( .A1(n149), .A2(B[29]), .ZN(n20) );
  NAND2_X4 U17 ( .A1(n149), .A2(B[29]), .ZN(n21) );
  NOR2_X4 U18 ( .A1(n148), .A2(B[28]), .ZN(n22) );
  NAND2_X4 U19 ( .A1(n148), .A2(B[28]), .ZN(n23) );
  NAND2_X4 U20 ( .A1(n30), .A2(n24), .ZN(n5) );
  AOI21_X4 U21 ( .B1(n24), .B2(n31), .A(n25), .ZN(n4) );
  NOR2_X4 U22 ( .A1(n28), .A2(n26), .ZN(n24) );
  OAI21_X4 U23 ( .B1(n26), .B2(n29), .A(n27), .ZN(n25) );
  NOR2_X4 U24 ( .A1(n147), .A2(B[27]), .ZN(n26) );
  NAND2_X4 U25 ( .A1(n147), .A2(B[27]), .ZN(n27) );
  NOR2_X4 U26 ( .A1(n146), .A2(B[26]), .ZN(n28) );
  NAND2_X4 U27 ( .A1(n146), .A2(B[26]), .ZN(n29) );
  NOR2_X4 U30 ( .A1(n145), .A2(B[25]), .ZN(n32) );
  NAND2_X4 U31 ( .A1(n145), .A2(B[25]), .ZN(n33) );
  NOR2_X4 U32 ( .A1(n144), .A2(B[24]), .ZN(n34) );
  NAND2_X4 U33 ( .A1(n144), .A2(B[24]), .ZN(n35) );
  NOR2_X4 U34 ( .A1(n50), .A2(n36), .ZN(n3) );
  NAND2_X4 U36 ( .A1(n44), .A2(n38), .ZN(n36) );
  AOI21_X4 U37 ( .B1(n38), .B2(n45), .A(n39), .ZN(n37) );
  NOR2_X4 U38 ( .A1(n42), .A2(n40), .ZN(n38) );
  OAI21_X4 U39 ( .B1(n40), .B2(n43), .A(n41), .ZN(n39) );
  NOR2_X4 U40 ( .A1(n143), .A2(B[23]), .ZN(n40) );
  NAND2_X4 U41 ( .A1(n143), .A2(B[23]), .ZN(n41) );
  NOR2_X4 U42 ( .A1(n142), .A2(B[22]), .ZN(n42) );
  NAND2_X4 U43 ( .A1(n142), .A2(B[22]), .ZN(n43) );
  NOR2_X4 U44 ( .A1(n48), .A2(n46), .ZN(n44) );
  OAI21_X4 U45 ( .B1(n46), .B2(n49), .A(n47), .ZN(n45) );
  NOR2_X4 U46 ( .A1(n141), .A2(B[21]), .ZN(n46) );
  NAND2_X4 U47 ( .A1(n141), .A2(B[21]), .ZN(n47) );
  NAND2_X4 U50 ( .A1(n58), .A2(n52), .ZN(n50) );
  AOI21_X4 U51 ( .B1(n52), .B2(n59), .A(n53), .ZN(n51) );
  NOR2_X4 U52 ( .A1(n56), .A2(n54), .ZN(n52) );
  OAI21_X4 U53 ( .B1(n54), .B2(n57), .A(n55), .ZN(n53) );
  NOR2_X4 U58 ( .A1(n62), .A2(n60), .ZN(n58) );
  OAI21_X4 U59 ( .B1(n60), .B2(n63), .A(n61), .ZN(n59) );
  AOI21_X4 U64 ( .B1(n94), .B2(n64), .A(n65), .ZN(n1) );
  NOR2_X4 U65 ( .A1(n80), .A2(n66), .ZN(n64) );
  OAI21_X4 U66 ( .B1(n81), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X4 U67 ( .A1(n74), .A2(n68), .ZN(n66) );
  AOI21_X4 U68 ( .B1(n68), .B2(n75), .A(n69), .ZN(n67) );
  NOR2_X4 U69 ( .A1(n72), .A2(n70), .ZN(n68) );
  OAI21_X4 U70 ( .B1(n70), .B2(n73), .A(n71), .ZN(n69) );
  NOR2_X4 U75 ( .A1(n78), .A2(n76), .ZN(n74) );
  OAI21_X4 U76 ( .B1(n76), .B2(n79), .A(n77), .ZN(n75) );
  NAND2_X4 U81 ( .A1(n88), .A2(n82), .ZN(n80) );
  AOI21_X4 U82 ( .B1(n82), .B2(n89), .A(n83), .ZN(n81) );
  NOR2_X4 U83 ( .A1(n86), .A2(n84), .ZN(n82) );
  OAI21_X4 U84 ( .B1(n84), .B2(n87), .A(n85), .ZN(n83) );
  NOR2_X4 U89 ( .A1(n92), .A2(n90), .ZN(n88) );
  OAI21_X4 U90 ( .B1(n90), .B2(n93), .A(n91), .ZN(n89) );
  OAI21_X4 U95 ( .B1(n109), .B2(n95), .A(n96), .ZN(n94) );
  NAND2_X4 U96 ( .A1(n103), .A2(n97), .ZN(n95) );
  AOI21_X4 U97 ( .B1(n97), .B2(n104), .A(n98), .ZN(n96) );
  NOR2_X4 U98 ( .A1(n101), .A2(n99), .ZN(n97) );
  OAI21_X4 U99 ( .B1(n99), .B2(n102), .A(n100), .ZN(n98) );
  NOR2_X4 U104 ( .A1(n107), .A2(n105), .ZN(n103) );
  OAI21_X4 U105 ( .B1(n105), .B2(n108), .A(n106), .ZN(n104) );
  AOI21_X4 U110 ( .B1(n110), .B2(n116), .A(n111), .ZN(n109) );
  NOR2_X4 U111 ( .A1(n114), .A2(n112), .ZN(n110) );
  OAI21_X4 U112 ( .B1(n112), .B2(n115), .A(n113), .ZN(n111) );
  NOR2_X4 U113 ( .A1(n123), .A2(B[3]), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n123), .A2(B[3]), .ZN(n113) );
  NOR2_X4 U115 ( .A1(n122), .A2(B[2]), .ZN(n114) );
  NAND2_X4 U116 ( .A1(n122), .A2(B[2]), .ZN(n115) );
  OAI21_X4 U117 ( .B1(n117), .B2(n119), .A(n118), .ZN(n116) );
  NOR2_X4 U118 ( .A1(n121), .A2(B[1]), .ZN(n117) );
  NAND2_X4 U119 ( .A1(n121), .A2(B[1]), .ZN(n118) );
  NAND2_X4 U120 ( .A1(n120), .A2(B[0]), .ZN(n119) );
  INV_X1 U157 ( .A(A[14]), .ZN(n134) );
  INV_X2 U158 ( .A(A[18]), .ZN(n138) );
  INV_X1 U159 ( .A(A[12]), .ZN(n132) );
  OAI21_X1 U160 ( .B1(n1), .B2(n6), .A(n7), .ZN(GE_LT_GT_LE) );
  INV_X1 U161 ( .A(A[28]), .ZN(n148) );
  INV_X1 U162 ( .A(A[27]), .ZN(n147) );
  INV_X1 U163 ( .A(A[24]), .ZN(n144) );
  INV_X4 U164 ( .A(A[1]), .ZN(n121) );
  INV_X4 U165 ( .A(A[0]), .ZN(n120) );
  OAI21_X2 U166 ( .B1(n32), .B2(n35), .A(n33), .ZN(n31) );
  NOR2_X1 U167 ( .A1(n34), .A2(n32), .ZN(n30) );
  INV_X4 U168 ( .A(A[25]), .ZN(n145) );
  INV_X4 U169 ( .A(A[2]), .ZN(n122) );
  AOI21_X2 U170 ( .B1(n12), .B2(n19), .A(n13), .ZN(n11) );
  INV_X4 U171 ( .A(A[30]), .ZN(n150) );
  OAI21_X1 U172 ( .B1(n51), .B2(n36), .A(n37), .ZN(n2) );
  INV_X4 U173 ( .A(A[22]), .ZN(n142) );
  INV_X1 U174 ( .A(A[10]), .ZN(n130) );
  INV_X1 U175 ( .A(A[6]), .ZN(n126) );
  INV_X2 U176 ( .A(A[13]), .ZN(n133) );
  INV_X1 U177 ( .A(A[8]), .ZN(n128) );
  INV_X1 U178 ( .A(A[4]), .ZN(n124) );
  NAND2_X1 U179 ( .A1(n124), .A2(B[4]), .ZN(n108) );
  NOR2_X1 U180 ( .A1(n124), .A2(B[4]), .ZN(n107) );
  INV_X1 U181 ( .A(A[7]), .ZN(n127) );
  INV_X1 U182 ( .A(A[19]), .ZN(n139) );
  INV_X1 U183 ( .A(A[29]), .ZN(n149) );
  INV_X4 U184 ( .A(A[21]), .ZN(n141) );
  OAI21_X1 U185 ( .B1(n14), .B2(n17), .A(n15), .ZN(n13) );
  INV_X1 U186 ( .A(B[31]), .ZN(n151) );
  NAND2_X1 U187 ( .A1(n151), .A2(A[31]), .ZN(n15) );
  NOR2_X1 U188 ( .A1(n151), .A2(A[31]), .ZN(n14) );
  INV_X2 U189 ( .A(A[17]), .ZN(n137) );
  INV_X1 U190 ( .A(A[5]), .ZN(n125) );
  NAND2_X1 U191 ( .A1(n133), .A2(B[13]), .ZN(n77) );
  NOR2_X1 U192 ( .A1(n133), .A2(B[13]), .ZN(n76) );
  NAND2_X1 U193 ( .A1(n129), .A2(B[9]), .ZN(n91) );
  NOR2_X1 U194 ( .A1(n129), .A2(B[9]), .ZN(n90) );
  NAND2_X1 U195 ( .A1(n127), .A2(B[7]), .ZN(n100) );
  NOR2_X1 U196 ( .A1(n127), .A2(B[7]), .ZN(n99) );
  NAND2_X1 U197 ( .A1(n135), .A2(B[15]), .ZN(n71) );
  NOR2_X1 U198 ( .A1(n135), .A2(B[15]), .ZN(n70) );
  NAND2_X1 U199 ( .A1(n137), .A2(B[17]), .ZN(n61) );
  NOR2_X1 U200 ( .A1(n137), .A2(B[17]), .ZN(n60) );
  NOR2_X1 U201 ( .A1(n136), .A2(B[16]), .ZN(n62) );
  NAND2_X1 U202 ( .A1(n136), .A2(B[16]), .ZN(n63) );
  NAND2_X1 U203 ( .A1(n131), .A2(B[11]), .ZN(n85) );
  NOR2_X1 U204 ( .A1(n131), .A2(B[11]), .ZN(n84) );
  INV_X2 U205 ( .A(A[9]), .ZN(n129) );
  NOR2_X1 U206 ( .A1(n138), .A2(B[18]), .ZN(n56) );
  NAND2_X1 U207 ( .A1(n126), .A2(B[6]), .ZN(n102) );
  NOR2_X1 U208 ( .A1(n126), .A2(B[6]), .ZN(n101) );
  NAND2_X1 U209 ( .A1(n125), .A2(B[5]), .ZN(n106) );
  NOR2_X1 U210 ( .A1(n125), .A2(B[5]), .ZN(n105) );
  INV_X1 U211 ( .A(A[11]), .ZN(n131) );
  NAND2_X1 U212 ( .A1(n139), .A2(B[19]), .ZN(n55) );
  NOR2_X1 U213 ( .A1(n139), .A2(B[19]), .ZN(n54) );
  NOR2_X1 U214 ( .A1(n130), .A2(B[10]), .ZN(n86) );
  NAND2_X1 U215 ( .A1(n130), .A2(B[10]), .ZN(n87) );
  NOR2_X1 U216 ( .A1(n132), .A2(B[12]), .ZN(n78) );
  NAND2_X1 U217 ( .A1(n132), .A2(B[12]), .ZN(n79) );
  NAND2_X1 U218 ( .A1(n134), .A2(B[14]), .ZN(n73) );
  NOR2_X1 U219 ( .A1(n134), .A2(B[14]), .ZN(n72) );
  NOR2_X1 U220 ( .A1(n140), .A2(B[20]), .ZN(n48) );
  NAND2_X1 U221 ( .A1(n140), .A2(B[20]), .ZN(n49) );
  INV_X1 U222 ( .A(A[26]), .ZN(n146) );
  NAND2_X1 U223 ( .A1(n138), .A2(B[18]), .ZN(n57) );
  INV_X1 U224 ( .A(A[3]), .ZN(n123) );
  INV_X1 U225 ( .A(A[23]), .ZN(n143) );
  NOR2_X1 U226 ( .A1(n128), .A2(B[8]), .ZN(n92) );
  NAND2_X1 U227 ( .A1(n128), .A2(B[8]), .ZN(n93) );
  INV_X2 U228 ( .A(A[16]), .ZN(n136) );
  INV_X4 U229 ( .A(A[15]), .ZN(n135) );
  INV_X4 U230 ( .A(A[20]), .ZN(n140) );
endmodule


module Xi_core_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636;

  INV_X4 U107 ( .A(n1179), .ZN(n1174) );
  INV_X1 U108 ( .A(A[24]), .ZN(n1421) );
  NAND2_X1 U109 ( .A1(A[4]), .A2(n1177), .ZN(n1626) );
  INV_X1 U110 ( .A(A[27]), .ZN(n1370) );
  NAND2_X1 U111 ( .A1(A[1]), .A2(n1175), .ZN(n1534) );
  INV_X1 U112 ( .A(A[1]), .ZN(n1620) );
  NAND2_X1 U113 ( .A1(A[0]), .A2(n1178), .ZN(n1636) );
  INV_X1 U114 ( .A(A[25]), .ZN(n1404) );
  NAND2_X1 U115 ( .A1(A[2]), .A2(n1175), .ZN(n1520) );
  INV_X1 U116 ( .A(A[2]), .ZN(n1634) );
  INV_X1 U117 ( .A(A[22]), .ZN(n1455) );
  INV_X1 U118 ( .A(A[0]), .ZN(n1628) );
  INV_X1 U119 ( .A(A[4]), .ZN(n1594) );
  INV_X1 U120 ( .A(A[21]), .ZN(n1472) );
  NAND2_X1 U121 ( .A1(A[6]), .A2(n1178), .ZN(n1632) );
  INV_X1 U122 ( .A(A[6]), .ZN(n1571) );
  NAND2_X1 U123 ( .A1(A[7]), .A2(n1176), .ZN(n1614) );
  INV_X1 U124 ( .A(A[7]), .ZN(n1559) );
  NAND2_X1 U125 ( .A1(A[5]), .A2(n1177), .ZN(n1618) );
  INV_X1 U126 ( .A(A[5]), .ZN(n1583) );
  INV_X1 U127 ( .A(A[19]), .ZN(n1371) );
  INV_X1 U128 ( .A(A[18]), .ZN(n1388) );
  INV_X1 U129 ( .A(A[16]), .ZN(n1422) );
  INV_X1 U130 ( .A(A[13]), .ZN(n1473) );
  INV_X1 U131 ( .A(A[17]), .ZN(n1405) );
  INV_X1 U132 ( .A(A[15]), .ZN(n1439) );
  INV_X1 U133 ( .A(A[14]), .ZN(n1456) );
  INV_X1 U134 ( .A(A[20]), .ZN(n1489) );
  INV_X1 U135 ( .A(A[12]), .ZN(n1490) );
  INV_X1 U136 ( .A(A[9]), .ZN(n1531) );
  INV_X1 U137 ( .A(A[11]), .ZN(n1504) );
  INV_X1 U138 ( .A(A[8]), .ZN(n1545) );
  INV_X1 U139 ( .A(A[10]), .ZN(n1517) );
  INV_X1 U140 ( .A(n1172), .ZN(n1162) );
  INV_X1 U141 ( .A(n1172), .ZN(n1163) );
  INV_X1 U142 ( .A(n1172), .ZN(n1164) );
  INV_X1 U143 ( .A(n1172), .ZN(n1165) );
  INV_X1 U144 ( .A(n1171), .ZN(n1166) );
  CLKBUF_X3 U145 ( .A(SH[4]), .Z(n1167) );
  CLKBUF_X3 U146 ( .A(SH[4]), .Z(n1168) );
  CLKBUF_X3 U147 ( .A(SH[4]), .Z(n1169) );
  CLKBUF_X3 U148 ( .A(SH[4]), .Z(n1170) );
  CLKBUF_X3 U149 ( .A(SH[4]), .Z(n1171) );
  CLKBUF_X3 U150 ( .A(SH[4]), .Z(n1172) );
  INV_X1 U151 ( .A(n1179), .ZN(n1173) );
  INV_X1 U152 ( .A(SH[3]), .ZN(n1175) );
  INV_X1 U153 ( .A(SH[3]), .ZN(n1176) );
  INV_X1 U154 ( .A(SH[3]), .ZN(n1177) );
  INV_X1 U155 ( .A(SH[3]), .ZN(n1178) );
  INV_X1 U156 ( .A(SH[3]), .ZN(n1179) );
  INV_X1 U157 ( .A(n1183), .ZN(n1180) );
  INV_X1 U158 ( .A(n1183), .ZN(n1181) );
  INV_X1 U159 ( .A(n1183), .ZN(n1182) );
  INV_X8 U160 ( .A(SH[2]), .ZN(n1183) );
  INV_X1 U161 ( .A(n1189), .ZN(n1184) );
  INV_X1 U162 ( .A(n1188), .ZN(n1185) );
  INV_X1 U163 ( .A(n1189), .ZN(n1186) );
  INV_X1 U164 ( .A(n1188), .ZN(n1187) );
  INV_X2 U165 ( .A(SH[1]), .ZN(n1188) );
  INV_X2 U166 ( .A(SH[1]), .ZN(n1189) );
  INV_X1 U167 ( .A(n1196), .ZN(n1190) );
  INV_X1 U168 ( .A(n1199), .ZN(n1191) );
  INV_X1 U169 ( .A(n1200), .ZN(n1192) );
  INV_X1 U170 ( .A(n1201), .ZN(n1193) );
  INV_X1 U171 ( .A(n1202), .ZN(n1194) );
  CLKBUF_X3 U172 ( .A(SH[0]), .Z(n1195) );
  CLKBUF_X3 U173 ( .A(SH[0]), .Z(n1196) );
  CLKBUF_X3 U174 ( .A(SH[0]), .Z(n1197) );
  CLKBUF_X3 U175 ( .A(SH[0]), .Z(n1198) );
  CLKBUF_X3 U176 ( .A(SH[0]), .Z(n1199) );
  CLKBUF_X3 U177 ( .A(SH[0]), .Z(n1200) );
  CLKBUF_X3 U178 ( .A(SH[0]), .Z(n1201) );
  CLKBUF_X3 U179 ( .A(SH[0]), .Z(n1202) );
  CLKBUF_X3 U180 ( .A(SH[0]), .Z(n1203) );
  CLKBUF_X3 U181 ( .A(SH[0]), .Z(n1204) );
  CLKBUF_X3 U182 ( .A(SH[0]), .Z(n1205) );
  CLKBUF_X3 U183 ( .A(SH[0]), .Z(n1206) );
  CLKBUF_X3 U184 ( .A(SH[0]), .Z(n1207) );
  CLKBUF_X3 U185 ( .A(SH[0]), .Z(n1208) );
  CLKBUF_X3 U186 ( .A(SH[0]), .Z(n1209) );
  NAND2_X2 U187 ( .A1(n1210), .A2(n1211), .ZN(B[9]) );
  MUX2_X1 U188 ( .A(n1212), .B(n1213), .S(n1184), .Z(n1211) );
  NAND2_X2 U189 ( .A1(n1208), .A2(n1214), .ZN(n1213) );
  NAND2_X2 U190 ( .A1(n1209), .A2(n1215), .ZN(n1212) );
  MUX2_X1 U191 ( .A(n1216), .B(n1217), .S(n1187), .Z(n1210) );
  NAND2_X2 U192 ( .A1(n1218), .A2(n1192), .ZN(n1217) );
  NAND2_X2 U193 ( .A1(n1219), .A2(n1190), .ZN(n1216) );
  NAND2_X2 U194 ( .A1(n1220), .A2(n1221), .ZN(B[8]) );
  MUX2_X1 U195 ( .A(n1222), .B(n1223), .S(n1187), .Z(n1221) );
  NAND2_X2 U196 ( .A1(n1209), .A2(n1224), .ZN(n1223) );
  NAND2_X2 U197 ( .A1(n1208), .A2(n1218), .ZN(n1222) );
  MUX2_X1 U198 ( .A(n1225), .B(n1226), .S(n1187), .Z(n1220) );
  NAND2_X2 U199 ( .A1(n1214), .A2(n1190), .ZN(n1226) );
  NAND2_X2 U200 ( .A1(n1215), .A2(n1190), .ZN(n1225) );
  NAND2_X2 U201 ( .A1(n1227), .A2(n1228), .ZN(B[7]) );
  MUX2_X1 U202 ( .A(n1229), .B(n1230), .S(n1187), .Z(n1228) );
  NAND2_X2 U203 ( .A1(n1208), .A2(n1231), .ZN(n1230) );
  NAND2_X2 U204 ( .A1(n1207), .A2(n1214), .ZN(n1229) );
  MUX2_X1 U205 ( .A(n1232), .B(n1233), .S(n1187), .Z(n1227) );
  NAND2_X2 U206 ( .A1(n1224), .A2(n1190), .ZN(n1233) );
  NAND2_X2 U207 ( .A1(n1218), .A2(n1190), .ZN(n1232) );
  NAND2_X2 U208 ( .A1(n1234), .A2(n1235), .ZN(B[6]) );
  MUX2_X1 U209 ( .A(n1236), .B(n1237), .S(n1186), .Z(n1235) );
  NAND2_X2 U210 ( .A1(n1238), .A2(n1195), .ZN(n1237) );
  NAND2_X2 U211 ( .A1(n1208), .A2(n1224), .ZN(n1236) );
  MUX2_X1 U212 ( .A(n1239), .B(n1240), .S(n1186), .Z(n1234) );
  NAND2_X2 U213 ( .A1(n1231), .A2(n1190), .ZN(n1240) );
  NAND2_X2 U214 ( .A1(n1214), .A2(n1190), .ZN(n1239) );
  INV_X2 U215 ( .A(n1241), .ZN(n1214) );
  MUX2_X1 U216 ( .A(n1242), .B(n1243), .S(n1180), .Z(n1241) );
  NAND2_X2 U217 ( .A1(n1244), .A2(n1164), .ZN(n1243) );
  NAND2_X2 U218 ( .A1(n1245), .A2(n1162), .ZN(n1242) );
  NAND2_X2 U219 ( .A1(n1246), .A2(n1247), .ZN(B[5]) );
  MUX2_X1 U220 ( .A(n1248), .B(n1249), .S(n1186), .Z(n1247) );
  NAND2_X2 U221 ( .A1(n1250), .A2(n1195), .ZN(n1249) );
  NAND2_X2 U222 ( .A1(n1207), .A2(n1231), .ZN(n1248) );
  MUX2_X1 U223 ( .A(n1251), .B(n1252), .S(n1186), .Z(n1246) );
  NAND2_X2 U224 ( .A1(n1238), .A2(n1190), .ZN(n1252) );
  NAND2_X2 U225 ( .A1(n1224), .A2(n1190), .ZN(n1251) );
  INV_X2 U226 ( .A(n1253), .ZN(n1224) );
  MUX2_X1 U227 ( .A(n1254), .B(n1255), .S(n1182), .Z(n1253) );
  NAND2_X2 U228 ( .A1(n1256), .A2(n1162), .ZN(n1255) );
  NAND2_X2 U229 ( .A1(n1257), .A2(n1162), .ZN(n1254) );
  NAND2_X2 U230 ( .A1(n1258), .A2(n1259), .ZN(B[4]) );
  MUX2_X1 U231 ( .A(n1260), .B(n1261), .S(n1186), .Z(n1259) );
  NAND2_X2 U232 ( .A1(n1262), .A2(n1195), .ZN(n1261) );
  NAND2_X2 U233 ( .A1(n1238), .A2(n1196), .ZN(n1260) );
  MUX2_X1 U234 ( .A(n1263), .B(n1264), .S(n1186), .Z(n1258) );
  NAND2_X2 U235 ( .A1(n1250), .A2(n1190), .ZN(n1264) );
  NAND2_X2 U236 ( .A1(n1231), .A2(n1190), .ZN(n1263) );
  INV_X2 U237 ( .A(n1265), .ZN(n1231) );
  MUX2_X1 U238 ( .A(n1266), .B(n1267), .S(n1182), .Z(n1265) );
  NAND2_X2 U239 ( .A1(n1268), .A2(n1162), .ZN(n1267) );
  NAND2_X2 U240 ( .A1(n1269), .A2(n1162), .ZN(n1266) );
  NAND2_X2 U241 ( .A1(n1270), .A2(n1271), .ZN(B[3]) );
  MUX2_X1 U242 ( .A(n1272), .B(n1273), .S(n1186), .Z(n1271) );
  NAND2_X2 U243 ( .A1(n1274), .A2(n1196), .ZN(n1273) );
  NAND2_X2 U244 ( .A1(n1250), .A2(n1195), .ZN(n1272) );
  MUX2_X1 U245 ( .A(n1275), .B(n1276), .S(n1186), .Z(n1270) );
  NAND2_X2 U246 ( .A1(n1262), .A2(n1190), .ZN(n1276) );
  NAND2_X2 U247 ( .A1(n1238), .A2(n1191), .ZN(n1275) );
  INV_X2 U248 ( .A(n1277), .ZN(n1238) );
  NAND3_X1 U249 ( .A1(n1183), .A2(n1166), .A3(n1278), .ZN(n1277) );
  NAND2_X2 U250 ( .A1(n1279), .A2(n1280), .ZN(B[31]) );
  MUX2_X1 U251 ( .A(n1281), .B(n1282), .S(n1186), .Z(n1280) );
  NAND2_X2 U252 ( .A1(n1207), .A2(n1283), .ZN(n1282) );
  NAND2_X2 U253 ( .A1(n1207), .A2(n1284), .ZN(n1281) );
  MUX2_X1 U254 ( .A(n1285), .B(n1286), .S(n1186), .Z(n1279) );
  NAND2_X2 U255 ( .A1(n1287), .A2(n1191), .ZN(n1286) );
  OAI21_X2 U256 ( .B1(n1288), .B2(n1289), .A(n1194), .ZN(n1285) );
  MUX2_X1 U257 ( .A(n1290), .B(n1291), .S(n1182), .Z(n1289) );
  AND2_X2 U258 ( .A1(n1292), .A2(n1165), .ZN(n1291) );
  AND2_X2 U259 ( .A1(n1293), .A2(n1165), .ZN(n1290) );
  MUX2_X1 U260 ( .A(A[31]), .B(A[23]), .S(n1173), .Z(n1293) );
  MUX2_X1 U261 ( .A(n1294), .B(n1295), .S(n1182), .Z(n1288) );
  AND2_X2 U262 ( .A1(n1172), .A2(n1296), .ZN(n1295) );
  AND2_X2 U263 ( .A1(n1172), .A2(n1297), .ZN(n1294) );
  NAND2_X2 U264 ( .A1(n1298), .A2(n1299), .ZN(B[30]) );
  MUX2_X1 U265 ( .A(n1300), .B(n1301), .S(n1186), .Z(n1299) );
  NAND2_X2 U266 ( .A1(n1206), .A2(n1302), .ZN(n1301) );
  NAND2_X2 U267 ( .A1(n1206), .A2(n1287), .ZN(n1300) );
  MUX2_X1 U268 ( .A(n1303), .B(n1304), .S(n1186), .Z(n1298) );
  NAND2_X2 U269 ( .A1(n1283), .A2(n1191), .ZN(n1304) );
  NAND2_X2 U270 ( .A1(n1284), .A2(n1191), .ZN(n1303) );
  NAND2_X2 U271 ( .A1(n1305), .A2(n1306), .ZN(n1284) );
  MUX2_X1 U272 ( .A(n1307), .B(n1308), .S(n1182), .Z(n1306) );
  NAND2_X2 U273 ( .A1(n1171), .A2(n1309), .ZN(n1308) );
  NAND2_X2 U274 ( .A1(n1171), .A2(n1310), .ZN(n1307) );
  MUX2_X1 U275 ( .A(n1311), .B(n1312), .S(n1182), .Z(n1305) );
  NAND2_X2 U276 ( .A1(n1313), .A2(n1162), .ZN(n1312) );
  NAND2_X2 U277 ( .A1(n1314), .A2(n1162), .ZN(n1311) );
  MUX2_X1 U278 ( .A(A[30]), .B(A[22]), .S(n1173), .Z(n1314) );
  NAND2_X2 U279 ( .A1(n1315), .A2(n1316), .ZN(B[2]) );
  NAND3_X1 U280 ( .A1(n1194), .A2(n1189), .A3(n1250), .ZN(n1316) );
  INV_X2 U281 ( .A(n1317), .ZN(n1250) );
  NAND3_X1 U282 ( .A1(n1183), .A2(n1166), .A3(n1244), .ZN(n1317) );
  MUX2_X1 U283 ( .A(n1318), .B(n1319), .S(n1197), .Z(n1315) );
  NAND2_X2 U284 ( .A1(n1262), .A2(n1188), .ZN(n1319) );
  NAND2_X2 U285 ( .A1(n1274), .A2(n1184), .ZN(n1318) );
  NAND2_X2 U286 ( .A1(n1320), .A2(n1321), .ZN(B[29]) );
  MUX2_X1 U287 ( .A(n1322), .B(n1323), .S(n1186), .Z(n1321) );
  NAND2_X2 U288 ( .A1(n1206), .A2(n1324), .ZN(n1323) );
  NAND2_X2 U289 ( .A1(n1206), .A2(n1283), .ZN(n1322) );
  MUX2_X1 U290 ( .A(n1325), .B(n1326), .S(n1186), .Z(n1320) );
  NAND2_X2 U291 ( .A1(n1302), .A2(n1191), .ZN(n1326) );
  NAND2_X2 U292 ( .A1(n1287), .A2(n1191), .ZN(n1325) );
  NAND2_X2 U293 ( .A1(n1327), .A2(n1328), .ZN(n1287) );
  MUX2_X1 U294 ( .A(n1329), .B(n1330), .S(n1182), .Z(n1328) );
  NAND2_X2 U295 ( .A1(n1170), .A2(n1331), .ZN(n1330) );
  NAND2_X2 U296 ( .A1(n1170), .A2(n1332), .ZN(n1329) );
  MUX2_X1 U297 ( .A(n1333), .B(n1334), .S(n1182), .Z(n1327) );
  NAND2_X2 U298 ( .A1(n1335), .A2(n1162), .ZN(n1334) );
  NAND2_X2 U299 ( .A1(n1336), .A2(n1162), .ZN(n1333) );
  MUX2_X1 U300 ( .A(A[29]), .B(A[21]), .S(n1173), .Z(n1336) );
  NAND2_X2 U301 ( .A1(n1337), .A2(n1338), .ZN(B[28]) );
  MUX2_X1 U302 ( .A(n1339), .B(n1340), .S(n1186), .Z(n1338) );
  NAND2_X2 U303 ( .A1(n1205), .A2(n1341), .ZN(n1340) );
  NAND2_X2 U304 ( .A1(n1205), .A2(n1302), .ZN(n1339) );
  MUX2_X1 U305 ( .A(n1342), .B(n1343), .S(n1186), .Z(n1337) );
  NAND2_X2 U306 ( .A1(n1324), .A2(n1191), .ZN(n1343) );
  NAND2_X2 U307 ( .A1(n1283), .A2(n1191), .ZN(n1342) );
  NAND2_X2 U308 ( .A1(n1344), .A2(n1345), .ZN(n1283) );
  MUX2_X1 U309 ( .A(n1346), .B(n1347), .S(n1181), .Z(n1345) );
  NAND2_X2 U310 ( .A1(n1170), .A2(n1348), .ZN(n1347) );
  NAND2_X2 U311 ( .A1(n1170), .A2(n1349), .ZN(n1346) );
  MUX2_X1 U312 ( .A(n1350), .B(n1351), .S(n1181), .Z(n1344) );
  NAND2_X2 U313 ( .A1(n1352), .A2(n1162), .ZN(n1351) );
  NAND2_X2 U314 ( .A1(n1353), .A2(n1162), .ZN(n1350) );
  MUX2_X1 U315 ( .A(A[28]), .B(A[20]), .S(n1173), .Z(n1353) );
  NAND2_X2 U316 ( .A1(n1354), .A2(n1355), .ZN(B[27]) );
  MUX2_X1 U317 ( .A(n1356), .B(n1357), .S(n1186), .Z(n1355) );
  NAND2_X2 U318 ( .A1(n1205), .A2(n1358), .ZN(n1357) );
  NAND2_X2 U319 ( .A1(n1205), .A2(n1324), .ZN(n1356) );
  MUX2_X1 U320 ( .A(n1359), .B(n1360), .S(n1186), .Z(n1354) );
  NAND2_X2 U321 ( .A1(n1341), .A2(n1191), .ZN(n1360) );
  NAND2_X2 U322 ( .A1(n1302), .A2(n1191), .ZN(n1359) );
  NAND2_X2 U323 ( .A1(n1361), .A2(n1362), .ZN(n1302) );
  MUX2_X1 U324 ( .A(n1363), .B(n1364), .S(n1181), .Z(n1362) );
  NAND2_X2 U325 ( .A1(n1170), .A2(n1365), .ZN(n1364) );
  NAND2_X2 U326 ( .A1(n1169), .A2(n1296), .ZN(n1363) );
  MUX2_X1 U327 ( .A(n1366), .B(n1367), .S(n1181), .Z(n1361) );
  NAND2_X2 U328 ( .A1(n1368), .A2(n1162), .ZN(n1367) );
  NAND2_X2 U329 ( .A1(n1292), .A2(n1163), .ZN(n1366) );
  INV_X2 U330 ( .A(n1369), .ZN(n1292) );
  MUX2_X1 U331 ( .A(n1370), .B(n1371), .S(n1173), .Z(n1369) );
  NAND2_X2 U332 ( .A1(n1372), .A2(n1373), .ZN(B[26]) );
  MUX2_X1 U333 ( .A(n1374), .B(n1375), .S(n1185), .Z(n1373) );
  NAND2_X2 U334 ( .A1(n1204), .A2(n1376), .ZN(n1375) );
  NAND2_X2 U335 ( .A1(n1204), .A2(n1341), .ZN(n1374) );
  MUX2_X1 U336 ( .A(n1377), .B(n1378), .S(n1185), .Z(n1372) );
  NAND2_X2 U337 ( .A1(n1358), .A2(n1191), .ZN(n1378) );
  NAND2_X2 U338 ( .A1(n1324), .A2(n1191), .ZN(n1377) );
  NAND2_X2 U339 ( .A1(n1379), .A2(n1380), .ZN(n1324) );
  MUX2_X1 U340 ( .A(n1381), .B(n1382), .S(n1181), .Z(n1380) );
  NAND2_X2 U341 ( .A1(n1169), .A2(n1245), .ZN(n1382) );
  NAND2_X2 U342 ( .A1(n1169), .A2(n1309), .ZN(n1381) );
  MUX2_X1 U343 ( .A(n1383), .B(n1384), .S(n1181), .Z(n1379) );
  NAND2_X2 U344 ( .A1(n1385), .A2(n1163), .ZN(n1384) );
  NAND2_X2 U345 ( .A1(n1313), .A2(n1163), .ZN(n1383) );
  INV_X2 U346 ( .A(n1386), .ZN(n1313) );
  MUX2_X1 U347 ( .A(n1387), .B(n1388), .S(n1173), .Z(n1386) );
  INV_X2 U348 ( .A(A[26]), .ZN(n1387) );
  NAND2_X2 U349 ( .A1(n1389), .A2(n1390), .ZN(B[25]) );
  MUX2_X1 U350 ( .A(n1391), .B(n1392), .S(n1185), .Z(n1390) );
  NAND2_X2 U351 ( .A1(n1204), .A2(n1393), .ZN(n1392) );
  NAND2_X2 U352 ( .A1(n1204), .A2(n1358), .ZN(n1391) );
  MUX2_X1 U353 ( .A(n1394), .B(n1395), .S(n1185), .Z(n1389) );
  NAND2_X2 U354 ( .A1(n1376), .A2(n1192), .ZN(n1395) );
  NAND2_X2 U355 ( .A1(n1341), .A2(n1192), .ZN(n1394) );
  NAND2_X2 U356 ( .A1(n1396), .A2(n1397), .ZN(n1341) );
  MUX2_X1 U357 ( .A(n1398), .B(n1399), .S(n1181), .Z(n1397) );
  NAND2_X2 U358 ( .A1(n1169), .A2(n1257), .ZN(n1399) );
  NAND2_X2 U359 ( .A1(n1169), .A2(n1331), .ZN(n1398) );
  MUX2_X1 U360 ( .A(n1400), .B(n1401), .S(n1181), .Z(n1396) );
  NAND2_X2 U361 ( .A1(n1402), .A2(n1163), .ZN(n1401) );
  NAND2_X2 U362 ( .A1(n1335), .A2(n1163), .ZN(n1400) );
  INV_X2 U363 ( .A(n1403), .ZN(n1335) );
  MUX2_X1 U364 ( .A(n1404), .B(n1405), .S(n1173), .Z(n1403) );
  NAND2_X2 U365 ( .A1(n1406), .A2(n1407), .ZN(B[24]) );
  MUX2_X1 U366 ( .A(n1408), .B(n1409), .S(n1185), .Z(n1407) );
  NAND2_X2 U367 ( .A1(n1203), .A2(n1410), .ZN(n1409) );
  NAND2_X2 U368 ( .A1(n1203), .A2(n1376), .ZN(n1408) );
  MUX2_X1 U369 ( .A(n1411), .B(n1412), .S(n1185), .Z(n1406) );
  NAND2_X2 U370 ( .A1(n1393), .A2(n1192), .ZN(n1412) );
  NAND2_X2 U371 ( .A1(n1358), .A2(n1192), .ZN(n1411) );
  NAND2_X2 U372 ( .A1(n1413), .A2(n1414), .ZN(n1358) );
  MUX2_X1 U373 ( .A(n1415), .B(n1416), .S(n1181), .Z(n1414) );
  NAND2_X2 U374 ( .A1(n1168), .A2(n1269), .ZN(n1416) );
  NAND2_X2 U375 ( .A1(n1168), .A2(n1348), .ZN(n1415) );
  MUX2_X1 U376 ( .A(n1417), .B(n1418), .S(n1181), .Z(n1413) );
  NAND2_X2 U377 ( .A1(n1419), .A2(n1163), .ZN(n1418) );
  NAND2_X2 U378 ( .A1(n1352), .A2(n1163), .ZN(n1417) );
  INV_X2 U379 ( .A(n1420), .ZN(n1352) );
  MUX2_X1 U380 ( .A(n1421), .B(n1422), .S(n1173), .Z(n1420) );
  NAND2_X2 U381 ( .A1(n1423), .A2(n1424), .ZN(B[23]) );
  MUX2_X1 U382 ( .A(n1425), .B(n1426), .S(n1185), .Z(n1424) );
  NAND2_X2 U383 ( .A1(n1203), .A2(n1427), .ZN(n1426) );
  NAND2_X2 U384 ( .A1(n1202), .A2(n1393), .ZN(n1425) );
  MUX2_X1 U385 ( .A(n1428), .B(n1429), .S(n1185), .Z(n1423) );
  NAND2_X2 U386 ( .A1(n1410), .A2(n1192), .ZN(n1429) );
  NAND2_X2 U387 ( .A1(n1376), .A2(n1192), .ZN(n1428) );
  NAND2_X2 U388 ( .A1(n1430), .A2(n1431), .ZN(n1376) );
  MUX2_X1 U389 ( .A(n1432), .B(n1433), .S(n1181), .Z(n1431) );
  NAND2_X2 U390 ( .A1(n1168), .A2(n1278), .ZN(n1433) );
  NAND2_X2 U391 ( .A1(n1168), .A2(n1365), .ZN(n1432) );
  MUX2_X1 U392 ( .A(n1434), .B(n1435), .S(n1181), .Z(n1430) );
  NAND2_X2 U393 ( .A1(n1436), .A2(n1163), .ZN(n1435) );
  NAND2_X2 U394 ( .A1(n1368), .A2(n1163), .ZN(n1434) );
  INV_X2 U395 ( .A(n1437), .ZN(n1368) );
  MUX2_X1 U396 ( .A(n1438), .B(n1439), .S(n1173), .Z(n1437) );
  INV_X2 U397 ( .A(A[23]), .ZN(n1438) );
  NAND2_X2 U398 ( .A1(n1440), .A2(n1441), .ZN(B[22]) );
  MUX2_X1 U399 ( .A(n1442), .B(n1443), .S(n1185), .Z(n1441) );
  NAND2_X2 U400 ( .A1(n1202), .A2(n1444), .ZN(n1443) );
  NAND2_X2 U401 ( .A1(n1202), .A2(n1410), .ZN(n1442) );
  MUX2_X1 U402 ( .A(n1445), .B(n1446), .S(n1185), .Z(n1440) );
  NAND2_X2 U403 ( .A1(n1427), .A2(n1192), .ZN(n1446) );
  NAND2_X2 U404 ( .A1(n1393), .A2(n1192), .ZN(n1445) );
  NAND2_X2 U405 ( .A1(n1447), .A2(n1448), .ZN(n1393) );
  MUX2_X1 U406 ( .A(n1449), .B(n1450), .S(n1181), .Z(n1448) );
  NAND2_X2 U407 ( .A1(n1168), .A2(n1244), .ZN(n1450) );
  NAND2_X2 U408 ( .A1(n1167), .A2(n1245), .ZN(n1449) );
  MUX2_X1 U409 ( .A(n1451), .B(n1452), .S(n1181), .Z(n1447) );
  NAND2_X2 U410 ( .A1(n1453), .A2(n1163), .ZN(n1452) );
  NAND2_X2 U411 ( .A1(n1385), .A2(n1163), .ZN(n1451) );
  INV_X2 U412 ( .A(n1454), .ZN(n1385) );
  MUX2_X1 U413 ( .A(n1455), .B(n1456), .S(n1173), .Z(n1454) );
  NAND2_X2 U414 ( .A1(n1457), .A2(n1458), .ZN(B[21]) );
  MUX2_X1 U415 ( .A(n1459), .B(n1460), .S(n1185), .Z(n1458) );
  NAND2_X2 U416 ( .A1(n1202), .A2(n1461), .ZN(n1460) );
  NAND2_X2 U417 ( .A1(n1201), .A2(n1427), .ZN(n1459) );
  MUX2_X1 U418 ( .A(n1462), .B(n1463), .S(n1185), .Z(n1457) );
  NAND2_X2 U419 ( .A1(n1444), .A2(n1192), .ZN(n1463) );
  NAND2_X2 U420 ( .A1(n1410), .A2(n1192), .ZN(n1462) );
  NAND2_X2 U421 ( .A1(n1464), .A2(n1465), .ZN(n1410) );
  MUX2_X1 U422 ( .A(n1466), .B(n1467), .S(n1181), .Z(n1465) );
  NAND2_X2 U423 ( .A1(n1167), .A2(n1256), .ZN(n1467) );
  NAND2_X2 U424 ( .A1(n1167), .A2(n1257), .ZN(n1466) );
  MUX2_X1 U425 ( .A(n1468), .B(n1469), .S(n1181), .Z(n1464) );
  NAND2_X2 U426 ( .A1(n1470), .A2(n1163), .ZN(n1469) );
  NAND2_X2 U427 ( .A1(n1402), .A2(n1164), .ZN(n1468) );
  INV_X2 U428 ( .A(n1471), .ZN(n1402) );
  MUX2_X1 U429 ( .A(n1472), .B(n1473), .S(n1173), .Z(n1471) );
  NAND2_X2 U430 ( .A1(n1474), .A2(n1475), .ZN(B[20]) );
  MUX2_X1 U431 ( .A(n1476), .B(n1477), .S(n1185), .Z(n1475) );
  NAND2_X2 U432 ( .A1(n1201), .A2(n1478), .ZN(n1477) );
  NAND2_X2 U433 ( .A1(n1201), .A2(n1444), .ZN(n1476) );
  MUX2_X1 U434 ( .A(n1479), .B(n1480), .S(n1185), .Z(n1474) );
  NAND2_X2 U435 ( .A1(n1461), .A2(n1192), .ZN(n1480) );
  NAND2_X2 U436 ( .A1(n1427), .A2(n1193), .ZN(n1479) );
  NAND2_X2 U437 ( .A1(n1481), .A2(n1482), .ZN(n1427) );
  MUX2_X1 U438 ( .A(n1483), .B(n1484), .S(n1180), .Z(n1482) );
  NAND2_X2 U439 ( .A1(n1167), .A2(n1268), .ZN(n1484) );
  NAND2_X2 U440 ( .A1(n1167), .A2(n1269), .ZN(n1483) );
  MUX2_X1 U441 ( .A(n1485), .B(n1486), .S(n1180), .Z(n1481) );
  NAND2_X2 U442 ( .A1(n1487), .A2(n1164), .ZN(n1486) );
  NAND2_X2 U443 ( .A1(n1419), .A2(n1164), .ZN(n1485) );
  INV_X2 U444 ( .A(n1488), .ZN(n1419) );
  MUX2_X1 U445 ( .A(n1489), .B(n1490), .S(n1173), .Z(n1488) );
  MUX2_X1 U446 ( .A(n1491), .B(n1492), .S(n1198), .Z(B[1]) );
  AND2_X2 U447 ( .A1(n1274), .A2(n1188), .ZN(n1492) );
  AND2_X2 U448 ( .A1(n1262), .A2(n1188), .ZN(n1491) );
  INV_X2 U449 ( .A(n1493), .ZN(n1262) );
  NAND3_X1 U450 ( .A1(n1183), .A2(n1165), .A3(n1256), .ZN(n1493) );
  NAND2_X2 U451 ( .A1(n1494), .A2(n1495), .ZN(B[19]) );
  MUX2_X1 U452 ( .A(n1496), .B(n1497), .S(n1185), .Z(n1495) );
  NAND2_X2 U453 ( .A1(n1201), .A2(n1498), .ZN(n1497) );
  NAND2_X2 U454 ( .A1(n1200), .A2(n1461), .ZN(n1496) );
  MUX2_X1 U455 ( .A(n1499), .B(n1500), .S(n1185), .Z(n1494) );
  NAND2_X2 U456 ( .A1(n1478), .A2(n1193), .ZN(n1500) );
  NAND2_X2 U457 ( .A1(n1444), .A2(n1193), .ZN(n1499) );
  NAND2_X2 U458 ( .A1(n1501), .A2(n1502), .ZN(n1444) );
  NAND3_X1 U459 ( .A1(n1183), .A2(n1166), .A3(n1436), .ZN(n1502) );
  INV_X2 U460 ( .A(n1503), .ZN(n1436) );
  MUX2_X1 U461 ( .A(n1371), .B(n1504), .S(n1174), .Z(n1503) );
  MUX2_X1 U462 ( .A(n1505), .B(n1506), .S(n1171), .Z(n1501) );
  NAND2_X2 U463 ( .A1(n1278), .A2(n1183), .ZN(n1506) );
  NAND2_X2 U464 ( .A1(n1180), .A2(n1297), .ZN(n1505) );
  NAND2_X2 U465 ( .A1(n1507), .A2(n1508), .ZN(B[18]) );
  MUX2_X1 U466 ( .A(n1509), .B(n1510), .S(n1185), .Z(n1508) );
  NAND2_X2 U467 ( .A1(n1200), .A2(n1511), .ZN(n1510) );
  NAND2_X2 U468 ( .A1(n1200), .A2(n1478), .ZN(n1509) );
  MUX2_X1 U469 ( .A(n1512), .B(n1513), .S(n1184), .Z(n1507) );
  NAND2_X2 U470 ( .A1(n1498), .A2(n1193), .ZN(n1513) );
  NAND2_X2 U471 ( .A1(n1461), .A2(n1193), .ZN(n1512) );
  NAND2_X2 U472 ( .A1(n1514), .A2(n1515), .ZN(n1461) );
  NAND3_X1 U473 ( .A1(n1183), .A2(n1166), .A3(n1453), .ZN(n1515) );
  INV_X2 U474 ( .A(n1516), .ZN(n1453) );
  MUX2_X1 U475 ( .A(n1388), .B(n1517), .S(n1174), .Z(n1516) );
  MUX2_X1 U476 ( .A(n1518), .B(n1519), .S(n1171), .Z(n1514) );
  NAND2_X2 U477 ( .A1(n1244), .A2(n1183), .ZN(n1519) );
  INV_X2 U478 ( .A(n1520), .ZN(n1244) );
  NAND2_X2 U479 ( .A1(n1180), .A2(n1310), .ZN(n1518) );
  NAND2_X2 U480 ( .A1(n1521), .A2(n1522), .ZN(B[17]) );
  MUX2_X1 U481 ( .A(n1523), .B(n1524), .S(n1184), .Z(n1522) );
  NAND2_X2 U482 ( .A1(n1200), .A2(n1525), .ZN(n1524) );
  NAND2_X2 U483 ( .A1(n1199), .A2(n1498), .ZN(n1523) );
  MUX2_X1 U484 ( .A(n1526), .B(n1527), .S(n1184), .Z(n1521) );
  NAND2_X2 U485 ( .A1(n1511), .A2(n1193), .ZN(n1527) );
  NAND2_X2 U486 ( .A1(n1478), .A2(n1193), .ZN(n1526) );
  NAND2_X2 U487 ( .A1(n1528), .A2(n1529), .ZN(n1478) );
  NAND3_X1 U488 ( .A1(n1183), .A2(n1166), .A3(n1470), .ZN(n1529) );
  INV_X2 U489 ( .A(n1530), .ZN(n1470) );
  MUX2_X1 U490 ( .A(n1405), .B(n1531), .S(n1174), .Z(n1530) );
  MUX2_X1 U491 ( .A(n1532), .B(n1533), .S(n1171), .Z(n1528) );
  NAND2_X2 U492 ( .A1(n1256), .A2(n1183), .ZN(n1533) );
  INV_X2 U493 ( .A(n1534), .ZN(n1256) );
  NAND2_X2 U494 ( .A1(n1180), .A2(n1332), .ZN(n1532) );
  NAND2_X2 U495 ( .A1(n1535), .A2(n1536), .ZN(B[16]) );
  MUX2_X1 U496 ( .A(n1537), .B(n1538), .S(n1184), .Z(n1536) );
  NAND2_X2 U497 ( .A1(n1198), .A2(n1539), .ZN(n1538) );
  NAND2_X2 U498 ( .A1(n1198), .A2(n1511), .ZN(n1537) );
  MUX2_X1 U499 ( .A(n1540), .B(n1541), .S(n1184), .Z(n1535) );
  NAND2_X2 U500 ( .A1(n1525), .A2(n1193), .ZN(n1541) );
  NAND2_X2 U501 ( .A1(n1498), .A2(n1193), .ZN(n1540) );
  NAND2_X2 U502 ( .A1(n1542), .A2(n1543), .ZN(n1498) );
  NAND3_X1 U503 ( .A1(n1183), .A2(n1166), .A3(n1487), .ZN(n1543) );
  INV_X2 U504 ( .A(n1544), .ZN(n1487) );
  MUX2_X1 U505 ( .A(n1422), .B(n1545), .S(n1174), .Z(n1544) );
  MUX2_X1 U506 ( .A(n1546), .B(n1547), .S(n1171), .Z(n1542) );
  NAND2_X2 U507 ( .A1(n1268), .A2(n1183), .ZN(n1547) );
  NAND2_X2 U508 ( .A1(n1180), .A2(n1349), .ZN(n1546) );
  NAND2_X2 U509 ( .A1(n1548), .A2(n1549), .ZN(B[15]) );
  MUX2_X1 U510 ( .A(n1550), .B(n1551), .S(n1184), .Z(n1549) );
  NAND2_X2 U511 ( .A1(n1197), .A2(n1552), .ZN(n1551) );
  NAND2_X2 U512 ( .A1(n1199), .A2(n1525), .ZN(n1550) );
  MUX2_X1 U513 ( .A(n1553), .B(n1554), .S(n1184), .Z(n1548) );
  NAND2_X2 U514 ( .A1(n1539), .A2(n1193), .ZN(n1554) );
  NAND2_X2 U515 ( .A1(n1511), .A2(n1193), .ZN(n1553) );
  INV_X2 U516 ( .A(n1555), .ZN(n1511) );
  MUX2_X1 U517 ( .A(n1556), .B(n1557), .S(n1180), .Z(n1555) );
  NAND2_X2 U518 ( .A1(n1296), .A2(n1164), .ZN(n1557) );
  NAND2_X2 U519 ( .A1(n1297), .A2(n1164), .ZN(n1556) );
  INV_X2 U520 ( .A(n1558), .ZN(n1297) );
  MUX2_X1 U521 ( .A(n1439), .B(n1559), .S(n1174), .Z(n1558) );
  NAND2_X2 U522 ( .A1(n1560), .A2(n1561), .ZN(B[14]) );
  MUX2_X1 U523 ( .A(n1562), .B(n1563), .S(n1184), .Z(n1561) );
  NAND2_X2 U524 ( .A1(n1197), .A2(n1564), .ZN(n1563) );
  NAND2_X2 U525 ( .A1(n1199), .A2(n1539), .ZN(n1562) );
  MUX2_X1 U526 ( .A(n1565), .B(n1566), .S(n1184), .Z(n1560) );
  NAND2_X2 U527 ( .A1(n1552), .A2(n1194), .ZN(n1566) );
  NAND2_X2 U528 ( .A1(n1525), .A2(n1194), .ZN(n1565) );
  INV_X2 U529 ( .A(n1567), .ZN(n1525) );
  MUX2_X1 U530 ( .A(n1568), .B(n1569), .S(n1180), .Z(n1567) );
  NAND2_X2 U531 ( .A1(n1309), .A2(n1164), .ZN(n1569) );
  NAND2_X2 U532 ( .A1(n1310), .A2(n1164), .ZN(n1568) );
  INV_X2 U533 ( .A(n1570), .ZN(n1310) );
  MUX2_X1 U534 ( .A(n1456), .B(n1571), .S(n1174), .Z(n1570) );
  NAND2_X2 U535 ( .A1(n1572), .A2(n1573), .ZN(B[13]) );
  MUX2_X1 U536 ( .A(n1574), .B(n1575), .S(n1184), .Z(n1573) );
  NAND2_X2 U537 ( .A1(n1197), .A2(n1576), .ZN(n1575) );
  NAND2_X2 U538 ( .A1(n1198), .A2(n1552), .ZN(n1574) );
  MUX2_X1 U539 ( .A(n1577), .B(n1578), .S(n1184), .Z(n1572) );
  NAND2_X2 U540 ( .A1(n1564), .A2(n1194), .ZN(n1578) );
  NAND2_X2 U541 ( .A1(n1539), .A2(n1194), .ZN(n1577) );
  INV_X2 U542 ( .A(n1579), .ZN(n1539) );
  MUX2_X1 U543 ( .A(n1580), .B(n1581), .S(n1180), .Z(n1579) );
  NAND2_X2 U544 ( .A1(n1331), .A2(n1164), .ZN(n1581) );
  NAND2_X2 U545 ( .A1(n1332), .A2(n1165), .ZN(n1580) );
  INV_X2 U546 ( .A(n1582), .ZN(n1332) );
  MUX2_X1 U547 ( .A(n1473), .B(n1583), .S(n1174), .Z(n1582) );
  NAND2_X2 U548 ( .A1(n1584), .A2(n1585), .ZN(B[12]) );
  MUX2_X1 U549 ( .A(n1586), .B(n1587), .S(n1184), .Z(n1585) );
  NAND2_X2 U550 ( .A1(n1197), .A2(n1219), .ZN(n1587) );
  NAND2_X2 U551 ( .A1(n1199), .A2(n1564), .ZN(n1586) );
  MUX2_X1 U552 ( .A(n1588), .B(n1589), .S(n1184), .Z(n1584) );
  NAND2_X2 U553 ( .A1(n1576), .A2(n1193), .ZN(n1589) );
  NAND2_X2 U554 ( .A1(n1552), .A2(n1194), .ZN(n1588) );
  INV_X2 U555 ( .A(n1590), .ZN(n1552) );
  MUX2_X1 U556 ( .A(n1591), .B(n1592), .S(n1180), .Z(n1590) );
  NAND2_X2 U557 ( .A1(n1348), .A2(n1164), .ZN(n1592) );
  NAND2_X2 U558 ( .A1(n1349), .A2(n1164), .ZN(n1591) );
  INV_X2 U559 ( .A(n1593), .ZN(n1349) );
  MUX2_X1 U560 ( .A(n1490), .B(n1594), .S(n1174), .Z(n1593) );
  NAND2_X2 U561 ( .A1(n1595), .A2(n1596), .ZN(B[11]) );
  MUX2_X1 U562 ( .A(n1597), .B(n1598), .S(n1184), .Z(n1596) );
  NAND2_X2 U563 ( .A1(n1196), .A2(n1215), .ZN(n1598) );
  NAND2_X2 U564 ( .A1(n1198), .A2(n1576), .ZN(n1597) );
  MUX2_X1 U565 ( .A(n1599), .B(n1600), .S(n1184), .Z(n1595) );
  NAND2_X2 U566 ( .A1(n1219), .A2(n1194), .ZN(n1600) );
  NAND2_X2 U567 ( .A1(n1564), .A2(n1194), .ZN(n1599) );
  INV_X2 U568 ( .A(n1601), .ZN(n1564) );
  MUX2_X1 U569 ( .A(n1602), .B(n1603), .S(n1180), .Z(n1601) );
  NAND2_X2 U570 ( .A1(n1365), .A2(n1165), .ZN(n1603) );
  NAND2_X2 U571 ( .A1(n1296), .A2(n1164), .ZN(n1602) );
  INV_X2 U572 ( .A(n1604), .ZN(n1296) );
  MUX2_X1 U573 ( .A(n1504), .B(n1605), .S(n1174), .Z(n1604) );
  INV_X2 U574 ( .A(A[3]), .ZN(n1605) );
  NAND2_X2 U575 ( .A1(n1606), .A2(n1607), .ZN(B[10]) );
  MUX2_X1 U576 ( .A(n1608), .B(n1609), .S(n1184), .Z(n1607) );
  NAND2_X2 U577 ( .A1(n1196), .A2(n1218), .ZN(n1609) );
  INV_X2 U578 ( .A(n1610), .ZN(n1218) );
  MUX2_X1 U579 ( .A(n1611), .B(n1612), .S(n1180), .Z(n1610) );
  NAND2_X2 U580 ( .A1(n1278), .A2(n1165), .ZN(n1612) );
  INV_X2 U581 ( .A(n1613), .ZN(n1278) );
  NAND2_X2 U582 ( .A1(A[3]), .A2(n1176), .ZN(n1613) );
  NAND2_X2 U583 ( .A1(n1365), .A2(n1165), .ZN(n1611) );
  INV_X2 U584 ( .A(n1614), .ZN(n1365) );
  NAND2_X2 U585 ( .A1(n1203), .A2(n1219), .ZN(n1608) );
  INV_X2 U586 ( .A(n1615), .ZN(n1219) );
  MUX2_X1 U587 ( .A(n1616), .B(n1617), .S(n1180), .Z(n1615) );
  NAND2_X2 U588 ( .A1(n1257), .A2(n1165), .ZN(n1617) );
  INV_X2 U589 ( .A(n1618), .ZN(n1257) );
  NAND2_X2 U590 ( .A1(n1331), .A2(n1165), .ZN(n1616) );
  INV_X2 U591 ( .A(n1619), .ZN(n1331) );
  MUX2_X1 U592 ( .A(n1531), .B(n1620), .S(n1174), .Z(n1619) );
  MUX2_X1 U593 ( .A(n1621), .B(n1622), .S(n1185), .Z(n1606) );
  NAND2_X2 U594 ( .A1(n1215), .A2(n1194), .ZN(n1622) );
  INV_X2 U595 ( .A(n1623), .ZN(n1215) );
  MUX2_X1 U596 ( .A(n1624), .B(n1625), .S(n1180), .Z(n1623) );
  NAND2_X2 U597 ( .A1(n1269), .A2(n1165), .ZN(n1625) );
  INV_X2 U598 ( .A(n1626), .ZN(n1269) );
  NAND2_X2 U599 ( .A1(n1348), .A2(n1165), .ZN(n1624) );
  INV_X2 U600 ( .A(n1627), .ZN(n1348) );
  MUX2_X1 U601 ( .A(n1545), .B(n1628), .S(n1174), .Z(n1627) );
  NAND2_X2 U602 ( .A1(n1576), .A2(n1194), .ZN(n1621) );
  INV_X2 U603 ( .A(n1629), .ZN(n1576) );
  MUX2_X1 U604 ( .A(n1630), .B(n1631), .S(n1181), .Z(n1629) );
  NAND2_X2 U605 ( .A1(n1245), .A2(n1165), .ZN(n1631) );
  INV_X2 U606 ( .A(n1632), .ZN(n1245) );
  NAND2_X2 U607 ( .A1(n1309), .A2(n1165), .ZN(n1630) );
  INV_X2 U608 ( .A(n1633), .ZN(n1309) );
  MUX2_X1 U609 ( .A(n1517), .B(n1634), .S(n1174), .Z(n1633) );
  AND3_X2 U610 ( .A1(n1194), .A2(n1189), .A3(n1274), .ZN(B[0]) );
  INV_X2 U611 ( .A(n1635), .ZN(n1274) );
  NAND3_X1 U612 ( .A1(n1183), .A2(n1166), .A3(n1268), .ZN(n1635) );
  INV_X2 U613 ( .A(n1636), .ZN(n1268) );
endmodule


module Xi_core_DW01_bsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671;

  INV_X1 U169 ( .A(A[24]), .ZN(n1595) );
  INV_X1 U170 ( .A(A[26]), .ZN(n1461) );
  INV_X1 U171 ( .A(A[28]), .ZN(n1591) );
  INV_X1 U172 ( .A(A[27]), .ZN(n1573) );
  INV_X1 U173 ( .A(A[1]), .ZN(n1479) );
  INV_X1 U174 ( .A(A[25]), .ZN(n1480) );
  INV_X1 U175 ( .A(A[30]), .ZN(n1623) );
  INV_X1 U176 ( .A(A[0]), .ZN(n1599) );
  INV_X1 U177 ( .A(A[2]), .ZN(n1460) );
  INV_X1 U178 ( .A(A[29]), .ZN(n1611) );
  INV_X1 U179 ( .A(A[4]), .ZN(n1590) );
  INV_X1 U180 ( .A(A[22]), .ZN(n1619) );
  INV_X1 U181 ( .A(A[21]), .ZN(n1607) );
  INV_X1 U182 ( .A(A[31]), .ZN(n1581) );
  INV_X1 U183 ( .A(A[6]), .ZN(n1622) );
  INV_X1 U184 ( .A(A[7]), .ZN(n1580) );
  INV_X1 U185 ( .A(A[5]), .ZN(n1610) );
  INV_X1 U186 ( .A(A[19]), .ZN(n1569) );
  INV_X1 U187 ( .A(A[18]), .ZN(n1463) );
  INV_X1 U188 ( .A(A[16]), .ZN(n1596) );
  INV_X1 U189 ( .A(A[13]), .ZN(n1608) );
  INV_X1 U190 ( .A(A[17]), .ZN(n1482) );
  INV_X1 U191 ( .A(A[15]), .ZN(n1578) );
  INV_X1 U192 ( .A(A[14]), .ZN(n1620) );
  INV_X1 U193 ( .A(A[20]), .ZN(n1587) );
  INV_X1 U194 ( .A(A[12]), .ZN(n1588) );
  INV_X1 U195 ( .A(A[9]), .ZN(n1483) );
  INV_X1 U196 ( .A(A[11]), .ZN(n1570) );
  INV_X1 U197 ( .A(A[8]), .ZN(n1598) );
  INV_X1 U198 ( .A(A[10]), .ZN(n1464) );
  CLKBUF_X3 U199 ( .A(SH[4]), .Z(n1105) );
  CLKBUF_X3 U200 ( .A(SH[4]), .Z(n1106) );
  CLKBUF_X3 U201 ( .A(SH[4]), .Z(n1107) );
  CLKBUF_X3 U202 ( .A(SH[4]), .Z(n1108) );
  CLKBUF_X3 U203 ( .A(SH[4]), .Z(n1109) );
  CLKBUF_X3 U204 ( .A(SH[4]), .Z(n1110) );
  CLKBUF_X3 U205 ( .A(SH[3]), .Z(n1111) );
  CLKBUF_X3 U206 ( .A(SH[3]), .Z(n1112) );
  CLKBUF_X3 U207 ( .A(SH[3]), .Z(n1113) );
  INV_X1 U208 ( .A(n1132), .ZN(n1114) );
  INV_X1 U209 ( .A(n1132), .ZN(n1115) );
  INV_X1 U210 ( .A(n1133), .ZN(n1116) );
  INV_X1 U211 ( .A(n1133), .ZN(n1117) );
  INV_X1 U212 ( .A(n1133), .ZN(n1118) );
  INV_X1 U213 ( .A(n1133), .ZN(n1119) );
  CLKBUF_X3 U214 ( .A(SH[2]), .Z(n1120) );
  CLKBUF_X3 U215 ( .A(SH[2]), .Z(n1121) );
  CLKBUF_X3 U216 ( .A(SH[2]), .Z(n1122) );
  CLKBUF_X3 U217 ( .A(SH[2]), .Z(n1123) );
  CLKBUF_X3 U218 ( .A(SH[2]), .Z(n1124) );
  CLKBUF_X3 U219 ( .A(SH[2]), .Z(n1125) );
  CLKBUF_X3 U220 ( .A(SH[2]), .Z(n1126) );
  CLKBUF_X3 U221 ( .A(SH[2]), .Z(n1127) );
  CLKBUF_X3 U222 ( .A(SH[2]), .Z(n1128) );
  CLKBUF_X3 U223 ( .A(SH[2]), .Z(n1129) );
  CLKBUF_X3 U224 ( .A(SH[2]), .Z(n1130) );
  CLKBUF_X3 U225 ( .A(SH[2]), .Z(n1131) );
  CLKBUF_X3 U226 ( .A(SH[2]), .Z(n1132) );
  CLKBUF_X3 U227 ( .A(SH[2]), .Z(n1133) );
  INV_X1 U228 ( .A(n1152), .ZN(n1134) );
  INV_X1 U229 ( .A(n1152), .ZN(n1135) );
  INV_X1 U230 ( .A(n1153), .ZN(n1136) );
  INV_X1 U231 ( .A(n1153), .ZN(n1137) );
  INV_X1 U232 ( .A(n1153), .ZN(n1138) );
  INV_X1 U233 ( .A(n1153), .ZN(n1139) );
  CLKBUF_X3 U234 ( .A(SH[1]), .Z(n1140) );
  CLKBUF_X3 U235 ( .A(SH[1]), .Z(n1141) );
  CLKBUF_X3 U236 ( .A(SH[1]), .Z(n1142) );
  CLKBUF_X3 U237 ( .A(SH[1]), .Z(n1143) );
  CLKBUF_X3 U238 ( .A(SH[1]), .Z(n1144) );
  CLKBUF_X3 U239 ( .A(SH[1]), .Z(n1145) );
  CLKBUF_X3 U240 ( .A(SH[1]), .Z(n1146) );
  CLKBUF_X3 U241 ( .A(SH[1]), .Z(n1147) );
  CLKBUF_X3 U242 ( .A(SH[1]), .Z(n1148) );
  CLKBUF_X3 U243 ( .A(SH[1]), .Z(n1149) );
  CLKBUF_X3 U244 ( .A(SH[1]), .Z(n1150) );
  CLKBUF_X3 U245 ( .A(SH[1]), .Z(n1151) );
  CLKBUF_X3 U246 ( .A(SH[1]), .Z(n1152) );
  CLKBUF_X3 U247 ( .A(SH[1]), .Z(n1153) );
  CLKBUF_X3 U248 ( .A(SH[0]), .Z(n1154) );
  CLKBUF_X3 U249 ( .A(SH[0]), .Z(n1155) );
  CLKBUF_X3 U250 ( .A(SH[0]), .Z(n1156) );
  CLKBUF_X3 U251 ( .A(SH[0]), .Z(n1157) );
  CLKBUF_X3 U252 ( .A(SH[0]), .Z(n1158) );
  CLKBUF_X3 U253 ( .A(SH[0]), .Z(n1159) );
  NAND2_X2 U254 ( .A1(n1160), .A2(n1161), .ZN(B[9]) );
  MUX2_X1 U255 ( .A(n1162), .B(n1163), .S(n1154), .Z(n1161) );
  NAND2_X2 U256 ( .A1(n1152), .A2(n1164), .ZN(n1163) );
  NAND2_X2 U257 ( .A1(n1152), .A2(n1165), .ZN(n1162) );
  MUX2_X1 U258 ( .A(n1166), .B(n1167), .S(n1154), .Z(n1160) );
  NAND2_X2 U259 ( .A1(n1168), .A2(n1139), .ZN(n1167) );
  NAND2_X2 U260 ( .A1(n1169), .A2(n1139), .ZN(n1166) );
  NAND2_X2 U261 ( .A1(n1170), .A2(n1171), .ZN(B[8]) );
  MUX2_X1 U262 ( .A(n1172), .B(n1173), .S(n1154), .Z(n1171) );
  NAND2_X2 U263 ( .A1(n1152), .A2(n1174), .ZN(n1173) );
  NAND2_X2 U264 ( .A1(n1152), .A2(n1164), .ZN(n1172) );
  MUX2_X1 U265 ( .A(n1175), .B(n1176), .S(n1154), .Z(n1170) );
  NAND2_X2 U266 ( .A1(n1165), .A2(n1139), .ZN(n1176) );
  NAND2_X2 U267 ( .A1(n1168), .A2(n1139), .ZN(n1175) );
  NAND2_X2 U268 ( .A1(n1177), .A2(n1178), .ZN(B[7]) );
  MUX2_X1 U269 ( .A(n1179), .B(n1180), .S(n1154), .Z(n1178) );
  NAND2_X2 U270 ( .A1(n1151), .A2(n1181), .ZN(n1180) );
  NAND2_X2 U271 ( .A1(n1151), .A2(n1174), .ZN(n1179) );
  MUX2_X1 U272 ( .A(n1182), .B(n1183), .S(n1154), .Z(n1177) );
  NAND2_X2 U273 ( .A1(n1164), .A2(n1138), .ZN(n1183) );
  NAND2_X2 U274 ( .A1(n1165), .A2(n1138), .ZN(n1182) );
  NAND2_X2 U275 ( .A1(n1184), .A2(n1185), .ZN(B[6]) );
  MUX2_X1 U276 ( .A(n1186), .B(n1187), .S(n1154), .Z(n1185) );
  NAND2_X2 U277 ( .A1(n1151), .A2(n1188), .ZN(n1187) );
  NAND2_X2 U278 ( .A1(n1151), .A2(n1181), .ZN(n1186) );
  MUX2_X1 U279 ( .A(n1189), .B(n1190), .S(n1154), .Z(n1184) );
  NAND2_X2 U280 ( .A1(n1174), .A2(n1138), .ZN(n1190) );
  NAND2_X2 U281 ( .A1(n1164), .A2(n1138), .ZN(n1189) );
  NAND2_X2 U282 ( .A1(n1191), .A2(n1192), .ZN(n1164) );
  MUX2_X1 U283 ( .A(n1193), .B(n1194), .S(n1105), .Z(n1192) );
  NAND2_X2 U284 ( .A1(n1132), .A2(n1195), .ZN(n1194) );
  NAND2_X2 U285 ( .A1(n1132), .A2(n1196), .ZN(n1193) );
  MUX2_X1 U286 ( .A(n1197), .B(n1198), .S(n1105), .Z(n1191) );
  NAND2_X2 U287 ( .A1(n1199), .A2(n1119), .ZN(n1198) );
  NAND2_X2 U288 ( .A1(n1200), .A2(n1119), .ZN(n1197) );
  NAND2_X2 U289 ( .A1(n1201), .A2(n1202), .ZN(B[5]) );
  MUX2_X1 U290 ( .A(n1203), .B(n1204), .S(n1154), .Z(n1202) );
  NAND2_X2 U291 ( .A1(n1151), .A2(n1205), .ZN(n1204) );
  NAND2_X2 U292 ( .A1(n1150), .A2(n1188), .ZN(n1203) );
  MUX2_X1 U293 ( .A(n1206), .B(n1207), .S(n1154), .Z(n1201) );
  NAND2_X2 U294 ( .A1(n1181), .A2(n1138), .ZN(n1207) );
  NAND2_X2 U295 ( .A1(n1174), .A2(n1138), .ZN(n1206) );
  NAND2_X2 U296 ( .A1(n1208), .A2(n1209), .ZN(n1174) );
  MUX2_X1 U297 ( .A(n1210), .B(n1211), .S(n1105), .Z(n1209) );
  NAND2_X2 U298 ( .A1(n1132), .A2(n1212), .ZN(n1211) );
  NAND2_X2 U299 ( .A1(n1132), .A2(n1213), .ZN(n1210) );
  MUX2_X1 U300 ( .A(n1214), .B(n1215), .S(n1105), .Z(n1208) );
  NAND2_X2 U301 ( .A1(n1216), .A2(n1119), .ZN(n1215) );
  NAND2_X2 U302 ( .A1(n1217), .A2(n1119), .ZN(n1214) );
  NAND2_X2 U303 ( .A1(n1218), .A2(n1219), .ZN(B[4]) );
  MUX2_X1 U304 ( .A(n1220), .B(n1221), .S(n1154), .Z(n1219) );
  NAND2_X2 U305 ( .A1(n1150), .A2(n1222), .ZN(n1221) );
  NAND2_X2 U306 ( .A1(n1150), .A2(n1205), .ZN(n1220) );
  MUX2_X1 U307 ( .A(n1223), .B(n1224), .S(n1154), .Z(n1218) );
  NAND2_X2 U308 ( .A1(n1188), .A2(n1138), .ZN(n1224) );
  NAND2_X2 U309 ( .A1(n1181), .A2(n1138), .ZN(n1223) );
  NAND2_X2 U310 ( .A1(n1225), .A2(n1226), .ZN(n1181) );
  MUX2_X1 U311 ( .A(n1227), .B(n1228), .S(n1105), .Z(n1226) );
  NAND2_X2 U312 ( .A1(n1131), .A2(n1229), .ZN(n1228) );
  NAND2_X2 U313 ( .A1(n1131), .A2(n1230), .ZN(n1227) );
  MUX2_X1 U314 ( .A(n1231), .B(n1232), .S(n1105), .Z(n1225) );
  NAND2_X2 U315 ( .A1(n1233), .A2(n1118), .ZN(n1232) );
  NAND2_X2 U316 ( .A1(n1234), .A2(n1118), .ZN(n1231) );
  NAND2_X2 U317 ( .A1(n1235), .A2(n1236), .ZN(B[3]) );
  MUX2_X1 U318 ( .A(n1237), .B(n1238), .S(n1155), .Z(n1236) );
  NAND2_X2 U319 ( .A1(n1150), .A2(n1239), .ZN(n1238) );
  NAND2_X2 U320 ( .A1(n1150), .A2(n1222), .ZN(n1237) );
  MUX2_X1 U321 ( .A(n1240), .B(n1241), .S(n1155), .Z(n1235) );
  NAND2_X2 U322 ( .A1(n1205), .A2(n1138), .ZN(n1241) );
  NAND2_X2 U323 ( .A1(n1188), .A2(n1138), .ZN(n1240) );
  NAND2_X2 U324 ( .A1(n1242), .A2(n1243), .ZN(n1188) );
  MUX2_X1 U325 ( .A(n1244), .B(n1245), .S(n1105), .Z(n1243) );
  NAND2_X2 U326 ( .A1(n1131), .A2(n1246), .ZN(n1245) );
  NAND2_X2 U327 ( .A1(n1131), .A2(n1247), .ZN(n1244) );
  MUX2_X1 U328 ( .A(n1248), .B(n1249), .S(n1105), .Z(n1242) );
  NAND2_X2 U329 ( .A1(n1250), .A2(n1118), .ZN(n1249) );
  NAND2_X2 U330 ( .A1(n1251), .A2(n1118), .ZN(n1248) );
  NAND2_X2 U331 ( .A1(n1252), .A2(n1253), .ZN(B[31]) );
  MUX2_X1 U332 ( .A(n1254), .B(n1255), .S(n1155), .Z(n1253) );
  NAND2_X2 U333 ( .A1(n1149), .A2(n1256), .ZN(n1255) );
  NAND2_X2 U334 ( .A1(n1149), .A2(n1257), .ZN(n1254) );
  MUX2_X1 U335 ( .A(n1258), .B(n1259), .S(n1155), .Z(n1252) );
  NAND2_X2 U336 ( .A1(n1260), .A2(n1138), .ZN(n1259) );
  NAND2_X2 U337 ( .A1(n1261), .A2(n1138), .ZN(n1258) );
  NAND2_X2 U338 ( .A1(n1262), .A2(n1263), .ZN(B[30]) );
  MUX2_X1 U339 ( .A(n1264), .B(n1265), .S(n1155), .Z(n1263) );
  NAND2_X2 U340 ( .A1(n1149), .A2(n1266), .ZN(n1265) );
  NAND2_X2 U341 ( .A1(n1149), .A2(n1256), .ZN(n1264) );
  MUX2_X1 U342 ( .A(n1267), .B(n1268), .S(n1155), .Z(n1262) );
  NAND2_X2 U343 ( .A1(n1257), .A2(n1137), .ZN(n1268) );
  NAND2_X2 U344 ( .A1(n1260), .A2(n1137), .ZN(n1267) );
  NAND2_X2 U345 ( .A1(n1269), .A2(n1270), .ZN(B[2]) );
  MUX2_X1 U346 ( .A(n1271), .B(n1272), .S(n1155), .Z(n1270) );
  NAND2_X2 U347 ( .A1(n1149), .A2(n1261), .ZN(n1272) );
  NAND2_X2 U348 ( .A1(n1148), .A2(n1239), .ZN(n1271) );
  MUX2_X1 U349 ( .A(n1273), .B(n1274), .S(n1155), .Z(n1269) );
  NAND2_X2 U350 ( .A1(n1222), .A2(n1137), .ZN(n1274) );
  NAND2_X2 U351 ( .A1(n1205), .A2(n1137), .ZN(n1273) );
  NAND2_X2 U352 ( .A1(n1275), .A2(n1276), .ZN(n1205) );
  MUX2_X1 U353 ( .A(n1277), .B(n1278), .S(n1105), .Z(n1276) );
  NAND2_X2 U354 ( .A1(n1131), .A2(n1279), .ZN(n1278) );
  NAND2_X2 U355 ( .A1(n1130), .A2(n1280), .ZN(n1277) );
  MUX2_X1 U356 ( .A(n1281), .B(n1282), .S(n1105), .Z(n1275) );
  NAND2_X2 U357 ( .A1(n1195), .A2(n1118), .ZN(n1282) );
  NAND2_X2 U358 ( .A1(n1196), .A2(n1118), .ZN(n1281) );
  NAND2_X2 U359 ( .A1(n1283), .A2(n1284), .ZN(B[29]) );
  MUX2_X1 U360 ( .A(n1285), .B(n1286), .S(n1155), .Z(n1284) );
  NAND2_X2 U361 ( .A1(n1148), .A2(n1287), .ZN(n1286) );
  NAND2_X2 U362 ( .A1(n1148), .A2(n1266), .ZN(n1285) );
  MUX2_X1 U363 ( .A(n1288), .B(n1289), .S(n1155), .Z(n1283) );
  NAND2_X2 U364 ( .A1(n1256), .A2(n1137), .ZN(n1289) );
  NAND2_X2 U365 ( .A1(n1257), .A2(n1137), .ZN(n1288) );
  NAND2_X2 U366 ( .A1(n1290), .A2(n1291), .ZN(B[28]) );
  MUX2_X1 U367 ( .A(n1292), .B(n1293), .S(n1155), .Z(n1291) );
  NAND2_X2 U368 ( .A1(n1148), .A2(n1294), .ZN(n1293) );
  NAND2_X2 U369 ( .A1(n1148), .A2(n1287), .ZN(n1292) );
  MUX2_X1 U370 ( .A(n1295), .B(n1296), .S(n1155), .Z(n1290) );
  NAND2_X2 U371 ( .A1(n1266), .A2(n1137), .ZN(n1296) );
  NAND2_X2 U372 ( .A1(n1256), .A2(n1137), .ZN(n1295) );
  NAND2_X2 U373 ( .A1(n1297), .A2(n1298), .ZN(n1256) );
  MUX2_X1 U374 ( .A(n1299), .B(n1300), .S(n1105), .Z(n1298) );
  NAND2_X2 U375 ( .A1(n1130), .A2(n1301), .ZN(n1300) );
  NAND2_X2 U376 ( .A1(n1130), .A2(n1302), .ZN(n1299) );
  MUX2_X1 U377 ( .A(n1303), .B(n1304), .S(n1105), .Z(n1297) );
  NAND2_X2 U378 ( .A1(n1305), .A2(n1118), .ZN(n1304) );
  NAND2_X2 U379 ( .A1(n1306), .A2(n1118), .ZN(n1303) );
  NAND2_X2 U380 ( .A1(n1307), .A2(n1308), .ZN(B[27]) );
  MUX2_X1 U381 ( .A(n1309), .B(n1310), .S(n1156), .Z(n1308) );
  NAND2_X2 U382 ( .A1(n1147), .A2(n1311), .ZN(n1310) );
  NAND2_X2 U383 ( .A1(n1147), .A2(n1294), .ZN(n1309) );
  MUX2_X1 U384 ( .A(n1312), .B(n1313), .S(n1156), .Z(n1307) );
  NAND2_X2 U385 ( .A1(n1287), .A2(n1137), .ZN(n1313) );
  NAND2_X2 U386 ( .A1(n1266), .A2(n1137), .ZN(n1312) );
  NAND2_X2 U387 ( .A1(n1314), .A2(n1315), .ZN(n1266) );
  MUX2_X1 U388 ( .A(n1316), .B(n1317), .S(n1106), .Z(n1315) );
  NAND2_X2 U389 ( .A1(n1130), .A2(n1318), .ZN(n1317) );
  NAND2_X2 U390 ( .A1(n1130), .A2(n1319), .ZN(n1316) );
  MUX2_X1 U391 ( .A(n1320), .B(n1321), .S(n1106), .Z(n1314) );
  NAND2_X2 U392 ( .A1(n1322), .A2(n1118), .ZN(n1321) );
  NAND2_X2 U393 ( .A1(n1323), .A2(n1118), .ZN(n1320) );
  NAND2_X2 U394 ( .A1(n1324), .A2(n1325), .ZN(B[26]) );
  MUX2_X1 U395 ( .A(n1326), .B(n1327), .S(n1156), .Z(n1325) );
  NAND2_X2 U396 ( .A1(n1147), .A2(n1328), .ZN(n1327) );
  NAND2_X2 U397 ( .A1(n1147), .A2(n1311), .ZN(n1326) );
  MUX2_X1 U398 ( .A(n1329), .B(n1330), .S(n1156), .Z(n1324) );
  NAND2_X2 U399 ( .A1(n1294), .A2(n1137), .ZN(n1330) );
  NAND2_X2 U400 ( .A1(n1287), .A2(n1137), .ZN(n1329) );
  NAND2_X2 U401 ( .A1(n1331), .A2(n1332), .ZN(n1287) );
  MUX2_X1 U402 ( .A(n1333), .B(n1334), .S(n1106), .Z(n1332) );
  NAND2_X2 U403 ( .A1(n1129), .A2(n1200), .ZN(n1334) );
  NAND2_X2 U404 ( .A1(n1129), .A2(n1199), .ZN(n1333) );
  MUX2_X1 U405 ( .A(n1335), .B(n1336), .S(n1106), .Z(n1331) );
  NAND2_X2 U406 ( .A1(n1337), .A2(n1118), .ZN(n1336) );
  NAND2_X2 U407 ( .A1(n1338), .A2(n1118), .ZN(n1335) );
  NAND2_X2 U408 ( .A1(n1339), .A2(n1340), .ZN(B[25]) );
  MUX2_X1 U409 ( .A(n1341), .B(n1342), .S(n1156), .Z(n1340) );
  NAND2_X2 U410 ( .A1(n1147), .A2(n1343), .ZN(n1342) );
  NAND2_X2 U411 ( .A1(n1146), .A2(n1328), .ZN(n1341) );
  MUX2_X1 U412 ( .A(n1344), .B(n1345), .S(n1156), .Z(n1339) );
  NAND2_X2 U413 ( .A1(n1311), .A2(n1136), .ZN(n1345) );
  NAND2_X2 U414 ( .A1(n1294), .A2(n1136), .ZN(n1344) );
  NAND2_X2 U415 ( .A1(n1346), .A2(n1347), .ZN(n1294) );
  MUX2_X1 U416 ( .A(n1348), .B(n1349), .S(n1106), .Z(n1347) );
  NAND2_X2 U417 ( .A1(n1129), .A2(n1217), .ZN(n1349) );
  NAND2_X2 U418 ( .A1(n1129), .A2(n1216), .ZN(n1348) );
  MUX2_X1 U419 ( .A(n1350), .B(n1351), .S(n1106), .Z(n1346) );
  NAND2_X2 U420 ( .A1(n1352), .A2(n1117), .ZN(n1351) );
  NAND2_X2 U421 ( .A1(n1353), .A2(n1117), .ZN(n1350) );
  NAND2_X2 U422 ( .A1(n1354), .A2(n1355), .ZN(B[24]) );
  MUX2_X1 U423 ( .A(n1356), .B(n1357), .S(n1156), .Z(n1355) );
  NAND2_X2 U424 ( .A1(n1146), .A2(n1358), .ZN(n1357) );
  NAND2_X2 U425 ( .A1(n1146), .A2(n1343), .ZN(n1356) );
  MUX2_X1 U426 ( .A(n1359), .B(n1360), .S(n1156), .Z(n1354) );
  NAND2_X2 U427 ( .A1(n1328), .A2(n1136), .ZN(n1360) );
  NAND2_X2 U428 ( .A1(n1311), .A2(n1136), .ZN(n1359) );
  NAND2_X2 U429 ( .A1(n1361), .A2(n1362), .ZN(n1311) );
  MUX2_X1 U430 ( .A(n1363), .B(n1364), .S(n1106), .Z(n1362) );
  NAND2_X2 U431 ( .A1(n1129), .A2(n1234), .ZN(n1364) );
  NAND2_X2 U432 ( .A1(n1128), .A2(n1233), .ZN(n1363) );
  MUX2_X1 U433 ( .A(n1365), .B(n1366), .S(n1106), .Z(n1361) );
  NAND2_X2 U434 ( .A1(n1301), .A2(n1117), .ZN(n1366) );
  NAND2_X2 U435 ( .A1(n1302), .A2(n1117), .ZN(n1365) );
  NAND2_X2 U436 ( .A1(n1367), .A2(n1368), .ZN(B[23]) );
  MUX2_X1 U437 ( .A(n1369), .B(n1370), .S(n1156), .Z(n1368) );
  NAND2_X2 U438 ( .A1(n1146), .A2(n1371), .ZN(n1370) );
  NAND2_X2 U439 ( .A1(n1146), .A2(n1358), .ZN(n1369) );
  MUX2_X1 U440 ( .A(n1372), .B(n1373), .S(n1156), .Z(n1367) );
  NAND2_X2 U441 ( .A1(n1343), .A2(n1136), .ZN(n1373) );
  NAND2_X2 U442 ( .A1(n1328), .A2(n1136), .ZN(n1372) );
  NAND2_X2 U443 ( .A1(n1374), .A2(n1375), .ZN(n1328) );
  MUX2_X1 U444 ( .A(n1376), .B(n1377), .S(n1106), .Z(n1375) );
  NAND2_X2 U445 ( .A1(n1128), .A2(n1251), .ZN(n1377) );
  NAND2_X2 U446 ( .A1(n1128), .A2(n1250), .ZN(n1376) );
  MUX2_X1 U447 ( .A(n1378), .B(n1379), .S(n1106), .Z(n1374) );
  NAND2_X2 U448 ( .A1(n1318), .A2(n1117), .ZN(n1379) );
  NAND2_X2 U449 ( .A1(n1319), .A2(n1117), .ZN(n1378) );
  NAND2_X2 U450 ( .A1(n1380), .A2(n1381), .ZN(B[22]) );
  MUX2_X1 U451 ( .A(n1382), .B(n1383), .S(n1156), .Z(n1381) );
  NAND2_X2 U452 ( .A1(n1145), .A2(n1384), .ZN(n1383) );
  NAND2_X2 U453 ( .A1(n1145), .A2(n1371), .ZN(n1382) );
  MUX2_X1 U454 ( .A(n1385), .B(n1386), .S(n1156), .Z(n1380) );
  NAND2_X2 U455 ( .A1(n1358), .A2(n1136), .ZN(n1386) );
  NAND2_X2 U456 ( .A1(n1343), .A2(n1136), .ZN(n1385) );
  NAND2_X2 U457 ( .A1(n1387), .A2(n1388), .ZN(n1343) );
  MUX2_X1 U458 ( .A(n1389), .B(n1390), .S(n1106), .Z(n1388) );
  NAND2_X2 U459 ( .A1(n1128), .A2(n1196), .ZN(n1390) );
  NAND2_X2 U460 ( .A1(n1128), .A2(n1195), .ZN(n1389) );
  MUX2_X1 U461 ( .A(n1391), .B(n1392), .S(n1106), .Z(n1387) );
  NAND2_X2 U462 ( .A1(n1200), .A2(n1117), .ZN(n1392) );
  NAND2_X2 U463 ( .A1(n1199), .A2(n1117), .ZN(n1391) );
  NAND2_X2 U464 ( .A1(n1393), .A2(n1394), .ZN(B[21]) );
  MUX2_X1 U465 ( .A(n1395), .B(n1396), .S(n1157), .Z(n1394) );
  NAND2_X2 U466 ( .A1(n1145), .A2(n1397), .ZN(n1396) );
  NAND2_X2 U467 ( .A1(n1145), .A2(n1384), .ZN(n1395) );
  MUX2_X1 U468 ( .A(n1398), .B(n1399), .S(n1157), .Z(n1393) );
  NAND2_X2 U469 ( .A1(n1371), .A2(n1136), .ZN(n1399) );
  NAND2_X2 U470 ( .A1(n1358), .A2(n1136), .ZN(n1398) );
  NAND2_X2 U471 ( .A1(n1400), .A2(n1401), .ZN(n1358) );
  MUX2_X1 U472 ( .A(n1402), .B(n1403), .S(n1107), .Z(n1401) );
  NAND2_X2 U473 ( .A1(n1127), .A2(n1213), .ZN(n1403) );
  NAND2_X2 U474 ( .A1(n1127), .A2(n1212), .ZN(n1402) );
  MUX2_X1 U475 ( .A(n1404), .B(n1405), .S(n1107), .Z(n1400) );
  NAND2_X2 U476 ( .A1(n1217), .A2(n1117), .ZN(n1405) );
  NAND2_X2 U477 ( .A1(n1216), .A2(n1117), .ZN(n1404) );
  NAND2_X2 U478 ( .A1(n1406), .A2(n1407), .ZN(B[20]) );
  MUX2_X1 U479 ( .A(n1408), .B(n1409), .S(n1157), .Z(n1407) );
  NAND2_X2 U480 ( .A1(n1145), .A2(n1410), .ZN(n1409) );
  NAND2_X2 U481 ( .A1(n1144), .A2(n1397), .ZN(n1408) );
  MUX2_X1 U482 ( .A(n1411), .B(n1412), .S(n1157), .Z(n1406) );
  NAND2_X2 U483 ( .A1(n1384), .A2(n1136), .ZN(n1412) );
  NAND2_X2 U484 ( .A1(n1371), .A2(n1136), .ZN(n1411) );
  NAND2_X2 U485 ( .A1(n1413), .A2(n1414), .ZN(n1371) );
  MUX2_X1 U486 ( .A(n1415), .B(n1416), .S(n1107), .Z(n1414) );
  NAND2_X2 U487 ( .A1(n1127), .A2(n1230), .ZN(n1416) );
  NAND2_X2 U488 ( .A1(n1127), .A2(n1229), .ZN(n1415) );
  MUX2_X1 U489 ( .A(n1417), .B(n1418), .S(n1107), .Z(n1413) );
  NAND2_X2 U490 ( .A1(n1234), .A2(n1117), .ZN(n1418) );
  NAND2_X2 U491 ( .A1(n1233), .A2(n1117), .ZN(n1417) );
  NAND2_X2 U492 ( .A1(n1419), .A2(n1420), .ZN(B[1]) );
  MUX2_X1 U493 ( .A(n1421), .B(n1422), .S(n1157), .Z(n1420) );
  NAND2_X2 U494 ( .A1(n1144), .A2(n1260), .ZN(n1422) );
  NAND2_X2 U495 ( .A1(n1144), .A2(n1261), .ZN(n1421) );
  MUX2_X1 U496 ( .A(n1423), .B(n1424), .S(n1157), .Z(n1419) );
  NAND2_X2 U497 ( .A1(n1239), .A2(n1135), .ZN(n1424) );
  NAND2_X2 U498 ( .A1(n1222), .A2(n1135), .ZN(n1423) );
  NAND2_X2 U499 ( .A1(n1425), .A2(n1426), .ZN(n1222) );
  MUX2_X1 U500 ( .A(n1427), .B(n1428), .S(n1107), .Z(n1426) );
  NAND2_X2 U501 ( .A1(n1127), .A2(n1429), .ZN(n1428) );
  NAND2_X2 U502 ( .A1(n1126), .A2(n1430), .ZN(n1427) );
  MUX2_X1 U503 ( .A(n1431), .B(n1432), .S(n1107), .Z(n1425) );
  NAND2_X2 U504 ( .A1(n1212), .A2(n1116), .ZN(n1432) );
  NAND2_X2 U505 ( .A1(n1213), .A2(n1116), .ZN(n1431) );
  NAND2_X2 U506 ( .A1(n1433), .A2(n1434), .ZN(B[19]) );
  MUX2_X1 U507 ( .A(n1435), .B(n1436), .S(n1157), .Z(n1434) );
  NAND2_X2 U508 ( .A1(n1144), .A2(n1437), .ZN(n1436) );
  NAND2_X2 U509 ( .A1(n1144), .A2(n1410), .ZN(n1435) );
  MUX2_X1 U510 ( .A(n1438), .B(n1439), .S(n1157), .Z(n1433) );
  NAND2_X2 U511 ( .A1(n1397), .A2(n1135), .ZN(n1439) );
  NAND2_X2 U512 ( .A1(n1384), .A2(n1135), .ZN(n1438) );
  NAND2_X2 U513 ( .A1(n1440), .A2(n1441), .ZN(n1384) );
  MUX2_X1 U514 ( .A(n1442), .B(n1443), .S(n1107), .Z(n1441) );
  NAND2_X2 U515 ( .A1(n1126), .A2(n1247), .ZN(n1443) );
  NAND2_X2 U516 ( .A1(n1126), .A2(n1246), .ZN(n1442) );
  MUX2_X1 U517 ( .A(n1444), .B(n1445), .S(n1107), .Z(n1440) );
  NAND2_X2 U518 ( .A1(n1251), .A2(n1116), .ZN(n1445) );
  NAND2_X2 U519 ( .A1(n1250), .A2(n1116), .ZN(n1444) );
  NAND2_X2 U520 ( .A1(n1446), .A2(n1447), .ZN(B[18]) );
  MUX2_X1 U521 ( .A(n1448), .B(n1449), .S(n1157), .Z(n1447) );
  NAND2_X2 U522 ( .A1(n1143), .A2(n1450), .ZN(n1449) );
  NAND2_X2 U523 ( .A1(n1143), .A2(n1437), .ZN(n1448) );
  MUX2_X1 U524 ( .A(n1451), .B(n1452), .S(n1157), .Z(n1446) );
  NAND2_X2 U525 ( .A1(n1410), .A2(n1135), .ZN(n1452) );
  NAND2_X2 U526 ( .A1(n1397), .A2(n1135), .ZN(n1451) );
  NAND2_X2 U527 ( .A1(n1453), .A2(n1454), .ZN(n1397) );
  MUX2_X1 U528 ( .A(n1455), .B(n1456), .S(n1107), .Z(n1454) );
  NAND2_X2 U529 ( .A1(n1126), .A2(n1280), .ZN(n1456) );
  NAND2_X2 U530 ( .A1(n1126), .A2(n1279), .ZN(n1455) );
  MUX2_X1 U531 ( .A(n1457), .B(n1458), .S(n1107), .Z(n1453) );
  NAND2_X2 U532 ( .A1(n1196), .A2(n1116), .ZN(n1458) );
  INV_X2 U533 ( .A(n1459), .ZN(n1196) );
  MUX2_X1 U534 ( .A(n1460), .B(n1461), .S(n1111), .Z(n1459) );
  NAND2_X2 U535 ( .A1(n1195), .A2(n1116), .ZN(n1457) );
  INV_X2 U536 ( .A(n1462), .ZN(n1195) );
  MUX2_X1 U537 ( .A(n1463), .B(n1464), .S(n1111), .Z(n1462) );
  NAND2_X2 U538 ( .A1(n1465), .A2(n1466), .ZN(B[17]) );
  MUX2_X1 U539 ( .A(n1467), .B(n1468), .S(n1157), .Z(n1466) );
  NAND2_X2 U540 ( .A1(n1143), .A2(n1469), .ZN(n1468) );
  NAND2_X2 U541 ( .A1(n1143), .A2(n1450), .ZN(n1467) );
  MUX2_X1 U542 ( .A(n1470), .B(n1471), .S(n1157), .Z(n1465) );
  NAND2_X2 U543 ( .A1(n1437), .A2(n1135), .ZN(n1471) );
  NAND2_X2 U544 ( .A1(n1410), .A2(n1135), .ZN(n1470) );
  NAND2_X2 U545 ( .A1(n1472), .A2(n1473), .ZN(n1410) );
  MUX2_X1 U546 ( .A(n1474), .B(n1475), .S(n1107), .Z(n1473) );
  NAND2_X2 U547 ( .A1(n1125), .A2(n1430), .ZN(n1475) );
  NAND2_X2 U548 ( .A1(n1125), .A2(n1429), .ZN(n1474) );
  MUX2_X1 U549 ( .A(n1476), .B(n1477), .S(n1107), .Z(n1472) );
  NAND2_X2 U550 ( .A1(n1213), .A2(n1116), .ZN(n1477) );
  INV_X2 U551 ( .A(n1478), .ZN(n1213) );
  MUX2_X1 U552 ( .A(n1479), .B(n1480), .S(n1111), .Z(n1478) );
  NAND2_X2 U553 ( .A1(n1212), .A2(n1116), .ZN(n1476) );
  INV_X2 U554 ( .A(n1481), .ZN(n1212) );
  MUX2_X1 U555 ( .A(n1482), .B(n1483), .S(n1111), .Z(n1481) );
  NAND2_X2 U556 ( .A1(n1484), .A2(n1485), .ZN(B[16]) );
  MUX2_X1 U557 ( .A(n1486), .B(n1487), .S(n1158), .Z(n1485) );
  NAND2_X2 U558 ( .A1(n1143), .A2(n1488), .ZN(n1487) );
  NAND2_X2 U559 ( .A1(n1142), .A2(n1469), .ZN(n1486) );
  MUX2_X1 U560 ( .A(n1489), .B(n1490), .S(n1158), .Z(n1484) );
  NAND2_X2 U561 ( .A1(n1450), .A2(n1135), .ZN(n1490) );
  NAND2_X2 U562 ( .A1(n1437), .A2(n1135), .ZN(n1489) );
  NAND2_X2 U563 ( .A1(n1491), .A2(n1492), .ZN(n1437) );
  MUX2_X1 U564 ( .A(n1493), .B(n1494), .S(n1108), .Z(n1492) );
  NAND2_X2 U565 ( .A1(n1125), .A2(n1306), .ZN(n1494) );
  NAND2_X2 U566 ( .A1(n1125), .A2(n1305), .ZN(n1493) );
  MUX2_X1 U567 ( .A(n1495), .B(n1496), .S(n1108), .Z(n1491) );
  NAND2_X2 U568 ( .A1(n1230), .A2(n1116), .ZN(n1496) );
  NAND2_X2 U569 ( .A1(n1229), .A2(n1116), .ZN(n1495) );
  NAND2_X2 U570 ( .A1(n1497), .A2(n1498), .ZN(B[15]) );
  MUX2_X1 U571 ( .A(n1499), .B(n1500), .S(n1158), .Z(n1498) );
  NAND2_X2 U572 ( .A1(n1142), .A2(n1501), .ZN(n1500) );
  NAND2_X2 U573 ( .A1(n1142), .A2(n1488), .ZN(n1499) );
  MUX2_X1 U574 ( .A(n1502), .B(n1503), .S(n1158), .Z(n1497) );
  NAND2_X2 U575 ( .A1(n1469), .A2(n1135), .ZN(n1503) );
  NAND2_X2 U576 ( .A1(n1450), .A2(n1135), .ZN(n1502) );
  NAND2_X2 U577 ( .A1(n1504), .A2(n1505), .ZN(n1450) );
  MUX2_X1 U578 ( .A(n1506), .B(n1507), .S(n1108), .Z(n1505) );
  NAND2_X2 U579 ( .A1(n1125), .A2(n1323), .ZN(n1507) );
  NAND2_X2 U580 ( .A1(n1124), .A2(n1322), .ZN(n1506) );
  MUX2_X1 U581 ( .A(n1508), .B(n1509), .S(n1108), .Z(n1504) );
  NAND2_X2 U582 ( .A1(n1247), .A2(n1116), .ZN(n1509) );
  NAND2_X2 U583 ( .A1(n1246), .A2(n1116), .ZN(n1508) );
  NAND2_X2 U584 ( .A1(n1510), .A2(n1511), .ZN(B[14]) );
  MUX2_X1 U585 ( .A(n1512), .B(n1513), .S(n1158), .Z(n1511) );
  NAND2_X2 U586 ( .A1(n1142), .A2(n1514), .ZN(n1513) );
  NAND2_X2 U587 ( .A1(n1142), .A2(n1501), .ZN(n1512) );
  MUX2_X1 U588 ( .A(n1515), .B(n1516), .S(n1158), .Z(n1510) );
  NAND2_X2 U589 ( .A1(n1488), .A2(n1134), .ZN(n1516) );
  NAND2_X2 U590 ( .A1(n1469), .A2(n1134), .ZN(n1515) );
  NAND2_X2 U591 ( .A1(n1517), .A2(n1518), .ZN(n1469) );
  MUX2_X1 U592 ( .A(n1519), .B(n1520), .S(n1108), .Z(n1518) );
  NAND2_X2 U593 ( .A1(n1124), .A2(n1338), .ZN(n1520) );
  NAND2_X2 U594 ( .A1(n1124), .A2(n1337), .ZN(n1519) );
  MUX2_X1 U595 ( .A(n1521), .B(n1522), .S(n1108), .Z(n1517) );
  NAND2_X2 U596 ( .A1(n1280), .A2(n1115), .ZN(n1522) );
  NAND2_X2 U597 ( .A1(n1279), .A2(n1115), .ZN(n1521) );
  NAND2_X2 U598 ( .A1(n1523), .A2(n1524), .ZN(B[13]) );
  MUX2_X1 U599 ( .A(n1525), .B(n1526), .S(n1158), .Z(n1524) );
  NAND2_X2 U600 ( .A1(n1141), .A2(n1527), .ZN(n1526) );
  NAND2_X2 U601 ( .A1(n1141), .A2(n1514), .ZN(n1525) );
  MUX2_X1 U602 ( .A(n1528), .B(n1529), .S(n1158), .Z(n1523) );
  NAND2_X2 U603 ( .A1(n1501), .A2(n1134), .ZN(n1529) );
  NAND2_X2 U604 ( .A1(n1488), .A2(n1134), .ZN(n1528) );
  NAND2_X2 U605 ( .A1(n1530), .A2(n1531), .ZN(n1488) );
  MUX2_X1 U606 ( .A(n1532), .B(n1533), .S(n1108), .Z(n1531) );
  NAND2_X2 U607 ( .A1(n1124), .A2(n1353), .ZN(n1533) );
  NAND2_X2 U608 ( .A1(n1124), .A2(n1352), .ZN(n1532) );
  MUX2_X1 U609 ( .A(n1534), .B(n1535), .S(n1108), .Z(n1530) );
  NAND2_X2 U610 ( .A1(n1430), .A2(n1115), .ZN(n1535) );
  NAND2_X2 U611 ( .A1(n1429), .A2(n1115), .ZN(n1534) );
  NAND2_X2 U612 ( .A1(n1536), .A2(n1537), .ZN(B[12]) );
  MUX2_X1 U613 ( .A(n1538), .B(n1539), .S(n1158), .Z(n1537) );
  NAND2_X2 U614 ( .A1(n1141), .A2(n1169), .ZN(n1539) );
  NAND2_X2 U615 ( .A1(n1141), .A2(n1527), .ZN(n1538) );
  MUX2_X1 U616 ( .A(n1540), .B(n1541), .S(n1158), .Z(n1536) );
  NAND2_X2 U617 ( .A1(n1514), .A2(n1134), .ZN(n1541) );
  NAND2_X2 U618 ( .A1(n1501), .A2(n1134), .ZN(n1540) );
  NAND2_X2 U619 ( .A1(n1542), .A2(n1543), .ZN(n1501) );
  MUX2_X1 U620 ( .A(n1544), .B(n1545), .S(n1108), .Z(n1543) );
  NAND2_X2 U621 ( .A1(n1123), .A2(n1302), .ZN(n1545) );
  NAND2_X2 U622 ( .A1(n1123), .A2(n1301), .ZN(n1544) );
  MUX2_X1 U623 ( .A(n1546), .B(n1547), .S(n1108), .Z(n1542) );
  NAND2_X2 U624 ( .A1(n1306), .A2(n1115), .ZN(n1547) );
  NAND2_X2 U625 ( .A1(n1305), .A2(n1115), .ZN(n1546) );
  NAND2_X2 U626 ( .A1(n1548), .A2(n1549), .ZN(B[11]) );
  MUX2_X1 U627 ( .A(n1550), .B(n1551), .S(n1158), .Z(n1549) );
  NAND2_X2 U628 ( .A1(n1141), .A2(n1168), .ZN(n1551) );
  NAND2_X2 U629 ( .A1(n1140), .A2(n1169), .ZN(n1550) );
  MUX2_X1 U630 ( .A(n1552), .B(n1553), .S(n1158), .Z(n1548) );
  NAND2_X2 U631 ( .A1(n1527), .A2(n1134), .ZN(n1553) );
  NAND2_X2 U632 ( .A1(n1514), .A2(n1134), .ZN(n1552) );
  NAND2_X2 U633 ( .A1(n1554), .A2(n1555), .ZN(n1514) );
  MUX2_X1 U634 ( .A(n1556), .B(n1557), .S(n1108), .Z(n1555) );
  NAND2_X2 U635 ( .A1(n1123), .A2(n1319), .ZN(n1557) );
  NAND2_X2 U636 ( .A1(n1123), .A2(n1318), .ZN(n1556) );
  MUX2_X1 U637 ( .A(n1558), .B(n1559), .S(n1108), .Z(n1554) );
  NAND2_X2 U638 ( .A1(n1323), .A2(n1115), .ZN(n1559) );
  NAND2_X2 U639 ( .A1(n1322), .A2(n1115), .ZN(n1558) );
  NAND2_X2 U640 ( .A1(n1560), .A2(n1561), .ZN(B[10]) );
  MUX2_X1 U641 ( .A(n1562), .B(n1563), .S(n1159), .Z(n1561) );
  NAND2_X2 U642 ( .A1(n1140), .A2(n1165), .ZN(n1563) );
  NAND2_X2 U643 ( .A1(n1564), .A2(n1565), .ZN(n1165) );
  MUX2_X1 U644 ( .A(n1566), .B(n1567), .S(n1109), .Z(n1565) );
  NAND2_X2 U645 ( .A1(n1123), .A2(n1250), .ZN(n1567) );
  INV_X2 U646 ( .A(n1568), .ZN(n1250) );
  MUX2_X1 U647 ( .A(n1569), .B(n1570), .S(n1111), .Z(n1568) );
  NAND2_X2 U648 ( .A1(n1122), .A2(n1251), .ZN(n1566) );
  INV_X2 U649 ( .A(n1571), .ZN(n1251) );
  MUX2_X1 U650 ( .A(n1572), .B(n1573), .S(n1111), .Z(n1571) );
  MUX2_X1 U651 ( .A(n1574), .B(n1575), .S(n1109), .Z(n1564) );
  NAND2_X2 U652 ( .A1(n1319), .A2(n1115), .ZN(n1575) );
  INV_X2 U653 ( .A(n1576), .ZN(n1319) );
  MUX2_X1 U654 ( .A(n1577), .B(n1578), .S(n1111), .Z(n1576) );
  NAND2_X2 U655 ( .A1(n1318), .A2(n1115), .ZN(n1574) );
  INV_X2 U656 ( .A(n1579), .ZN(n1318) );
  MUX2_X1 U657 ( .A(n1580), .B(n1581), .S(n1111), .Z(n1579) );
  NAND2_X2 U658 ( .A1(n1140), .A2(n1168), .ZN(n1562) );
  NAND2_X2 U659 ( .A1(n1582), .A2(n1583), .ZN(n1168) );
  MUX2_X1 U660 ( .A(n1584), .B(n1585), .S(n1109), .Z(n1583) );
  NAND2_X2 U661 ( .A1(n1122), .A2(n1233), .ZN(n1585) );
  INV_X2 U662 ( .A(n1586), .ZN(n1233) );
  MUX2_X1 U663 ( .A(n1587), .B(n1588), .S(n1111), .Z(n1586) );
  NAND2_X2 U664 ( .A1(n1122), .A2(n1234), .ZN(n1584) );
  INV_X2 U665 ( .A(n1589), .ZN(n1234) );
  MUX2_X1 U666 ( .A(n1590), .B(n1591), .S(n1111), .Z(n1589) );
  MUX2_X1 U667 ( .A(n1592), .B(n1593), .S(n1109), .Z(n1582) );
  NAND2_X2 U668 ( .A1(n1302), .A2(n1115), .ZN(n1593) );
  INV_X2 U669 ( .A(n1594), .ZN(n1302) );
  MUX2_X1 U670 ( .A(n1595), .B(n1596), .S(n1111), .Z(n1594) );
  NAND2_X2 U671 ( .A1(n1301), .A2(n1115), .ZN(n1592) );
  INV_X2 U672 ( .A(n1597), .ZN(n1301) );
  MUX2_X1 U673 ( .A(n1598), .B(n1599), .S(n1111), .Z(n1597) );
  MUX2_X1 U674 ( .A(n1600), .B(n1601), .S(n1159), .Z(n1560) );
  NAND2_X2 U675 ( .A1(n1169), .A2(n1134), .ZN(n1601) );
  NAND2_X2 U676 ( .A1(n1602), .A2(n1603), .ZN(n1169) );
  MUX2_X1 U677 ( .A(n1604), .B(n1605), .S(n1109), .Z(n1603) );
  NAND2_X2 U678 ( .A1(n1122), .A2(n1216), .ZN(n1605) );
  INV_X2 U679 ( .A(n1606), .ZN(n1216) );
  MUX2_X1 U680 ( .A(n1607), .B(n1608), .S(n1112), .Z(n1606) );
  NAND2_X2 U681 ( .A1(n1122), .A2(n1217), .ZN(n1604) );
  INV_X2 U682 ( .A(n1609), .ZN(n1217) );
  MUX2_X1 U683 ( .A(n1610), .B(n1611), .S(n1112), .Z(n1609) );
  MUX2_X1 U684 ( .A(n1612), .B(n1613), .S(n1109), .Z(n1602) );
  NAND2_X2 U685 ( .A1(n1353), .A2(n1114), .ZN(n1613) );
  NAND2_X2 U686 ( .A1(n1352), .A2(n1114), .ZN(n1612) );
  NAND2_X2 U687 ( .A1(n1527), .A2(n1134), .ZN(n1600) );
  NAND2_X2 U688 ( .A1(n1614), .A2(n1615), .ZN(n1527) );
  MUX2_X1 U689 ( .A(n1616), .B(n1617), .S(n1109), .Z(n1615) );
  NAND2_X2 U690 ( .A1(n1121), .A2(n1199), .ZN(n1617) );
  INV_X2 U691 ( .A(n1618), .ZN(n1199) );
  MUX2_X1 U692 ( .A(n1619), .B(n1620), .S(n1112), .Z(n1618) );
  NAND2_X2 U693 ( .A1(n1121), .A2(n1200), .ZN(n1616) );
  INV_X2 U694 ( .A(n1621), .ZN(n1200) );
  MUX2_X1 U695 ( .A(n1622), .B(n1623), .S(n1112), .Z(n1621) );
  MUX2_X1 U696 ( .A(n1624), .B(n1625), .S(n1109), .Z(n1614) );
  NAND2_X2 U697 ( .A1(n1338), .A2(n1114), .ZN(n1625) );
  NAND2_X2 U698 ( .A1(n1337), .A2(n1114), .ZN(n1624) );
  NAND2_X2 U699 ( .A1(n1626), .A2(n1627), .ZN(B[0]) );
  MUX2_X1 U700 ( .A(n1628), .B(n1629), .S(n1159), .Z(n1627) );
  NAND2_X2 U701 ( .A1(n1140), .A2(n1257), .ZN(n1629) );
  NAND2_X2 U702 ( .A1(n1630), .A2(n1631), .ZN(n1257) );
  MUX2_X1 U703 ( .A(n1632), .B(n1633), .S(n1109), .Z(n1631) );
  NAND2_X2 U704 ( .A1(n1121), .A2(n1352), .ZN(n1633) );
  INV_X2 U705 ( .A(n1634), .ZN(n1352) );
  MUX2_X1 U706 ( .A(n1483), .B(n1479), .S(n1112), .Z(n1634) );
  NAND2_X2 U707 ( .A1(n1121), .A2(n1353), .ZN(n1632) );
  INV_X2 U708 ( .A(n1635), .ZN(n1353) );
  MUX2_X1 U709 ( .A(n1480), .B(n1482), .S(n1112), .Z(n1635) );
  MUX2_X1 U710 ( .A(n1636), .B(n1637), .S(n1109), .Z(n1630) );
  NAND2_X2 U711 ( .A1(n1429), .A2(n1114), .ZN(n1637) );
  INV_X2 U712 ( .A(n1638), .ZN(n1429) );
  MUX2_X1 U713 ( .A(n1608), .B(n1610), .S(n1112), .Z(n1638) );
  NAND2_X2 U714 ( .A1(n1430), .A2(n1114), .ZN(n1636) );
  INV_X2 U715 ( .A(n1639), .ZN(n1430) );
  MUX2_X1 U716 ( .A(n1611), .B(n1607), .S(n1112), .Z(n1639) );
  NAND2_X2 U717 ( .A1(n1140), .A2(n1260), .ZN(n1628) );
  NAND2_X2 U718 ( .A1(n1640), .A2(n1641), .ZN(n1260) );
  MUX2_X1 U719 ( .A(n1642), .B(n1643), .S(n1109), .Z(n1641) );
  NAND2_X2 U720 ( .A1(n1121), .A2(n1337), .ZN(n1643) );
  INV_X2 U721 ( .A(n1644), .ZN(n1337) );
  MUX2_X1 U722 ( .A(n1464), .B(n1460), .S(n1112), .Z(n1644) );
  NAND2_X2 U723 ( .A1(n1120), .A2(n1338), .ZN(n1642) );
  INV_X2 U724 ( .A(n1645), .ZN(n1338) );
  MUX2_X1 U725 ( .A(n1461), .B(n1463), .S(n1112), .Z(n1645) );
  MUX2_X1 U726 ( .A(n1646), .B(n1647), .S(n1109), .Z(n1640) );
  NAND2_X2 U727 ( .A1(n1279), .A2(n1114), .ZN(n1647) );
  INV_X2 U728 ( .A(n1648), .ZN(n1279) );
  MUX2_X1 U729 ( .A(n1620), .B(n1622), .S(n1112), .Z(n1648) );
  NAND2_X2 U730 ( .A1(n1280), .A2(n1114), .ZN(n1646) );
  INV_X2 U731 ( .A(n1649), .ZN(n1280) );
  MUX2_X1 U732 ( .A(n1623), .B(n1619), .S(n1112), .Z(n1649) );
  MUX2_X1 U733 ( .A(n1650), .B(n1651), .S(n1159), .Z(n1626) );
  NAND2_X2 U734 ( .A1(n1261), .A2(n1134), .ZN(n1651) );
  NAND2_X2 U735 ( .A1(n1652), .A2(n1653), .ZN(n1261) );
  MUX2_X1 U736 ( .A(n1654), .B(n1655), .S(n1110), .Z(n1653) );
  NAND2_X2 U737 ( .A1(n1120), .A2(n1322), .ZN(n1655) );
  INV_X2 U738 ( .A(n1656), .ZN(n1322) );
  MUX2_X1 U739 ( .A(n1570), .B(n1572), .S(n1113), .Z(n1656) );
  INV_X2 U740 ( .A(A[3]), .ZN(n1572) );
  NAND2_X2 U741 ( .A1(n1120), .A2(n1323), .ZN(n1654) );
  INV_X2 U742 ( .A(n1657), .ZN(n1323) );
  MUX2_X1 U743 ( .A(n1573), .B(n1569), .S(n1113), .Z(n1657) );
  MUX2_X1 U744 ( .A(n1658), .B(n1659), .S(n1110), .Z(n1652) );
  NAND2_X2 U745 ( .A1(n1246), .A2(n1114), .ZN(n1659) );
  INV_X2 U746 ( .A(n1660), .ZN(n1246) );
  MUX2_X1 U747 ( .A(n1578), .B(n1580), .S(n1113), .Z(n1660) );
  NAND2_X2 U748 ( .A1(n1247), .A2(n1114), .ZN(n1658) );
  INV_X2 U749 ( .A(n1661), .ZN(n1247) );
  MUX2_X1 U750 ( .A(n1581), .B(n1577), .S(n1113), .Z(n1661) );
  INV_X2 U751 ( .A(A[23]), .ZN(n1577) );
  NAND2_X2 U752 ( .A1(n1239), .A2(n1134), .ZN(n1650) );
  NAND2_X2 U753 ( .A1(n1662), .A2(n1663), .ZN(n1239) );
  MUX2_X1 U754 ( .A(n1664), .B(n1665), .S(n1110), .Z(n1663) );
  NAND2_X2 U755 ( .A1(n1120), .A2(n1305), .ZN(n1665) );
  INV_X2 U756 ( .A(n1666), .ZN(n1305) );
  MUX2_X1 U757 ( .A(n1588), .B(n1590), .S(n1113), .Z(n1666) );
  NAND2_X2 U758 ( .A1(n1120), .A2(n1306), .ZN(n1664) );
  INV_X2 U759 ( .A(n1667), .ZN(n1306) );
  MUX2_X1 U760 ( .A(n1591), .B(n1587), .S(n1113), .Z(n1667) );
  MUX2_X1 U761 ( .A(n1668), .B(n1669), .S(n1110), .Z(n1662) );
  NAND2_X2 U762 ( .A1(n1229), .A2(n1114), .ZN(n1669) );
  INV_X2 U763 ( .A(n1670), .ZN(n1229) );
  MUX2_X1 U764 ( .A(n1596), .B(n1598), .S(n1113), .Z(n1670) );
  NAND2_X2 U765 ( .A1(n1230), .A2(n1114), .ZN(n1668) );
  INV_X2 U766 ( .A(n1671), .ZN(n1230) );
  MUX2_X1 U767 ( .A(n1599), .B(n1595), .S(n1113), .Z(n1671) );
endmodule


module Xi_core_DW_rbsh_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672;

  INV_X1 U170 ( .A(A[24]), .ZN(n1480) );
  INV_X1 U171 ( .A(A[26]), .ZN(n1617) );
  INV_X1 U172 ( .A(A[28]), .ZN(n1602) );
  INV_X1 U173 ( .A(A[1]), .ZN(n1462) );
  INV_X1 U174 ( .A(A[25]), .ZN(n1461) );
  INV_X1 U175 ( .A(A[30]), .ZN(n1614) );
  INV_X1 U176 ( .A(A[0]), .ZN(n1481) );
  INV_X1 U177 ( .A(A[2]), .ZN(n1618) );
  INV_X1 U178 ( .A(A[29]), .ZN(n1570) );
  INV_X1 U179 ( .A(A[4]), .ZN(n1603) );
  INV_X1 U180 ( .A(A[22]), .ZN(n1623) );
  INV_X1 U181 ( .A(A[27]), .ZN(n1585) );
  INV_X1 U182 ( .A(A[21]), .ZN(n1576) );
  INV_X1 U183 ( .A(A[31]), .ZN(n1582) );
  INV_X1 U184 ( .A(A[6]), .ZN(n1615) );
  INV_X1 U185 ( .A(A[7]), .ZN(n1583) );
  INV_X1 U186 ( .A(A[5]), .ZN(n1571) );
  INV_X1 U187 ( .A(A[19]), .ZN(n1594) );
  INV_X1 U188 ( .A(A[18]), .ZN(n1626) );
  INV_X1 U189 ( .A(A[16]), .ZN(n1476) );
  INV_X1 U190 ( .A(A[13]), .ZN(n1575) );
  INV_X1 U191 ( .A(A[17]), .ZN(n1457) );
  INV_X1 U192 ( .A(A[15]), .ZN(n1590) );
  INV_X1 U193 ( .A(A[14]), .ZN(n1622) );
  INV_X1 U194 ( .A(A[20]), .ZN(n1608) );
  INV_X1 U195 ( .A(A[12]), .ZN(n1607) );
  INV_X1 U196 ( .A(A[9]), .ZN(n1456) );
  INV_X1 U197 ( .A(A[11]), .ZN(n1593) );
  INV_X1 U198 ( .A(A[8]), .ZN(n1475) );
  INV_X1 U199 ( .A(A[10]), .ZN(n1625) );
  INV_X1 U200 ( .A(n1124), .ZN(n1106) );
  INV_X1 U201 ( .A(n1124), .ZN(n1107) );
  INV_X1 U202 ( .A(n1125), .ZN(n1108) );
  INV_X1 U203 ( .A(n1125), .ZN(n1109) );
  INV_X1 U204 ( .A(n1125), .ZN(n1110) );
  INV_X1 U205 ( .A(n1125), .ZN(n1111) );
  CLKBUF_X3 U206 ( .A(SH[4]), .Z(n1112) );
  CLKBUF_X3 U207 ( .A(SH[4]), .Z(n1113) );
  CLKBUF_X3 U208 ( .A(SH[4]), .Z(n1114) );
  CLKBUF_X3 U209 ( .A(SH[4]), .Z(n1115) );
  CLKBUF_X3 U210 ( .A(SH[4]), .Z(n1116) );
  CLKBUF_X3 U211 ( .A(SH[4]), .Z(n1117) );
  CLKBUF_X3 U212 ( .A(SH[4]), .Z(n1118) );
  CLKBUF_X3 U213 ( .A(SH[4]), .Z(n1119) );
  CLKBUF_X3 U214 ( .A(SH[4]), .Z(n1120) );
  CLKBUF_X3 U215 ( .A(SH[4]), .Z(n1121) );
  CLKBUF_X3 U216 ( .A(SH[4]), .Z(n1122) );
  CLKBUF_X3 U217 ( .A(SH[4]), .Z(n1123) );
  CLKBUF_X3 U218 ( .A(SH[4]), .Z(n1124) );
  CLKBUF_X3 U219 ( .A(SH[4]), .Z(n1125) );
  CLKBUF_X3 U220 ( .A(SH[3]), .Z(n1126) );
  CLKBUF_X3 U221 ( .A(SH[3]), .Z(n1127) );
  CLKBUF_X3 U222 ( .A(SH[3]), .Z(n1128) );
  CLKBUF_X3 U223 ( .A(SH[2]), .Z(n1129) );
  CLKBUF_X3 U224 ( .A(SH[2]), .Z(n1130) );
  CLKBUF_X3 U225 ( .A(SH[2]), .Z(n1131) );
  CLKBUF_X3 U226 ( .A(SH[2]), .Z(n1132) );
  CLKBUF_X3 U227 ( .A(SH[2]), .Z(n1133) );
  CLKBUF_X3 U228 ( .A(SH[2]), .Z(n1134) );
  CLKBUF_X3 U229 ( .A(SH[1]), .Z(n1135) );
  CLKBUF_X3 U230 ( .A(SH[1]), .Z(n1136) );
  CLKBUF_X3 U231 ( .A(SH[1]), .Z(n1137) );
  CLKBUF_X3 U232 ( .A(SH[1]), .Z(n1138) );
  CLKBUF_X3 U233 ( .A(SH[1]), .Z(n1139) );
  CLKBUF_X3 U234 ( .A(SH[1]), .Z(n1140) );
  INV_X1 U235 ( .A(n1159), .ZN(n1141) );
  INV_X1 U236 ( .A(n1159), .ZN(n1142) );
  INV_X1 U237 ( .A(n1160), .ZN(n1143) );
  INV_X1 U238 ( .A(n1160), .ZN(n1144) );
  INV_X1 U239 ( .A(n1160), .ZN(n1145) );
  INV_X1 U240 ( .A(n1160), .ZN(n1146) );
  CLKBUF_X3 U241 ( .A(SH[0]), .Z(n1147) );
  CLKBUF_X3 U242 ( .A(SH[0]), .Z(n1148) );
  CLKBUF_X3 U243 ( .A(SH[0]), .Z(n1149) );
  CLKBUF_X3 U244 ( .A(SH[0]), .Z(n1150) );
  CLKBUF_X3 U245 ( .A(SH[0]), .Z(n1151) );
  CLKBUF_X3 U246 ( .A(SH[0]), .Z(n1152) );
  CLKBUF_X3 U247 ( .A(SH[0]), .Z(n1153) );
  CLKBUF_X3 U248 ( .A(SH[0]), .Z(n1154) );
  CLKBUF_X3 U249 ( .A(SH[0]), .Z(n1155) );
  CLKBUF_X3 U250 ( .A(SH[0]), .Z(n1156) );
  CLKBUF_X3 U251 ( .A(SH[0]), .Z(n1157) );
  CLKBUF_X3 U252 ( .A(SH[0]), .Z(n1158) );
  CLKBUF_X3 U253 ( .A(SH[0]), .Z(n1159) );
  CLKBUF_X3 U254 ( .A(SH[0]), .Z(n1160) );
  NAND2_X2 U255 ( .A1(n1161), .A2(n1162), .ZN(B[9]) );
  MUX2_X1 U256 ( .A(n1163), .B(n1164), .S(n1135), .Z(n1162) );
  NAND2_X2 U257 ( .A1(n1159), .A2(n1165), .ZN(n1164) );
  NAND2_X2 U258 ( .A1(n1159), .A2(n1166), .ZN(n1163) );
  MUX2_X1 U259 ( .A(n1167), .B(n1168), .S(n1135), .Z(n1161) );
  NAND2_X2 U260 ( .A1(n1169), .A2(n1146), .ZN(n1168) );
  NAND2_X2 U261 ( .A1(n1170), .A2(n1146), .ZN(n1167) );
  NAND2_X2 U262 ( .A1(n1171), .A2(n1172), .ZN(B[8]) );
  MUX2_X1 U263 ( .A(n1173), .B(n1174), .S(n1135), .Z(n1172) );
  NAND2_X2 U264 ( .A1(n1159), .A2(n1169), .ZN(n1174) );
  NAND2_X2 U265 ( .A1(n1159), .A2(n1170), .ZN(n1173) );
  MUX2_X1 U266 ( .A(n1175), .B(n1176), .S(n1135), .Z(n1171) );
  NAND2_X2 U267 ( .A1(n1166), .A2(n1146), .ZN(n1176) );
  NAND2_X2 U268 ( .A1(n1177), .A2(n1146), .ZN(n1175) );
  NAND2_X2 U269 ( .A1(n1178), .A2(n1179), .ZN(B[7]) );
  MUX2_X1 U270 ( .A(n1180), .B(n1181), .S(n1135), .Z(n1179) );
  NAND2_X2 U271 ( .A1(n1158), .A2(n1166), .ZN(n1181) );
  NAND2_X2 U272 ( .A1(n1158), .A2(n1177), .ZN(n1180) );
  MUX2_X1 U273 ( .A(n1182), .B(n1183), .S(n1135), .Z(n1178) );
  NAND2_X2 U274 ( .A1(n1170), .A2(n1145), .ZN(n1183) );
  NAND2_X2 U275 ( .A1(n1184), .A2(n1145), .ZN(n1182) );
  NAND2_X2 U276 ( .A1(n1185), .A2(n1186), .ZN(B[6]) );
  MUX2_X1 U277 ( .A(n1187), .B(n1188), .S(n1135), .Z(n1186) );
  NAND2_X2 U278 ( .A1(n1158), .A2(n1170), .ZN(n1188) );
  NAND2_X2 U279 ( .A1(n1189), .A2(n1190), .ZN(n1170) );
  MUX2_X1 U280 ( .A(n1191), .B(n1192), .S(n1129), .Z(n1190) );
  NAND2_X2 U281 ( .A1(n1124), .A2(n1193), .ZN(n1192) );
  NAND2_X2 U282 ( .A1(n1124), .A2(n1194), .ZN(n1191) );
  MUX2_X1 U283 ( .A(n1195), .B(n1196), .S(n1129), .Z(n1189) );
  NAND2_X2 U284 ( .A1(n1197), .A2(n1111), .ZN(n1196) );
  NAND2_X2 U285 ( .A1(n1198), .A2(n1111), .ZN(n1195) );
  NAND2_X2 U286 ( .A1(n1158), .A2(n1184), .ZN(n1187) );
  MUX2_X1 U287 ( .A(n1199), .B(n1200), .S(n1135), .Z(n1185) );
  NAND2_X2 U288 ( .A1(n1177), .A2(n1145), .ZN(n1200) );
  NAND2_X2 U289 ( .A1(n1201), .A2(n1145), .ZN(n1199) );
  NAND2_X2 U290 ( .A1(n1202), .A2(n1203), .ZN(B[5]) );
  MUX2_X1 U291 ( .A(n1204), .B(n1205), .S(n1135), .Z(n1203) );
  NAND2_X2 U292 ( .A1(n1158), .A2(n1177), .ZN(n1205) );
  NAND2_X2 U293 ( .A1(n1206), .A2(n1207), .ZN(n1177) );
  MUX2_X1 U294 ( .A(n1208), .B(n1209), .S(n1129), .Z(n1207) );
  NAND2_X2 U295 ( .A1(n1124), .A2(n1210), .ZN(n1209) );
  NAND2_X2 U296 ( .A1(n1124), .A2(n1211), .ZN(n1208) );
  MUX2_X1 U297 ( .A(n1212), .B(n1213), .S(n1129), .Z(n1206) );
  NAND2_X2 U298 ( .A1(n1214), .A2(n1111), .ZN(n1213) );
  NAND2_X2 U299 ( .A1(n1215), .A2(n1111), .ZN(n1212) );
  NAND2_X2 U300 ( .A1(n1157), .A2(n1201), .ZN(n1204) );
  MUX2_X1 U301 ( .A(n1216), .B(n1217), .S(n1135), .Z(n1202) );
  NAND2_X2 U302 ( .A1(n1184), .A2(n1145), .ZN(n1217) );
  NAND2_X2 U303 ( .A1(n1218), .A2(n1145), .ZN(n1216) );
  NAND2_X2 U304 ( .A1(n1219), .A2(n1220), .ZN(B[4]) );
  MUX2_X1 U305 ( .A(n1221), .B(n1222), .S(n1135), .Z(n1220) );
  NAND2_X2 U306 ( .A1(n1157), .A2(n1184), .ZN(n1222) );
  NAND2_X2 U307 ( .A1(n1223), .A2(n1224), .ZN(n1184) );
  MUX2_X1 U308 ( .A(n1225), .B(n1226), .S(n1129), .Z(n1224) );
  NAND2_X2 U309 ( .A1(n1123), .A2(n1227), .ZN(n1226) );
  NAND2_X2 U310 ( .A1(n1123), .A2(n1228), .ZN(n1225) );
  MUX2_X1 U311 ( .A(n1229), .B(n1230), .S(n1129), .Z(n1223) );
  NAND2_X2 U312 ( .A1(n1231), .A2(n1110), .ZN(n1230) );
  NAND2_X2 U313 ( .A1(n1232), .A2(n1110), .ZN(n1229) );
  NAND2_X2 U314 ( .A1(n1157), .A2(n1218), .ZN(n1221) );
  MUX2_X1 U315 ( .A(n1233), .B(n1234), .S(n1135), .Z(n1219) );
  NAND2_X2 U316 ( .A1(n1201), .A2(n1145), .ZN(n1234) );
  NAND2_X2 U317 ( .A1(n1235), .A2(n1145), .ZN(n1233) );
  NAND2_X2 U318 ( .A1(n1236), .A2(n1237), .ZN(B[3]) );
  MUX2_X1 U319 ( .A(n1238), .B(n1239), .S(n1136), .Z(n1237) );
  NAND2_X2 U320 ( .A1(n1157), .A2(n1201), .ZN(n1239) );
  NAND2_X2 U321 ( .A1(n1240), .A2(n1241), .ZN(n1201) );
  MUX2_X1 U322 ( .A(n1242), .B(n1243), .S(n1129), .Z(n1241) );
  NAND2_X2 U323 ( .A1(n1123), .A2(n1244), .ZN(n1243) );
  NAND2_X2 U324 ( .A1(n1123), .A2(n1245), .ZN(n1242) );
  MUX2_X1 U325 ( .A(n1246), .B(n1247), .S(n1129), .Z(n1240) );
  NAND2_X2 U326 ( .A1(n1248), .A2(n1110), .ZN(n1247) );
  NAND2_X2 U327 ( .A1(n1249), .A2(n1110), .ZN(n1246) );
  NAND2_X2 U328 ( .A1(n1157), .A2(n1235), .ZN(n1238) );
  MUX2_X1 U329 ( .A(n1250), .B(n1251), .S(n1136), .Z(n1236) );
  NAND2_X2 U330 ( .A1(n1218), .A2(n1145), .ZN(n1251) );
  NAND2_X2 U331 ( .A1(n1252), .A2(n1145), .ZN(n1250) );
  NAND2_X2 U332 ( .A1(n1253), .A2(n1254), .ZN(B[31]) );
  MUX2_X1 U333 ( .A(n1255), .B(n1256), .S(n1136), .Z(n1254) );
  NAND2_X2 U334 ( .A1(n1156), .A2(n1257), .ZN(n1256) );
  NAND2_X2 U335 ( .A1(n1156), .A2(n1258), .ZN(n1255) );
  MUX2_X1 U336 ( .A(n1259), .B(n1260), .S(n1136), .Z(n1253) );
  NAND2_X2 U337 ( .A1(n1261), .A2(n1145), .ZN(n1260) );
  NAND2_X2 U338 ( .A1(n1262), .A2(n1145), .ZN(n1259) );
  NAND2_X2 U339 ( .A1(n1263), .A2(n1264), .ZN(B[30]) );
  MUX2_X1 U340 ( .A(n1265), .B(n1266), .S(n1136), .Z(n1264) );
  NAND2_X2 U341 ( .A1(n1156), .A2(n1261), .ZN(n1266) );
  NAND2_X2 U342 ( .A1(n1156), .A2(n1262), .ZN(n1265) );
  MUX2_X1 U343 ( .A(n1267), .B(n1268), .S(n1136), .Z(n1263) );
  NAND2_X2 U344 ( .A1(n1258), .A2(n1144), .ZN(n1268) );
  NAND2_X2 U345 ( .A1(n1269), .A2(n1144), .ZN(n1267) );
  NAND2_X2 U346 ( .A1(n1270), .A2(n1271), .ZN(B[2]) );
  MUX2_X1 U347 ( .A(n1272), .B(n1273), .S(n1136), .Z(n1271) );
  NAND2_X2 U348 ( .A1(n1156), .A2(n1218), .ZN(n1273) );
  NAND2_X2 U349 ( .A1(n1274), .A2(n1275), .ZN(n1218) );
  MUX2_X1 U350 ( .A(n1276), .B(n1277), .S(n1129), .Z(n1275) );
  NAND2_X2 U351 ( .A1(n1123), .A2(n1194), .ZN(n1277) );
  NAND2_X2 U352 ( .A1(n1122), .A2(n1278), .ZN(n1276) );
  MUX2_X1 U353 ( .A(n1279), .B(n1280), .S(n1129), .Z(n1274) );
  NAND2_X2 U354 ( .A1(n1198), .A2(n1110), .ZN(n1280) );
  NAND2_X2 U355 ( .A1(n1281), .A2(n1110), .ZN(n1279) );
  NAND2_X2 U356 ( .A1(n1155), .A2(n1252), .ZN(n1272) );
  MUX2_X1 U357 ( .A(n1282), .B(n1283), .S(n1136), .Z(n1270) );
  NAND2_X2 U358 ( .A1(n1235), .A2(n1144), .ZN(n1283) );
  NAND2_X2 U359 ( .A1(n1257), .A2(n1144), .ZN(n1282) );
  NAND2_X2 U360 ( .A1(n1284), .A2(n1285), .ZN(B[29]) );
  MUX2_X1 U361 ( .A(n1286), .B(n1287), .S(n1136), .Z(n1285) );
  NAND2_X2 U362 ( .A1(n1155), .A2(n1258), .ZN(n1287) );
  NAND2_X2 U363 ( .A1(n1155), .A2(n1269), .ZN(n1286) );
  MUX2_X1 U364 ( .A(n1288), .B(n1289), .S(n1136), .Z(n1284) );
  NAND2_X2 U365 ( .A1(n1262), .A2(n1144), .ZN(n1289) );
  NAND2_X2 U366 ( .A1(n1290), .A2(n1144), .ZN(n1288) );
  NAND2_X2 U367 ( .A1(n1291), .A2(n1292), .ZN(B[28]) );
  MUX2_X1 U368 ( .A(n1293), .B(n1294), .S(n1136), .Z(n1292) );
  NAND2_X2 U369 ( .A1(n1155), .A2(n1262), .ZN(n1294) );
  NAND2_X2 U370 ( .A1(n1295), .A2(n1296), .ZN(n1262) );
  MUX2_X1 U371 ( .A(n1297), .B(n1298), .S(n1129), .Z(n1296) );
  NAND2_X2 U372 ( .A1(n1122), .A2(n1299), .ZN(n1298) );
  NAND2_X2 U373 ( .A1(n1122), .A2(n1300), .ZN(n1297) );
  MUX2_X1 U374 ( .A(n1301), .B(n1302), .S(n1129), .Z(n1295) );
  NAND2_X2 U375 ( .A1(n1303), .A2(n1110), .ZN(n1302) );
  NAND2_X2 U376 ( .A1(n1304), .A2(n1110), .ZN(n1301) );
  NAND2_X2 U377 ( .A1(n1155), .A2(n1290), .ZN(n1293) );
  MUX2_X1 U378 ( .A(n1305), .B(n1306), .S(n1136), .Z(n1291) );
  NAND2_X2 U379 ( .A1(n1269), .A2(n1144), .ZN(n1306) );
  NAND2_X2 U380 ( .A1(n1307), .A2(n1144), .ZN(n1305) );
  NAND2_X2 U381 ( .A1(n1308), .A2(n1309), .ZN(B[27]) );
  MUX2_X1 U382 ( .A(n1310), .B(n1311), .S(n1137), .Z(n1309) );
  NAND2_X2 U383 ( .A1(n1154), .A2(n1269), .ZN(n1311) );
  NAND2_X2 U384 ( .A1(n1312), .A2(n1313), .ZN(n1269) );
  MUX2_X1 U385 ( .A(n1314), .B(n1315), .S(n1130), .Z(n1313) );
  NAND2_X2 U386 ( .A1(n1122), .A2(n1316), .ZN(n1315) );
  NAND2_X2 U387 ( .A1(n1122), .A2(n1317), .ZN(n1314) );
  MUX2_X1 U388 ( .A(n1318), .B(n1319), .S(n1130), .Z(n1312) );
  NAND2_X2 U389 ( .A1(n1320), .A2(n1110), .ZN(n1319) );
  NAND2_X2 U390 ( .A1(n1321), .A2(n1110), .ZN(n1318) );
  NAND2_X2 U391 ( .A1(n1154), .A2(n1307), .ZN(n1310) );
  MUX2_X1 U392 ( .A(n1322), .B(n1323), .S(n1137), .Z(n1308) );
  NAND2_X2 U393 ( .A1(n1290), .A2(n1144), .ZN(n1323) );
  NAND2_X2 U394 ( .A1(n1324), .A2(n1144), .ZN(n1322) );
  NAND2_X2 U395 ( .A1(n1325), .A2(n1326), .ZN(B[26]) );
  MUX2_X1 U396 ( .A(n1327), .B(n1328), .S(n1137), .Z(n1326) );
  NAND2_X2 U397 ( .A1(n1154), .A2(n1290), .ZN(n1328) );
  NAND2_X2 U398 ( .A1(n1329), .A2(n1330), .ZN(n1290) );
  MUX2_X1 U399 ( .A(n1331), .B(n1332), .S(n1130), .Z(n1330) );
  NAND2_X2 U400 ( .A1(n1121), .A2(n1333), .ZN(n1332) );
  NAND2_X2 U401 ( .A1(n1121), .A2(n1197), .ZN(n1331) );
  MUX2_X1 U402 ( .A(n1334), .B(n1335), .S(n1130), .Z(n1329) );
  NAND2_X2 U403 ( .A1(n1336), .A2(n1110), .ZN(n1335) );
  NAND2_X2 U404 ( .A1(n1193), .A2(n1110), .ZN(n1334) );
  NAND2_X2 U405 ( .A1(n1154), .A2(n1324), .ZN(n1327) );
  MUX2_X1 U406 ( .A(n1337), .B(n1338), .S(n1137), .Z(n1325) );
  NAND2_X2 U407 ( .A1(n1307), .A2(n1144), .ZN(n1338) );
  NAND2_X2 U408 ( .A1(n1339), .A2(n1144), .ZN(n1337) );
  NAND2_X2 U409 ( .A1(n1340), .A2(n1341), .ZN(B[25]) );
  MUX2_X1 U410 ( .A(n1342), .B(n1343), .S(n1137), .Z(n1341) );
  NAND2_X2 U411 ( .A1(n1154), .A2(n1307), .ZN(n1343) );
  NAND2_X2 U412 ( .A1(n1344), .A2(n1345), .ZN(n1307) );
  MUX2_X1 U413 ( .A(n1346), .B(n1347), .S(n1130), .Z(n1345) );
  NAND2_X2 U414 ( .A1(n1121), .A2(n1348), .ZN(n1347) );
  NAND2_X2 U415 ( .A1(n1121), .A2(n1214), .ZN(n1346) );
  MUX2_X1 U416 ( .A(n1349), .B(n1350), .S(n1130), .Z(n1344) );
  NAND2_X2 U417 ( .A1(n1351), .A2(n1109), .ZN(n1350) );
  NAND2_X2 U418 ( .A1(n1210), .A2(n1109), .ZN(n1349) );
  NAND2_X2 U419 ( .A1(n1153), .A2(n1339), .ZN(n1342) );
  MUX2_X1 U420 ( .A(n1352), .B(n1353), .S(n1137), .Z(n1340) );
  NAND2_X2 U421 ( .A1(n1324), .A2(n1143), .ZN(n1353) );
  NAND2_X2 U422 ( .A1(n1354), .A2(n1143), .ZN(n1352) );
  NAND2_X2 U423 ( .A1(n1355), .A2(n1356), .ZN(B[24]) );
  MUX2_X1 U424 ( .A(n1357), .B(n1358), .S(n1137), .Z(n1356) );
  NAND2_X2 U425 ( .A1(n1153), .A2(n1324), .ZN(n1358) );
  NAND2_X2 U426 ( .A1(n1359), .A2(n1360), .ZN(n1324) );
  MUX2_X1 U427 ( .A(n1361), .B(n1362), .S(n1130), .Z(n1360) );
  NAND2_X2 U428 ( .A1(n1121), .A2(n1300), .ZN(n1362) );
  NAND2_X2 U429 ( .A1(n1120), .A2(n1231), .ZN(n1361) );
  MUX2_X1 U430 ( .A(n1363), .B(n1364), .S(n1130), .Z(n1359) );
  NAND2_X2 U431 ( .A1(n1304), .A2(n1109), .ZN(n1364) );
  NAND2_X2 U432 ( .A1(n1227), .A2(n1109), .ZN(n1363) );
  NAND2_X2 U433 ( .A1(n1153), .A2(n1354), .ZN(n1357) );
  MUX2_X1 U434 ( .A(n1365), .B(n1366), .S(n1137), .Z(n1355) );
  NAND2_X2 U435 ( .A1(n1339), .A2(n1143), .ZN(n1366) );
  NAND2_X2 U436 ( .A1(n1367), .A2(n1143), .ZN(n1365) );
  NAND2_X2 U437 ( .A1(n1368), .A2(n1369), .ZN(B[23]) );
  MUX2_X1 U438 ( .A(n1370), .B(n1371), .S(n1137), .Z(n1369) );
  NAND2_X2 U439 ( .A1(n1153), .A2(n1339), .ZN(n1371) );
  NAND2_X2 U440 ( .A1(n1372), .A2(n1373), .ZN(n1339) );
  MUX2_X1 U441 ( .A(n1374), .B(n1375), .S(n1130), .Z(n1373) );
  NAND2_X2 U442 ( .A1(n1120), .A2(n1317), .ZN(n1375) );
  NAND2_X2 U443 ( .A1(n1120), .A2(n1248), .ZN(n1374) );
  MUX2_X1 U444 ( .A(n1376), .B(n1377), .S(n1130), .Z(n1372) );
  NAND2_X2 U445 ( .A1(n1321), .A2(n1109), .ZN(n1377) );
  NAND2_X2 U446 ( .A1(n1244), .A2(n1109), .ZN(n1376) );
  NAND2_X2 U447 ( .A1(n1153), .A2(n1367), .ZN(n1370) );
  MUX2_X1 U448 ( .A(n1378), .B(n1379), .S(n1137), .Z(n1368) );
  NAND2_X2 U449 ( .A1(n1354), .A2(n1143), .ZN(n1379) );
  NAND2_X2 U450 ( .A1(n1380), .A2(n1143), .ZN(n1378) );
  NAND2_X2 U451 ( .A1(n1381), .A2(n1382), .ZN(B[22]) );
  MUX2_X1 U452 ( .A(n1383), .B(n1384), .S(n1137), .Z(n1382) );
  NAND2_X2 U453 ( .A1(n1152), .A2(n1354), .ZN(n1384) );
  NAND2_X2 U454 ( .A1(n1385), .A2(n1386), .ZN(n1354) );
  MUX2_X1 U455 ( .A(n1387), .B(n1388), .S(n1130), .Z(n1386) );
  NAND2_X2 U456 ( .A1(n1120), .A2(n1197), .ZN(n1388) );
  NAND2_X2 U457 ( .A1(n1120), .A2(n1198), .ZN(n1387) );
  MUX2_X1 U458 ( .A(n1389), .B(n1390), .S(n1130), .Z(n1385) );
  NAND2_X2 U459 ( .A1(n1193), .A2(n1109), .ZN(n1390) );
  NAND2_X2 U460 ( .A1(n1194), .A2(n1109), .ZN(n1389) );
  NAND2_X2 U461 ( .A1(n1152), .A2(n1380), .ZN(n1383) );
  MUX2_X1 U462 ( .A(n1391), .B(n1392), .S(n1137), .Z(n1381) );
  NAND2_X2 U463 ( .A1(n1367), .A2(n1143), .ZN(n1392) );
  NAND2_X2 U464 ( .A1(n1393), .A2(n1143), .ZN(n1391) );
  NAND2_X2 U465 ( .A1(n1394), .A2(n1395), .ZN(B[21]) );
  MUX2_X1 U466 ( .A(n1396), .B(n1397), .S(n1138), .Z(n1395) );
  NAND2_X2 U467 ( .A1(n1152), .A2(n1367), .ZN(n1397) );
  NAND2_X2 U468 ( .A1(n1398), .A2(n1399), .ZN(n1367) );
  MUX2_X1 U469 ( .A(n1400), .B(n1401), .S(n1131), .Z(n1399) );
  NAND2_X2 U470 ( .A1(n1119), .A2(n1214), .ZN(n1401) );
  NAND2_X2 U471 ( .A1(n1119), .A2(n1215), .ZN(n1400) );
  MUX2_X1 U472 ( .A(n1402), .B(n1403), .S(n1131), .Z(n1398) );
  NAND2_X2 U473 ( .A1(n1210), .A2(n1109), .ZN(n1403) );
  NAND2_X2 U474 ( .A1(n1211), .A2(n1109), .ZN(n1402) );
  NAND2_X2 U475 ( .A1(n1152), .A2(n1393), .ZN(n1396) );
  MUX2_X1 U476 ( .A(n1404), .B(n1405), .S(n1138), .Z(n1394) );
  NAND2_X2 U477 ( .A1(n1380), .A2(n1143), .ZN(n1405) );
  NAND2_X2 U478 ( .A1(n1406), .A2(n1143), .ZN(n1404) );
  NAND2_X2 U479 ( .A1(n1407), .A2(n1408), .ZN(B[20]) );
  MUX2_X1 U480 ( .A(n1409), .B(n1410), .S(n1138), .Z(n1408) );
  NAND2_X2 U481 ( .A1(n1152), .A2(n1380), .ZN(n1410) );
  NAND2_X2 U482 ( .A1(n1411), .A2(n1412), .ZN(n1380) );
  MUX2_X1 U483 ( .A(n1413), .B(n1414), .S(n1131), .Z(n1412) );
  NAND2_X2 U484 ( .A1(n1119), .A2(n1231), .ZN(n1414) );
  NAND2_X2 U485 ( .A1(n1119), .A2(n1232), .ZN(n1413) );
  MUX2_X1 U486 ( .A(n1415), .B(n1416), .S(n1131), .Z(n1411) );
  NAND2_X2 U487 ( .A1(n1227), .A2(n1109), .ZN(n1416) );
  NAND2_X2 U488 ( .A1(n1228), .A2(n1109), .ZN(n1415) );
  NAND2_X2 U489 ( .A1(n1151), .A2(n1406), .ZN(n1409) );
  MUX2_X1 U490 ( .A(n1417), .B(n1418), .S(n1138), .Z(n1407) );
  NAND2_X2 U491 ( .A1(n1393), .A2(n1143), .ZN(n1418) );
  NAND2_X2 U492 ( .A1(n1419), .A2(n1143), .ZN(n1417) );
  NAND2_X2 U493 ( .A1(n1420), .A2(n1421), .ZN(B[1]) );
  MUX2_X1 U494 ( .A(n1422), .B(n1423), .S(n1138), .Z(n1421) );
  NAND2_X2 U495 ( .A1(n1151), .A2(n1235), .ZN(n1423) );
  NAND2_X2 U496 ( .A1(n1424), .A2(n1425), .ZN(n1235) );
  MUX2_X1 U497 ( .A(n1426), .B(n1427), .S(n1131), .Z(n1425) );
  NAND2_X2 U498 ( .A1(n1119), .A2(n1211), .ZN(n1427) );
  NAND2_X2 U499 ( .A1(n1118), .A2(n1428), .ZN(n1426) );
  MUX2_X1 U500 ( .A(n1429), .B(n1430), .S(n1131), .Z(n1424) );
  NAND2_X2 U501 ( .A1(n1215), .A2(n1108), .ZN(n1430) );
  NAND2_X2 U502 ( .A1(n1431), .A2(n1108), .ZN(n1429) );
  NAND2_X2 U503 ( .A1(n1151), .A2(n1257), .ZN(n1422) );
  MUX2_X1 U504 ( .A(n1432), .B(n1433), .S(n1138), .Z(n1420) );
  NAND2_X2 U505 ( .A1(n1252), .A2(n1142), .ZN(n1433) );
  NAND2_X2 U506 ( .A1(n1261), .A2(n1142), .ZN(n1432) );
  NAND2_X2 U507 ( .A1(n1434), .A2(n1435), .ZN(B[19]) );
  MUX2_X1 U508 ( .A(n1436), .B(n1437), .S(n1138), .Z(n1435) );
  NAND2_X2 U509 ( .A1(n1151), .A2(n1393), .ZN(n1437) );
  NAND2_X2 U510 ( .A1(n1438), .A2(n1439), .ZN(n1393) );
  MUX2_X1 U511 ( .A(n1440), .B(n1441), .S(n1131), .Z(n1439) );
  NAND2_X2 U512 ( .A1(n1118), .A2(n1248), .ZN(n1441) );
  NAND2_X2 U513 ( .A1(n1118), .A2(n1249), .ZN(n1440) );
  MUX2_X1 U514 ( .A(n1442), .B(n1443), .S(n1131), .Z(n1438) );
  NAND2_X2 U515 ( .A1(n1244), .A2(n1108), .ZN(n1443) );
  NAND2_X2 U516 ( .A1(n1245), .A2(n1108), .ZN(n1442) );
  NAND2_X2 U517 ( .A1(n1151), .A2(n1419), .ZN(n1436) );
  MUX2_X1 U518 ( .A(n1444), .B(n1445), .S(n1138), .Z(n1434) );
  NAND2_X2 U519 ( .A1(n1406), .A2(n1142), .ZN(n1445) );
  NAND2_X2 U520 ( .A1(n1446), .A2(n1142), .ZN(n1444) );
  NAND2_X2 U521 ( .A1(n1447), .A2(n1448), .ZN(B[18]) );
  MUX2_X1 U522 ( .A(n1449), .B(n1450), .S(n1138), .Z(n1448) );
  NAND2_X2 U523 ( .A1(n1150), .A2(n1406), .ZN(n1450) );
  NAND2_X2 U524 ( .A1(n1451), .A2(n1452), .ZN(n1406) );
  MUX2_X1 U525 ( .A(n1453), .B(n1454), .S(n1131), .Z(n1452) );
  NAND2_X2 U526 ( .A1(n1118), .A2(n1198), .ZN(n1454) );
  INV_X2 U527 ( .A(n1455), .ZN(n1198) );
  MUX2_X1 U528 ( .A(n1456), .B(n1457), .S(n1126), .Z(n1455) );
  NAND2_X2 U529 ( .A1(n1118), .A2(n1281), .ZN(n1453) );
  MUX2_X1 U530 ( .A(n1458), .B(n1459), .S(n1131), .Z(n1451) );
  NAND2_X2 U531 ( .A1(n1194), .A2(n1108), .ZN(n1459) );
  INV_X2 U532 ( .A(n1460), .ZN(n1194) );
  MUX2_X1 U533 ( .A(n1461), .B(n1462), .S(n1126), .Z(n1460) );
  NAND2_X2 U534 ( .A1(n1278), .A2(n1108), .ZN(n1458) );
  NAND2_X2 U535 ( .A1(n1150), .A2(n1446), .ZN(n1449) );
  MUX2_X1 U536 ( .A(n1463), .B(n1464), .S(n1138), .Z(n1447) );
  NAND2_X2 U537 ( .A1(n1419), .A2(n1142), .ZN(n1464) );
  NAND2_X2 U538 ( .A1(n1465), .A2(n1142), .ZN(n1463) );
  NAND2_X2 U539 ( .A1(n1466), .A2(n1467), .ZN(B[17]) );
  MUX2_X1 U540 ( .A(n1468), .B(n1469), .S(n1138), .Z(n1467) );
  NAND2_X2 U541 ( .A1(n1150), .A2(n1419), .ZN(n1469) );
  NAND2_X2 U542 ( .A1(n1470), .A2(n1471), .ZN(n1419) );
  MUX2_X1 U543 ( .A(n1472), .B(n1473), .S(n1131), .Z(n1471) );
  NAND2_X2 U544 ( .A1(n1117), .A2(n1215), .ZN(n1473) );
  INV_X2 U545 ( .A(n1474), .ZN(n1215) );
  MUX2_X1 U546 ( .A(n1475), .B(n1476), .S(n1126), .Z(n1474) );
  NAND2_X2 U547 ( .A1(n1117), .A2(n1431), .ZN(n1472) );
  MUX2_X1 U548 ( .A(n1477), .B(n1478), .S(n1131), .Z(n1470) );
  NAND2_X2 U549 ( .A1(n1211), .A2(n1108), .ZN(n1478) );
  INV_X2 U550 ( .A(n1479), .ZN(n1211) );
  MUX2_X1 U551 ( .A(n1480), .B(n1481), .S(n1126), .Z(n1479) );
  NAND2_X2 U552 ( .A1(n1428), .A2(n1108), .ZN(n1477) );
  NAND2_X2 U553 ( .A1(n1150), .A2(n1465), .ZN(n1468) );
  MUX2_X1 U554 ( .A(n1482), .B(n1483), .S(n1138), .Z(n1466) );
  NAND2_X2 U555 ( .A1(n1446), .A2(n1142), .ZN(n1483) );
  NAND2_X2 U556 ( .A1(n1484), .A2(n1142), .ZN(n1482) );
  NAND2_X2 U557 ( .A1(n1485), .A2(n1486), .ZN(B[16]) );
  MUX2_X1 U558 ( .A(n1487), .B(n1488), .S(n1139), .Z(n1486) );
  NAND2_X2 U559 ( .A1(n1150), .A2(n1446), .ZN(n1488) );
  NAND2_X2 U560 ( .A1(n1489), .A2(n1490), .ZN(n1446) );
  MUX2_X1 U561 ( .A(n1491), .B(n1492), .S(n1132), .Z(n1490) );
  NAND2_X2 U562 ( .A1(n1117), .A2(n1232), .ZN(n1492) );
  NAND2_X2 U563 ( .A1(n1117), .A2(n1303), .ZN(n1491) );
  MUX2_X1 U564 ( .A(n1493), .B(n1494), .S(n1132), .Z(n1489) );
  NAND2_X2 U565 ( .A1(n1228), .A2(n1108), .ZN(n1494) );
  NAND2_X2 U566 ( .A1(n1299), .A2(n1108), .ZN(n1493) );
  NAND2_X2 U567 ( .A1(n1149), .A2(n1484), .ZN(n1487) );
  MUX2_X1 U568 ( .A(n1495), .B(n1496), .S(n1139), .Z(n1485) );
  NAND2_X2 U569 ( .A1(n1465), .A2(n1142), .ZN(n1496) );
  NAND2_X2 U570 ( .A1(n1497), .A2(n1142), .ZN(n1495) );
  NAND2_X2 U571 ( .A1(n1498), .A2(n1499), .ZN(B[15]) );
  MUX2_X1 U572 ( .A(n1500), .B(n1501), .S(n1139), .Z(n1499) );
  NAND2_X2 U573 ( .A1(n1149), .A2(n1465), .ZN(n1501) );
  NAND2_X2 U574 ( .A1(n1502), .A2(n1503), .ZN(n1465) );
  MUX2_X1 U575 ( .A(n1504), .B(n1505), .S(n1132), .Z(n1503) );
  NAND2_X2 U576 ( .A1(n1117), .A2(n1249), .ZN(n1505) );
  NAND2_X2 U577 ( .A1(n1116), .A2(n1320), .ZN(n1504) );
  MUX2_X1 U578 ( .A(n1506), .B(n1507), .S(n1132), .Z(n1502) );
  NAND2_X2 U579 ( .A1(n1245), .A2(n1108), .ZN(n1507) );
  NAND2_X2 U580 ( .A1(n1316), .A2(n1108), .ZN(n1506) );
  NAND2_X2 U581 ( .A1(n1149), .A2(n1497), .ZN(n1500) );
  MUX2_X1 U582 ( .A(n1508), .B(n1509), .S(n1139), .Z(n1498) );
  NAND2_X2 U583 ( .A1(n1484), .A2(n1142), .ZN(n1509) );
  NAND2_X2 U584 ( .A1(n1510), .A2(n1142), .ZN(n1508) );
  NAND2_X2 U585 ( .A1(n1511), .A2(n1512), .ZN(B[14]) );
  MUX2_X1 U586 ( .A(n1513), .B(n1514), .S(n1139), .Z(n1512) );
  NAND2_X2 U587 ( .A1(n1149), .A2(n1484), .ZN(n1514) );
  NAND2_X2 U588 ( .A1(n1515), .A2(n1516), .ZN(n1484) );
  MUX2_X1 U589 ( .A(n1517), .B(n1518), .S(n1132), .Z(n1516) );
  NAND2_X2 U590 ( .A1(n1116), .A2(n1281), .ZN(n1518) );
  NAND2_X2 U591 ( .A1(n1116), .A2(n1336), .ZN(n1517) );
  MUX2_X1 U592 ( .A(n1519), .B(n1520), .S(n1132), .Z(n1515) );
  NAND2_X2 U593 ( .A1(n1278), .A2(n1107), .ZN(n1520) );
  NAND2_X2 U594 ( .A1(n1333), .A2(n1107), .ZN(n1519) );
  NAND2_X2 U595 ( .A1(n1149), .A2(n1510), .ZN(n1513) );
  MUX2_X1 U596 ( .A(n1521), .B(n1522), .S(n1139), .Z(n1511) );
  NAND2_X2 U597 ( .A1(n1497), .A2(n1141), .ZN(n1522) );
  NAND2_X2 U598 ( .A1(n1523), .A2(n1141), .ZN(n1521) );
  NAND2_X2 U599 ( .A1(n1524), .A2(n1525), .ZN(B[13]) );
  MUX2_X1 U600 ( .A(n1526), .B(n1527), .S(n1139), .Z(n1525) );
  NAND2_X2 U601 ( .A1(n1148), .A2(n1497), .ZN(n1527) );
  NAND2_X2 U602 ( .A1(n1528), .A2(n1529), .ZN(n1497) );
  MUX2_X1 U603 ( .A(n1530), .B(n1531), .S(n1132), .Z(n1529) );
  NAND2_X2 U604 ( .A1(n1116), .A2(n1431), .ZN(n1531) );
  NAND2_X2 U605 ( .A1(n1116), .A2(n1351), .ZN(n1530) );
  MUX2_X1 U606 ( .A(n1532), .B(n1533), .S(n1132), .Z(n1528) );
  NAND2_X2 U607 ( .A1(n1428), .A2(n1107), .ZN(n1533) );
  NAND2_X2 U608 ( .A1(n1348), .A2(n1107), .ZN(n1532) );
  NAND2_X2 U609 ( .A1(n1148), .A2(n1523), .ZN(n1526) );
  MUX2_X1 U610 ( .A(n1534), .B(n1535), .S(n1139), .Z(n1524) );
  NAND2_X2 U611 ( .A1(n1510), .A2(n1141), .ZN(n1535) );
  NAND2_X2 U612 ( .A1(n1536), .A2(n1141), .ZN(n1534) );
  NAND2_X2 U613 ( .A1(n1537), .A2(n1538), .ZN(B[12]) );
  MUX2_X1 U614 ( .A(n1539), .B(n1540), .S(n1139), .Z(n1538) );
  NAND2_X2 U615 ( .A1(n1148), .A2(n1510), .ZN(n1540) );
  NAND2_X2 U616 ( .A1(n1541), .A2(n1542), .ZN(n1510) );
  MUX2_X1 U617 ( .A(n1543), .B(n1544), .S(n1132), .Z(n1542) );
  NAND2_X2 U618 ( .A1(n1115), .A2(n1303), .ZN(n1544) );
  NAND2_X2 U619 ( .A1(n1115), .A2(n1304), .ZN(n1543) );
  MUX2_X1 U620 ( .A(n1545), .B(n1546), .S(n1132), .Z(n1541) );
  NAND2_X2 U621 ( .A1(n1299), .A2(n1107), .ZN(n1546) );
  NAND2_X2 U622 ( .A1(n1300), .A2(n1107), .ZN(n1545) );
  NAND2_X2 U623 ( .A1(n1148), .A2(n1536), .ZN(n1539) );
  MUX2_X1 U624 ( .A(n1547), .B(n1548), .S(n1139), .Z(n1537) );
  NAND2_X2 U625 ( .A1(n1523), .A2(n1141), .ZN(n1548) );
  NAND2_X2 U626 ( .A1(n1165), .A2(n1141), .ZN(n1547) );
  NAND2_X2 U627 ( .A1(n1549), .A2(n1550), .ZN(B[11]) );
  MUX2_X1 U628 ( .A(n1551), .B(n1552), .S(n1139), .Z(n1550) );
  NAND2_X2 U629 ( .A1(n1148), .A2(n1523), .ZN(n1552) );
  NAND2_X2 U630 ( .A1(n1553), .A2(n1554), .ZN(n1523) );
  MUX2_X1 U631 ( .A(n1555), .B(n1556), .S(n1132), .Z(n1554) );
  NAND2_X2 U632 ( .A1(n1115), .A2(n1320), .ZN(n1556) );
  NAND2_X2 U633 ( .A1(n1115), .A2(n1321), .ZN(n1555) );
  MUX2_X1 U634 ( .A(n1557), .B(n1558), .S(n1132), .Z(n1553) );
  NAND2_X2 U635 ( .A1(n1316), .A2(n1107), .ZN(n1558) );
  NAND2_X2 U636 ( .A1(n1317), .A2(n1107), .ZN(n1557) );
  NAND2_X2 U637 ( .A1(n1147), .A2(n1165), .ZN(n1551) );
  MUX2_X1 U638 ( .A(n1559), .B(n1560), .S(n1139), .Z(n1549) );
  NAND2_X2 U639 ( .A1(n1536), .A2(n1141), .ZN(n1560) );
  NAND2_X2 U640 ( .A1(n1169), .A2(n1141), .ZN(n1559) );
  NAND2_X2 U641 ( .A1(n1561), .A2(n1562), .ZN(B[10]) );
  MUX2_X1 U642 ( .A(n1563), .B(n1564), .S(n1140), .Z(n1562) );
  NAND2_X2 U643 ( .A1(n1147), .A2(n1536), .ZN(n1564) );
  NAND2_X2 U644 ( .A1(n1565), .A2(n1566), .ZN(n1536) );
  MUX2_X1 U645 ( .A(n1567), .B(n1568), .S(n1133), .Z(n1566) );
  NAND2_X2 U646 ( .A1(n1115), .A2(n1336), .ZN(n1568) );
  NAND2_X2 U647 ( .A1(n1114), .A2(n1193), .ZN(n1567) );
  INV_X2 U648 ( .A(n1569), .ZN(n1193) );
  MUX2_X1 U649 ( .A(n1570), .B(n1571), .S(n1126), .Z(n1569) );
  MUX2_X1 U650 ( .A(n1572), .B(n1573), .S(n1133), .Z(n1565) );
  NAND2_X2 U651 ( .A1(n1333), .A2(n1107), .ZN(n1573) );
  NAND2_X2 U652 ( .A1(n1197), .A2(n1107), .ZN(n1572) );
  INV_X2 U653 ( .A(n1574), .ZN(n1197) );
  MUX2_X1 U654 ( .A(n1575), .B(n1576), .S(n1126), .Z(n1574) );
  NAND2_X2 U655 ( .A1(n1147), .A2(n1169), .ZN(n1563) );
  NAND2_X2 U656 ( .A1(n1577), .A2(n1578), .ZN(n1169) );
  MUX2_X1 U657 ( .A(n1579), .B(n1580), .S(n1133), .Z(n1578) );
  NAND2_X2 U658 ( .A1(n1114), .A2(n1304), .ZN(n1580) );
  INV_X2 U659 ( .A(n1581), .ZN(n1304) );
  MUX2_X1 U660 ( .A(n1582), .B(n1583), .S(n1126), .Z(n1581) );
  NAND2_X2 U661 ( .A1(n1114), .A2(n1227), .ZN(n1579) );
  INV_X2 U662 ( .A(n1584), .ZN(n1227) );
  MUX2_X1 U663 ( .A(n1585), .B(n1586), .S(n1126), .Z(n1584) );
  MUX2_X1 U664 ( .A(n1587), .B(n1588), .S(n1133), .Z(n1577) );
  NAND2_X2 U665 ( .A1(n1300), .A2(n1107), .ZN(n1588) );
  INV_X2 U666 ( .A(n1589), .ZN(n1300) );
  MUX2_X1 U667 ( .A(n1590), .B(n1591), .S(n1126), .Z(n1589) );
  NAND2_X2 U668 ( .A1(n1231), .A2(n1107), .ZN(n1587) );
  INV_X2 U669 ( .A(n1592), .ZN(n1231) );
  MUX2_X1 U670 ( .A(n1593), .B(n1594), .S(n1126), .Z(n1592) );
  MUX2_X1 U671 ( .A(n1595), .B(n1596), .S(n1140), .Z(n1561) );
  NAND2_X2 U672 ( .A1(n1165), .A2(n1141), .ZN(n1596) );
  NAND2_X2 U673 ( .A1(n1597), .A2(n1598), .ZN(n1165) );
  MUX2_X1 U674 ( .A(n1599), .B(n1600), .S(n1133), .Z(n1598) );
  NAND2_X2 U675 ( .A1(n1114), .A2(n1351), .ZN(n1600) );
  NAND2_X2 U676 ( .A1(n1114), .A2(n1210), .ZN(n1599) );
  INV_X2 U677 ( .A(n1601), .ZN(n1210) );
  MUX2_X1 U678 ( .A(n1602), .B(n1603), .S(n1126), .Z(n1601) );
  MUX2_X1 U679 ( .A(n1604), .B(n1605), .S(n1133), .Z(n1597) );
  NAND2_X2 U680 ( .A1(n1348), .A2(n1106), .ZN(n1605) );
  NAND2_X2 U681 ( .A1(n1214), .A2(n1106), .ZN(n1604) );
  INV_X2 U682 ( .A(n1606), .ZN(n1214) );
  MUX2_X1 U683 ( .A(n1607), .B(n1608), .S(n1126), .Z(n1606) );
  NAND2_X2 U684 ( .A1(n1166), .A2(n1141), .ZN(n1595) );
  NAND2_X2 U685 ( .A1(n1609), .A2(n1610), .ZN(n1166) );
  MUX2_X1 U686 ( .A(n1611), .B(n1612), .S(n1133), .Z(n1610) );
  NAND2_X2 U687 ( .A1(n1113), .A2(n1321), .ZN(n1612) );
  INV_X2 U688 ( .A(n1613), .ZN(n1321) );
  MUX2_X1 U689 ( .A(n1614), .B(n1615), .S(n1127), .Z(n1613) );
  NAND2_X2 U690 ( .A1(n1113), .A2(n1244), .ZN(n1611) );
  INV_X2 U691 ( .A(n1616), .ZN(n1244) );
  MUX2_X1 U692 ( .A(n1617), .B(n1618), .S(n1127), .Z(n1616) );
  MUX2_X1 U693 ( .A(n1619), .B(n1620), .S(n1133), .Z(n1609) );
  NAND2_X2 U694 ( .A1(n1317), .A2(n1106), .ZN(n1620) );
  INV_X2 U695 ( .A(n1621), .ZN(n1317) );
  MUX2_X1 U696 ( .A(n1622), .B(n1623), .S(n1127), .Z(n1621) );
  NAND2_X2 U697 ( .A1(n1248), .A2(n1106), .ZN(n1619) );
  INV_X2 U698 ( .A(n1624), .ZN(n1248) );
  MUX2_X1 U699 ( .A(n1625), .B(n1626), .S(n1127), .Z(n1624) );
  NAND2_X2 U700 ( .A1(n1627), .A2(n1628), .ZN(B[0]) );
  MUX2_X1 U701 ( .A(n1629), .B(n1630), .S(n1140), .Z(n1628) );
  NAND2_X2 U702 ( .A1(n1147), .A2(n1252), .ZN(n1630) );
  NAND2_X2 U703 ( .A1(n1631), .A2(n1632), .ZN(n1252) );
  MUX2_X1 U704 ( .A(n1633), .B(n1634), .S(n1133), .Z(n1632) );
  NAND2_X2 U705 ( .A1(n1113), .A2(n1228), .ZN(n1634) );
  INV_X2 U706 ( .A(n1635), .ZN(n1228) );
  MUX2_X1 U707 ( .A(n1591), .B(n1582), .S(n1127), .Z(n1635) );
  INV_X2 U708 ( .A(A[23]), .ZN(n1591) );
  NAND2_X2 U709 ( .A1(n1113), .A2(n1299), .ZN(n1633) );
  INV_X2 U710 ( .A(n1636), .ZN(n1299) );
  MUX2_X1 U711 ( .A(n1594), .B(n1585), .S(n1127), .Z(n1636) );
  MUX2_X1 U712 ( .A(n1637), .B(n1638), .S(n1133), .Z(n1631) );
  NAND2_X2 U713 ( .A1(n1232), .A2(n1106), .ZN(n1638) );
  INV_X2 U714 ( .A(n1639), .ZN(n1232) );
  MUX2_X1 U715 ( .A(n1583), .B(n1590), .S(n1127), .Z(n1639) );
  NAND2_X2 U716 ( .A1(n1303), .A2(n1106), .ZN(n1637) );
  INV_X2 U717 ( .A(n1640), .ZN(n1303) );
  MUX2_X1 U718 ( .A(n1586), .B(n1593), .S(n1127), .Z(n1640) );
  INV_X2 U719 ( .A(A[3]), .ZN(n1586) );
  NAND2_X2 U720 ( .A1(n1147), .A2(n1261), .ZN(n1629) );
  NAND2_X2 U721 ( .A1(n1641), .A2(n1642), .ZN(n1261) );
  MUX2_X1 U722 ( .A(n1643), .B(n1644), .S(n1133), .Z(n1642) );
  NAND2_X2 U723 ( .A1(n1113), .A2(n1278), .ZN(n1644) );
  INV_X2 U724 ( .A(n1645), .ZN(n1278) );
  MUX2_X1 U725 ( .A(n1576), .B(n1570), .S(n1127), .Z(n1645) );
  NAND2_X2 U726 ( .A1(n1112), .A2(n1333), .ZN(n1643) );
  INV_X2 U727 ( .A(n1646), .ZN(n1333) );
  MUX2_X1 U728 ( .A(n1457), .B(n1461), .S(n1127), .Z(n1646) );
  MUX2_X1 U729 ( .A(n1647), .B(n1648), .S(n1133), .Z(n1641) );
  NAND2_X2 U730 ( .A1(n1281), .A2(n1106), .ZN(n1648) );
  INV_X2 U731 ( .A(n1649), .ZN(n1281) );
  MUX2_X1 U732 ( .A(n1571), .B(n1575), .S(n1127), .Z(n1649) );
  NAND2_X2 U733 ( .A1(n1336), .A2(n1106), .ZN(n1647) );
  INV_X2 U734 ( .A(n1650), .ZN(n1336) );
  MUX2_X1 U735 ( .A(n1462), .B(n1456), .S(n1127), .Z(n1650) );
  MUX2_X1 U736 ( .A(n1651), .B(n1652), .S(n1140), .Z(n1627) );
  NAND2_X2 U737 ( .A1(n1257), .A2(n1141), .ZN(n1652) );
  NAND2_X2 U738 ( .A1(n1653), .A2(n1654), .ZN(n1257) );
  MUX2_X1 U739 ( .A(n1655), .B(n1656), .S(n1134), .Z(n1654) );
  NAND2_X2 U740 ( .A1(n1112), .A2(n1245), .ZN(n1656) );
  INV_X2 U741 ( .A(n1657), .ZN(n1245) );
  MUX2_X1 U742 ( .A(n1623), .B(n1614), .S(n1128), .Z(n1657) );
  NAND2_X2 U743 ( .A1(n1112), .A2(n1316), .ZN(n1655) );
  INV_X2 U744 ( .A(n1658), .ZN(n1316) );
  MUX2_X1 U745 ( .A(n1626), .B(n1617), .S(n1128), .Z(n1658) );
  MUX2_X1 U746 ( .A(n1659), .B(n1660), .S(n1134), .Z(n1653) );
  NAND2_X2 U747 ( .A1(n1249), .A2(n1106), .ZN(n1660) );
  INV_X2 U748 ( .A(n1661), .ZN(n1249) );
  MUX2_X1 U749 ( .A(n1615), .B(n1622), .S(n1128), .Z(n1661) );
  NAND2_X2 U750 ( .A1(n1320), .A2(n1106), .ZN(n1659) );
  INV_X2 U751 ( .A(n1662), .ZN(n1320) );
  MUX2_X1 U752 ( .A(n1618), .B(n1625), .S(n1128), .Z(n1662) );
  NAND2_X2 U753 ( .A1(n1258), .A2(n1141), .ZN(n1651) );
  NAND2_X2 U754 ( .A1(n1663), .A2(n1664), .ZN(n1258) );
  MUX2_X1 U755 ( .A(n1665), .B(n1666), .S(n1134), .Z(n1664) );
  NAND2_X2 U756 ( .A1(n1112), .A2(n1428), .ZN(n1666) );
  INV_X2 U757 ( .A(n1667), .ZN(n1428) );
  MUX2_X1 U758 ( .A(n1608), .B(n1602), .S(n1128), .Z(n1667) );
  NAND2_X2 U759 ( .A1(n1112), .A2(n1348), .ZN(n1665) );
  INV_X2 U760 ( .A(n1668), .ZN(n1348) );
  MUX2_X1 U761 ( .A(n1476), .B(n1480), .S(n1128), .Z(n1668) );
  MUX2_X1 U762 ( .A(n1669), .B(n1670), .S(n1134), .Z(n1663) );
  NAND2_X2 U763 ( .A1(n1431), .A2(n1106), .ZN(n1670) );
  INV_X2 U764 ( .A(n1671), .ZN(n1431) );
  MUX2_X1 U765 ( .A(n1603), .B(n1607), .S(n1128), .Z(n1671) );
  NAND2_X2 U766 ( .A1(n1351), .A2(n1106), .ZN(n1669) );
  INV_X2 U767 ( .A(n1672), .ZN(n1351) );
  MUX2_X1 U768 ( .A(n1481), .B(n1475), .S(n1128), .Z(n1672) );
endmodule


module Xi_core_DW_sra_1 ( A, SH, B, SH_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  INV_X1 U170 ( .A(A[24]), .ZN(n1409) );
  INV_X1 U171 ( .A(A[26]), .ZN(n1534) );
  INV_X4 U172 ( .A(n1130), .ZN(n1119) );
  BUF_X4 U173 ( .A(n1133), .Z(n1130) );
  NAND2_X1 U174 ( .A1(n1121), .A2(n1191), .ZN(n1188) );
  NAND2_X1 U175 ( .A1(n1121), .A2(n1224), .ZN(n1223) );
  NAND2_X1 U176 ( .A1(n1121), .A2(n1242), .ZN(n1239) );
  NAND2_X1 U177 ( .A1(n1121), .A2(n1194), .ZN(n1262) );
  NAND2_X1 U178 ( .A1(n1121), .A2(n1195), .ZN(n1261) );
  NAND2_X1 U179 ( .A1(n1121), .A2(n1207), .ZN(n1347) );
  NAND2_X1 U180 ( .A1(n1139), .A2(n1445), .ZN(n1470) );
  NAND2_X1 U181 ( .A1(n1140), .A2(n1445), .ZN(n1459) );
  NAND2_X1 U182 ( .A1(n1445), .A2(n1138), .ZN(n1455) );
  NAND2_X1 U183 ( .A1(n1445), .A2(n1137), .ZN(n1443) );
  NAND2_X1 U184 ( .A1(n1120), .A2(n1463), .ZN(n1510) );
  NAND2_X1 U185 ( .A1(n1120), .A2(n1211), .ZN(n1407) );
  NAND2_X1 U186 ( .A1(n1120), .A2(n1245), .ZN(n1431) );
  NAND2_X1 U187 ( .A1(n1120), .A2(n1228), .ZN(n1420) );
  NAND2_X1 U188 ( .A1(n1120), .A2(n1441), .ZN(n1486) );
  NAND2_X1 U189 ( .A1(n1120), .A2(n1194), .ZN(n1395) );
  NAND2_X1 U190 ( .A1(n1120), .A2(n1419), .ZN(n1464) );
  NAND2_X1 U191 ( .A1(n1120), .A2(n1374), .ZN(n1453) );
  NAND2_X1 U192 ( .A1(n1120), .A2(n1268), .ZN(n1442) );
  NAND2_X1 U193 ( .A1(n1120), .A2(n1430), .ZN(n1473) );
  INV_X1 U194 ( .A(A[28]), .ZN(n1502) );
  INV_X1 U195 ( .A(A[4]), .ZN(n1587) );
  INV_X1 U196 ( .A(A[30]), .ZN(n1527) );
  INV_X1 U197 ( .A(A[22]), .ZN(n1530) );
  INV_X1 U198 ( .A(A[25]), .ZN(n1397) );
  INV_X1 U199 ( .A(A[29]), .ZN(n1491) );
  INV_X1 U200 ( .A(A[27]), .ZN(n1518) );
  INV_X1 U201 ( .A(A[21]), .ZN(n1494) );
  NAND2_X1 U202 ( .A1(n1147), .A2(\A[31] ), .ZN(n1280) );
  OAI21_X1 U203 ( .B1(n1253), .B2(n1111), .A(n1316), .ZN(n1293) );
  OAI21_X1 U204 ( .B1(n1253), .B2(n1111), .A(n1307), .ZN(n1283) );
  OAI21_X1 U205 ( .B1(n1253), .B2(n1111), .A(n1298), .ZN(n1275) );
  NAND2_X1 U206 ( .A1(n1152), .A2(\A[31] ), .ZN(n1251) );
  OAI21_X1 U207 ( .B1(n1253), .B2(n1111), .A(n1288), .ZN(n1254) );
  NAND2_X1 U208 ( .A1(n1120), .A2(\A[31] ), .ZN(n1487) );
  NAND2_X1 U209 ( .A1(n1120), .A2(\A[31] ), .ZN(n1474) );
  NAND2_X1 U210 ( .A1(n1119), .A2(\A[31] ), .ZN(n1511) );
  NAND2_X1 U211 ( .A1(n1119), .A2(\A[31] ), .ZN(n1498) );
  INV_X4 U212 ( .A(\A[31] ), .ZN(n1253) );
  INV_X1 U213 ( .A(A[6]), .ZN(n1559) );
  INV_X1 U214 ( .A(A[7]), .ZN(n1548) );
  INV_X1 U215 ( .A(A[5]), .ZN(n1572) );
  INV_X1 U216 ( .A(A[19]), .ZN(n1521) );
  INV_X1 U217 ( .A(A[18]), .ZN(n1537) );
  INV_X1 U218 ( .A(A[16]), .ZN(n1371) );
  INV_X1 U219 ( .A(A[13]), .ZN(n1493) );
  INV_X1 U220 ( .A(A[17]), .ZN(n1265) );
  INV_X1 U221 ( .A(A[15]), .ZN(n1513) );
  INV_X1 U222 ( .A(A[14]), .ZN(n1529) );
  INV_X1 U223 ( .A(A[20]), .ZN(n1505) );
  INV_X1 U224 ( .A(A[12]), .ZN(n1504) );
  INV_X1 U225 ( .A(A[9]), .ZN(n1264) );
  INV_X1 U226 ( .A(A[11]), .ZN(n1520) );
  INV_X1 U227 ( .A(A[8]), .ZN(n1370) );
  INV_X1 U228 ( .A(A[10]), .ZN(n1536) );
  INV_X1 U229 ( .A(n1112), .ZN(n1106) );
  INV_X1 U230 ( .A(n1112), .ZN(n1107) );
  INV_X1 U231 ( .A(n1112), .ZN(n1108) );
  INV_X1 U232 ( .A(n1112), .ZN(n1109) );
  CLKBUF_X3 U233 ( .A(n1115), .Z(n1110) );
  CLKBUF_X3 U234 ( .A(n1115), .Z(n1111) );
  CLKBUF_X3 U235 ( .A(n1115), .Z(n1112) );
  CLKBUF_X3 U236 ( .A(n1115), .Z(n1113) );
  CLKBUF_X3 U237 ( .A(n1115), .Z(n1114) );
  INV_X8 U238 ( .A(SH[4]), .ZN(n1115) );
  CLKBUF_X3 U239 ( .A(SH[3]), .Z(n1116) );
  CLKBUF_X3 U240 ( .A(SH[3]), .Z(n1117) );
  CLKBUF_X3 U241 ( .A(SH[3]), .Z(n1118) );
  INV_X1 U242 ( .A(n1130), .ZN(n1120) );
  INV_X1 U243 ( .A(n1130), .ZN(n1121) );
  INV_X1 U244 ( .A(n1130), .ZN(n1122) );
  CLKBUF_X3 U245 ( .A(n1133), .Z(n1123) );
  CLKBUF_X3 U246 ( .A(n1133), .Z(n1124) );
  CLKBUF_X3 U247 ( .A(n1133), .Z(n1125) );
  CLKBUF_X3 U248 ( .A(n1133), .Z(n1126) );
  CLKBUF_X3 U249 ( .A(n1133), .Z(n1127) );
  CLKBUF_X3 U250 ( .A(n1133), .Z(n1128) );
  CLKBUF_X3 U251 ( .A(n1133), .Z(n1129) );
  CLKBUF_X3 U252 ( .A(n1133), .Z(n1131) );
  CLKBUF_X3 U253 ( .A(n1133), .Z(n1132) );
  INV_X16 U254 ( .A(SH[2]), .ZN(n1133) );
  INV_X1 U255 ( .A(n1150), .ZN(n1134) );
  INV_X1 U256 ( .A(n1151), .ZN(n1135) );
  INV_X1 U257 ( .A(n1151), .ZN(n1136) );
  INV_X1 U258 ( .A(n1151), .ZN(n1137) );
  INV_X1 U259 ( .A(n1151), .ZN(n1138) );
  CLKBUF_X3 U260 ( .A(SH[1]), .Z(n1139) );
  CLKBUF_X3 U261 ( .A(SH[1]), .Z(n1140) );
  CLKBUF_X3 U262 ( .A(SH[1]), .Z(n1141) );
  CLKBUF_X3 U263 ( .A(SH[1]), .Z(n1142) );
  CLKBUF_X3 U264 ( .A(SH[1]), .Z(n1143) );
  CLKBUF_X3 U265 ( .A(SH[1]), .Z(n1144) );
  CLKBUF_X3 U266 ( .A(SH[1]), .Z(n1145) );
  CLKBUF_X3 U267 ( .A(SH[1]), .Z(n1146) );
  CLKBUF_X3 U268 ( .A(SH[1]), .Z(n1147) );
  CLKBUF_X3 U269 ( .A(SH[1]), .Z(n1148) );
  CLKBUF_X3 U270 ( .A(SH[1]), .Z(n1149) );
  CLKBUF_X3 U271 ( .A(SH[1]), .Z(n1150) );
  CLKBUF_X3 U272 ( .A(SH[1]), .Z(n1151) );
  INV_X1 U273 ( .A(n1157), .ZN(n1152) );
  INV_X1 U274 ( .A(n1157), .ZN(n1153) );
  INV_X1 U275 ( .A(n1156), .ZN(n1154) );
  INV_X1 U276 ( .A(n1157), .ZN(n1155) );
  INV_X1 U277 ( .A(SH[0]), .ZN(n1156) );
  INV_X1 U278 ( .A(SH[0]), .ZN(n1157) );
  NAND2_X2 U279 ( .A1(n1158), .A2(n1159), .ZN(B[9]) );
  MUX2_X1 U280 ( .A(n1160), .B(n1161), .S(n1152), .Z(n1159) );
  NAND2_X2 U281 ( .A1(n1150), .A2(n1162), .ZN(n1161) );
  NAND2_X2 U282 ( .A1(n1150), .A2(n1163), .ZN(n1160) );
  MUX2_X1 U283 ( .A(n1164), .B(n1165), .S(n1155), .Z(n1158) );
  NAND2_X2 U284 ( .A1(n1166), .A2(n1136), .ZN(n1165) );
  NAND2_X2 U285 ( .A1(n1167), .A2(n1134), .ZN(n1164) );
  NAND2_X2 U286 ( .A1(n1168), .A2(n1169), .ZN(B[8]) );
  MUX2_X1 U287 ( .A(n1170), .B(n1171), .S(n1155), .Z(n1169) );
  NAND2_X2 U288 ( .A1(n1150), .A2(n1163), .ZN(n1171) );
  NAND2_X2 U289 ( .A1(n1149), .A2(n1166), .ZN(n1170) );
  MUX2_X1 U290 ( .A(n1172), .B(n1173), .S(n1155), .Z(n1168) );
  NAND2_X2 U291 ( .A1(n1167), .A2(n1134), .ZN(n1173) );
  NAND2_X2 U292 ( .A1(n1174), .A2(n1134), .ZN(n1172) );
  NAND2_X2 U293 ( .A1(n1175), .A2(n1176), .ZN(B[7]) );
  MUX2_X1 U294 ( .A(n1177), .B(n1178), .S(n1155), .Z(n1176) );
  NAND2_X2 U295 ( .A1(n1149), .A2(n1166), .ZN(n1178) );
  NAND2_X2 U296 ( .A1(n1149), .A2(n1167), .ZN(n1177) );
  MUX2_X1 U297 ( .A(n1179), .B(n1180), .S(n1155), .Z(n1175) );
  NAND2_X2 U298 ( .A1(n1174), .A2(n1134), .ZN(n1180) );
  NAND2_X2 U299 ( .A1(n1181), .A2(n1134), .ZN(n1179) );
  NAND2_X2 U300 ( .A1(n1182), .A2(n1183), .ZN(B[6]) );
  MUX2_X1 U301 ( .A(n1184), .B(n1185), .S(n1155), .Z(n1183) );
  NAND2_X2 U302 ( .A1(n1149), .A2(n1167), .ZN(n1185) );
  NAND2_X2 U303 ( .A1(n1186), .A2(n1187), .ZN(n1167) );
  MUX2_X1 U304 ( .A(n1188), .B(n1189), .S(n1106), .Z(n1187) );
  NAND2_X2 U305 ( .A1(n1119), .A2(n1190), .ZN(n1189) );
  MUX2_X1 U306 ( .A(n1192), .B(n1193), .S(n1106), .Z(n1186) );
  NAND2_X2 U307 ( .A1(n1194), .A2(n1124), .ZN(n1193) );
  NAND2_X2 U308 ( .A1(n1195), .A2(n1123), .ZN(n1192) );
  NAND2_X2 U309 ( .A1(n1148), .A2(n1174), .ZN(n1184) );
  MUX2_X1 U310 ( .A(n1196), .B(n1197), .S(n1155), .Z(n1182) );
  NAND2_X2 U311 ( .A1(n1181), .A2(n1134), .ZN(n1197) );
  NAND2_X2 U312 ( .A1(n1198), .A2(n1134), .ZN(n1196) );
  NAND2_X2 U313 ( .A1(n1199), .A2(n1200), .ZN(B[5]) );
  MUX2_X1 U314 ( .A(n1201), .B(n1202), .S(n1155), .Z(n1200) );
  NAND2_X2 U315 ( .A1(n1149), .A2(n1174), .ZN(n1202) );
  NAND2_X2 U316 ( .A1(n1203), .A2(n1204), .ZN(n1174) );
  MUX2_X1 U317 ( .A(n1205), .B(n1206), .S(n1106), .Z(n1204) );
  NAND2_X2 U318 ( .A1(n1122), .A2(n1207), .ZN(n1206) );
  NAND2_X2 U319 ( .A1(n1122), .A2(n1208), .ZN(n1205) );
  MUX2_X1 U320 ( .A(n1209), .B(n1210), .S(n1106), .Z(n1203) );
  NAND2_X2 U321 ( .A1(n1211), .A2(n1123), .ZN(n1210) );
  NAND2_X2 U322 ( .A1(n1212), .A2(n1123), .ZN(n1209) );
  NAND2_X2 U323 ( .A1(n1148), .A2(n1181), .ZN(n1201) );
  MUX2_X1 U324 ( .A(n1213), .B(n1214), .S(n1155), .Z(n1199) );
  NAND2_X2 U325 ( .A1(n1198), .A2(n1134), .ZN(n1214) );
  NAND2_X2 U326 ( .A1(n1215), .A2(n1134), .ZN(n1213) );
  NAND2_X2 U327 ( .A1(n1216), .A2(n1217), .ZN(B[4]) );
  MUX2_X1 U328 ( .A(n1218), .B(n1219), .S(n1155), .Z(n1217) );
  NAND2_X2 U329 ( .A1(n1148), .A2(n1181), .ZN(n1219) );
  NAND2_X2 U330 ( .A1(n1220), .A2(n1221), .ZN(n1181) );
  MUX2_X1 U331 ( .A(n1222), .B(n1223), .S(n1106), .Z(n1221) );
  NAND2_X2 U332 ( .A1(n1122), .A2(n1225), .ZN(n1222) );
  MUX2_X1 U333 ( .A(n1226), .B(n1227), .S(n1106), .Z(n1220) );
  NAND2_X2 U334 ( .A1(n1228), .A2(n1123), .ZN(n1227) );
  NAND2_X2 U335 ( .A1(n1229), .A2(n1124), .ZN(n1226) );
  NAND2_X2 U336 ( .A1(n1148), .A2(n1198), .ZN(n1218) );
  MUX2_X1 U337 ( .A(n1230), .B(n1231), .S(n1154), .Z(n1216) );
  NAND2_X2 U338 ( .A1(n1215), .A2(n1134), .ZN(n1231) );
  NAND2_X2 U339 ( .A1(n1232), .A2(n1134), .ZN(n1230) );
  NAND2_X2 U340 ( .A1(n1233), .A2(n1234), .ZN(B[3]) );
  MUX2_X1 U341 ( .A(n1235), .B(n1236), .S(n1154), .Z(n1234) );
  NAND2_X2 U342 ( .A1(n1148), .A2(n1198), .ZN(n1236) );
  NAND2_X2 U343 ( .A1(n1237), .A2(n1238), .ZN(n1198) );
  MUX2_X1 U344 ( .A(n1239), .B(n1240), .S(n1106), .Z(n1238) );
  NAND2_X2 U345 ( .A1(n1122), .A2(n1241), .ZN(n1240) );
  MUX2_X1 U346 ( .A(n1243), .B(n1244), .S(n1106), .Z(n1237) );
  NAND2_X2 U347 ( .A1(n1245), .A2(n1128), .ZN(n1244) );
  NAND2_X2 U348 ( .A1(n1246), .A2(n1128), .ZN(n1243) );
  NAND2_X2 U349 ( .A1(n1147), .A2(n1215), .ZN(n1235) );
  MUX2_X1 U350 ( .A(n1247), .B(n1248), .S(n1154), .Z(n1233) );
  NAND2_X2 U351 ( .A1(n1232), .A2(n1134), .ZN(n1248) );
  NAND2_X2 U352 ( .A1(n1249), .A2(n1135), .ZN(n1247) );
  NAND2_X2 U353 ( .A1(n1250), .A2(n1251), .ZN(B[30]) );
  MUX2_X1 U354 ( .A(n1252), .B(n1253), .S(n1150), .Z(n1250) );
  NAND2_X2 U355 ( .A1(n1254), .A2(n1156), .ZN(n1252) );
  NAND2_X2 U356 ( .A1(n1255), .A2(n1256), .ZN(B[2]) );
  MUX2_X1 U357 ( .A(n1257), .B(n1258), .S(n1154), .Z(n1256) );
  NAND2_X2 U358 ( .A1(n1147), .A2(n1215), .ZN(n1258) );
  NAND2_X2 U359 ( .A1(n1259), .A2(n1260), .ZN(n1215) );
  MUX2_X1 U360 ( .A(n1261), .B(n1262), .S(n1106), .Z(n1260) );
  INV_X2 U361 ( .A(n1263), .ZN(n1195) );
  MUX2_X1 U362 ( .A(n1264), .B(n1265), .S(n1116), .Z(n1263) );
  MUX2_X1 U363 ( .A(n1266), .B(n1267), .S(n1106), .Z(n1259) );
  NAND2_X2 U364 ( .A1(n1268), .A2(n1129), .ZN(n1267) );
  NAND2_X2 U365 ( .A1(n1269), .A2(n1129), .ZN(n1266) );
  NAND2_X2 U366 ( .A1(n1147), .A2(n1232), .ZN(n1257) );
  MUX2_X1 U367 ( .A(n1270), .B(n1271), .S(n1154), .Z(n1255) );
  NAND2_X2 U368 ( .A1(n1249), .A2(n1135), .ZN(n1271) );
  NAND2_X2 U369 ( .A1(n1272), .A2(n1135), .ZN(n1270) );
  NAND2_X2 U370 ( .A1(n1273), .A2(n1274), .ZN(B[29]) );
  NAND3_X1 U371 ( .A1(n1156), .A2(n1138), .A3(n1275), .ZN(n1274) );
  MUX2_X1 U372 ( .A(n1276), .B(n1253), .S(n1150), .Z(n1273) );
  NAND2_X2 U373 ( .A1(n1152), .A2(n1254), .ZN(n1276) );
  NAND2_X2 U374 ( .A1(n1277), .A2(n1278), .ZN(B[28]) );
  MUX2_X1 U375 ( .A(n1279), .B(n1280), .S(n1154), .Z(n1278) );
  NAND2_X2 U376 ( .A1(n1147), .A2(n1254), .ZN(n1279) );
  MUX2_X1 U377 ( .A(n1281), .B(n1282), .S(n1154), .Z(n1277) );
  NAND2_X2 U378 ( .A1(n1275), .A2(n1135), .ZN(n1282) );
  NAND2_X2 U379 ( .A1(n1283), .A2(n1135), .ZN(n1281) );
  NAND2_X2 U380 ( .A1(n1284), .A2(n1285), .ZN(B[27]) );
  MUX2_X1 U381 ( .A(n1286), .B(n1287), .S(n1154), .Z(n1285) );
  NAND2_X2 U382 ( .A1(n1146), .A2(n1254), .ZN(n1287) );
  MUX2_X1 U383 ( .A(n1289), .B(n1253), .S(n1122), .Z(n1288) );
  NAND2_X2 U384 ( .A1(n1290), .A2(n1110), .ZN(n1289) );
  NAND2_X2 U385 ( .A1(n1146), .A2(n1275), .ZN(n1286) );
  MUX2_X1 U386 ( .A(n1291), .B(n1292), .S(n1154), .Z(n1284) );
  NAND2_X2 U387 ( .A1(n1283), .A2(n1135), .ZN(n1292) );
  NAND2_X2 U388 ( .A1(n1293), .A2(n1135), .ZN(n1291) );
  NAND2_X2 U389 ( .A1(n1294), .A2(n1295), .ZN(B[26]) );
  MUX2_X1 U390 ( .A(n1296), .B(n1297), .S(n1154), .Z(n1295) );
  NAND2_X2 U391 ( .A1(n1146), .A2(n1275), .ZN(n1297) );
  MUX2_X1 U392 ( .A(n1299), .B(n1253), .S(n1122), .Z(n1298) );
  NAND2_X2 U393 ( .A1(n1190), .A2(n1110), .ZN(n1299) );
  NAND2_X2 U394 ( .A1(n1146), .A2(n1283), .ZN(n1296) );
  MUX2_X1 U395 ( .A(n1300), .B(n1301), .S(n1154), .Z(n1294) );
  NAND2_X2 U396 ( .A1(n1293), .A2(n1135), .ZN(n1301) );
  NAND2_X2 U397 ( .A1(n1302), .A2(n1135), .ZN(n1300) );
  NAND2_X2 U398 ( .A1(n1303), .A2(n1304), .ZN(B[25]) );
  MUX2_X1 U399 ( .A(n1305), .B(n1306), .S(n1154), .Z(n1304) );
  NAND2_X2 U400 ( .A1(n1146), .A2(n1283), .ZN(n1306) );
  MUX2_X1 U401 ( .A(n1308), .B(n1253), .S(n1122), .Z(n1307) );
  NAND2_X2 U402 ( .A1(n1207), .A2(n1110), .ZN(n1308) );
  NAND2_X2 U403 ( .A1(n1145), .A2(n1293), .ZN(n1305) );
  MUX2_X1 U404 ( .A(n1309), .B(n1310), .S(n1154), .Z(n1303) );
  NAND2_X2 U405 ( .A1(n1302), .A2(n1135), .ZN(n1310) );
  NAND2_X2 U406 ( .A1(n1311), .A2(n1135), .ZN(n1309) );
  NAND2_X2 U407 ( .A1(n1312), .A2(n1313), .ZN(B[24]) );
  MUX2_X1 U408 ( .A(n1314), .B(n1315), .S(n1154), .Z(n1313) );
  NAND2_X2 U409 ( .A1(n1145), .A2(n1293), .ZN(n1315) );
  MUX2_X1 U410 ( .A(n1317), .B(n1253), .S(n1122), .Z(n1316) );
  NAND2_X2 U411 ( .A1(n1224), .A2(n1110), .ZN(n1317) );
  NAND2_X2 U412 ( .A1(n1145), .A2(n1302), .ZN(n1314) );
  MUX2_X1 U413 ( .A(n1318), .B(n1319), .S(n1154), .Z(n1312) );
  NAND2_X2 U414 ( .A1(n1311), .A2(n1135), .ZN(n1319) );
  NAND2_X2 U415 ( .A1(n1320), .A2(n1136), .ZN(n1318) );
  NAND2_X2 U416 ( .A1(n1321), .A2(n1322), .ZN(B[23]) );
  MUX2_X1 U417 ( .A(n1323), .B(n1324), .S(n1154), .Z(n1322) );
  NAND2_X2 U418 ( .A1(n1145), .A2(n1302), .ZN(n1324) );
  NAND2_X2 U419 ( .A1(n1325), .A2(n1326), .ZN(n1302) );
  NAND3_X1 U420 ( .A1(n1131), .A2(n1113), .A3(n1241), .ZN(n1326) );
  MUX2_X1 U421 ( .A(n1327), .B(n1253), .S(n1106), .Z(n1325) );
  NAND2_X2 U422 ( .A1(n1121), .A2(n1290), .ZN(n1327) );
  NAND2_X2 U423 ( .A1(n1144), .A2(n1311), .ZN(n1323) );
  MUX2_X1 U424 ( .A(n1328), .B(n1329), .S(n1154), .Z(n1321) );
  NAND2_X2 U425 ( .A1(n1320), .A2(n1136), .ZN(n1329) );
  NAND2_X2 U426 ( .A1(n1330), .A2(n1136), .ZN(n1328) );
  NAND2_X2 U427 ( .A1(n1331), .A2(n1332), .ZN(B[22]) );
  MUX2_X1 U428 ( .A(n1333), .B(n1334), .S(n1153), .Z(n1332) );
  NAND2_X2 U429 ( .A1(n1144), .A2(n1311), .ZN(n1334) );
  NAND2_X2 U430 ( .A1(n1335), .A2(n1336), .ZN(n1311) );
  NAND3_X1 U431 ( .A1(n1131), .A2(n1113), .A3(n1194), .ZN(n1336) );
  MUX2_X1 U432 ( .A(n1337), .B(n1253), .S(n1106), .Z(n1335) );
  NAND2_X2 U433 ( .A1(n1121), .A2(n1190), .ZN(n1337) );
  NAND2_X2 U434 ( .A1(n1144), .A2(n1320), .ZN(n1333) );
  MUX2_X1 U435 ( .A(n1338), .B(n1339), .S(n1153), .Z(n1331) );
  NAND2_X2 U436 ( .A1(n1330), .A2(n1136), .ZN(n1339) );
  NAND2_X2 U437 ( .A1(n1340), .A2(n1136), .ZN(n1338) );
  NAND2_X2 U438 ( .A1(n1341), .A2(n1342), .ZN(B[21]) );
  MUX2_X1 U439 ( .A(n1343), .B(n1344), .S(n1153), .Z(n1342) );
  NAND2_X2 U440 ( .A1(n1144), .A2(n1320), .ZN(n1344) );
  NAND2_X2 U441 ( .A1(n1345), .A2(n1346), .ZN(n1320) );
  NAND3_X1 U442 ( .A1(n1131), .A2(n1112), .A3(n1211), .ZN(n1346) );
  MUX2_X1 U443 ( .A(n1347), .B(n1253), .S(n1107), .Z(n1345) );
  NAND2_X2 U444 ( .A1(n1144), .A2(n1330), .ZN(n1343) );
  MUX2_X1 U445 ( .A(n1348), .B(n1349), .S(n1153), .Z(n1341) );
  NAND2_X2 U446 ( .A1(n1340), .A2(n1136), .ZN(n1349) );
  NAND2_X2 U447 ( .A1(n1350), .A2(n1136), .ZN(n1348) );
  NAND2_X2 U448 ( .A1(n1351), .A2(n1352), .ZN(B[20]) );
  MUX2_X1 U449 ( .A(n1353), .B(n1354), .S(n1153), .Z(n1352) );
  NAND2_X2 U450 ( .A1(n1143), .A2(n1330), .ZN(n1354) );
  NAND2_X2 U451 ( .A1(n1355), .A2(n1356), .ZN(n1330) );
  NAND3_X1 U452 ( .A1(n1131), .A2(n1112), .A3(n1228), .ZN(n1356) );
  MUX2_X1 U453 ( .A(n1357), .B(n1253), .S(n1107), .Z(n1355) );
  NAND2_X2 U454 ( .A1(n1121), .A2(n1224), .ZN(n1357) );
  NAND2_X2 U455 ( .A1(n1143), .A2(n1340), .ZN(n1353) );
  MUX2_X1 U456 ( .A(n1358), .B(n1359), .S(n1153), .Z(n1351) );
  NAND2_X2 U457 ( .A1(n1350), .A2(n1136), .ZN(n1359) );
  NAND2_X2 U458 ( .A1(n1360), .A2(n1136), .ZN(n1358) );
  NAND2_X2 U459 ( .A1(n1361), .A2(n1362), .ZN(B[1]) );
  MUX2_X1 U460 ( .A(n1363), .B(n1364), .S(n1153), .Z(n1362) );
  NAND2_X2 U461 ( .A1(n1143), .A2(n1232), .ZN(n1364) );
  NAND2_X2 U462 ( .A1(n1365), .A2(n1366), .ZN(n1232) );
  MUX2_X1 U463 ( .A(n1367), .B(n1368), .S(n1107), .Z(n1366) );
  NAND2_X2 U464 ( .A1(n1121), .A2(n1211), .ZN(n1368) );
  NAND2_X2 U465 ( .A1(n1121), .A2(n1212), .ZN(n1367) );
  INV_X2 U466 ( .A(n1369), .ZN(n1212) );
  MUX2_X1 U467 ( .A(n1370), .B(n1371), .S(n1116), .Z(n1369) );
  MUX2_X1 U468 ( .A(n1372), .B(n1373), .S(n1107), .Z(n1365) );
  NAND2_X2 U469 ( .A1(n1374), .A2(n1129), .ZN(n1373) );
  NAND2_X2 U470 ( .A1(n1375), .A2(n1129), .ZN(n1372) );
  NAND2_X2 U471 ( .A1(n1143), .A2(n1249), .ZN(n1363) );
  MUX2_X1 U472 ( .A(n1376), .B(n1377), .S(n1153), .Z(n1361) );
  NAND2_X2 U473 ( .A1(n1272), .A2(n1136), .ZN(n1377) );
  NAND2_X2 U474 ( .A1(n1378), .A2(n1136), .ZN(n1376) );
  NAND2_X2 U475 ( .A1(n1379), .A2(n1380), .ZN(B[19]) );
  MUX2_X1 U476 ( .A(n1381), .B(n1382), .S(n1153), .Z(n1380) );
  NAND2_X2 U477 ( .A1(n1143), .A2(n1340), .ZN(n1382) );
  NAND2_X2 U478 ( .A1(n1383), .A2(n1384), .ZN(n1340) );
  NAND3_X1 U479 ( .A1(n1130), .A2(n1113), .A3(n1245), .ZN(n1384) );
  MUX2_X1 U480 ( .A(n1385), .B(n1253), .S(n1107), .Z(n1383) );
  NAND2_X2 U481 ( .A1(n1121), .A2(n1241), .ZN(n1385) );
  NAND2_X2 U482 ( .A1(n1142), .A2(n1350), .ZN(n1381) );
  MUX2_X1 U483 ( .A(n1386), .B(n1387), .S(n1153), .Z(n1379) );
  NAND2_X2 U484 ( .A1(n1360), .A2(n1137), .ZN(n1387) );
  NAND2_X2 U485 ( .A1(n1388), .A2(n1137), .ZN(n1386) );
  NAND2_X2 U486 ( .A1(n1389), .A2(n1390), .ZN(B[18]) );
  MUX2_X1 U487 ( .A(n1391), .B(n1392), .S(n1153), .Z(n1390) );
  NAND2_X2 U488 ( .A1(n1142), .A2(n1350), .ZN(n1392) );
  NAND2_X2 U489 ( .A1(n1393), .A2(n1394), .ZN(n1350) );
  NAND3_X1 U490 ( .A1(n1131), .A2(n1112), .A3(n1268), .ZN(n1394) );
  MUX2_X1 U491 ( .A(n1395), .B(n1253), .S(n1107), .Z(n1393) );
  INV_X2 U492 ( .A(n1396), .ZN(n1194) );
  MUX2_X1 U493 ( .A(n1397), .B(n1253), .S(n1116), .Z(n1396) );
  NAND2_X2 U494 ( .A1(n1142), .A2(n1360), .ZN(n1391) );
  MUX2_X1 U495 ( .A(n1398), .B(n1399), .S(n1153), .Z(n1389) );
  NAND2_X2 U496 ( .A1(n1388), .A2(n1137), .ZN(n1399) );
  NAND2_X2 U497 ( .A1(n1400), .A2(n1137), .ZN(n1398) );
  NAND2_X2 U498 ( .A1(n1401), .A2(n1402), .ZN(B[17]) );
  MUX2_X1 U499 ( .A(n1403), .B(n1404), .S(n1153), .Z(n1402) );
  NAND2_X2 U500 ( .A1(n1142), .A2(n1360), .ZN(n1404) );
  NAND2_X2 U501 ( .A1(n1405), .A2(n1406), .ZN(n1360) );
  NAND3_X1 U502 ( .A1(n1131), .A2(n1113), .A3(n1374), .ZN(n1406) );
  MUX2_X1 U503 ( .A(n1407), .B(n1253), .S(n1107), .Z(n1405) );
  INV_X2 U504 ( .A(n1408), .ZN(n1211) );
  MUX2_X1 U505 ( .A(n1409), .B(n1253), .S(n1116), .Z(n1408) );
  NAND2_X2 U506 ( .A1(n1142), .A2(n1388), .ZN(n1403) );
  MUX2_X1 U507 ( .A(n1410), .B(n1411), .S(n1153), .Z(n1401) );
  NAND2_X2 U508 ( .A1(n1400), .A2(n1137), .ZN(n1411) );
  NAND2_X2 U509 ( .A1(n1412), .A2(n1137), .ZN(n1410) );
  NAND2_X2 U510 ( .A1(n1413), .A2(n1414), .ZN(B[16]) );
  MUX2_X1 U511 ( .A(n1415), .B(n1416), .S(n1153), .Z(n1414) );
  NAND2_X2 U512 ( .A1(n1141), .A2(n1388), .ZN(n1416) );
  NAND2_X2 U513 ( .A1(n1417), .A2(n1418), .ZN(n1388) );
  NAND3_X1 U514 ( .A1(n1132), .A2(n1114), .A3(n1419), .ZN(n1418) );
  MUX2_X1 U515 ( .A(n1420), .B(n1253), .S(n1107), .Z(n1417) );
  NAND2_X2 U516 ( .A1(n1141), .A2(n1400), .ZN(n1415) );
  MUX2_X1 U517 ( .A(n1421), .B(n1422), .S(n1152), .Z(n1413) );
  NAND2_X2 U518 ( .A1(n1412), .A2(n1137), .ZN(n1422) );
  NAND2_X2 U519 ( .A1(n1423), .A2(n1137), .ZN(n1421) );
  NAND2_X2 U520 ( .A1(n1424), .A2(n1425), .ZN(B[15]) );
  MUX2_X1 U521 ( .A(n1426), .B(n1427), .S(n1152), .Z(n1425) );
  NAND2_X2 U522 ( .A1(n1141), .A2(n1400), .ZN(n1427) );
  NAND2_X2 U523 ( .A1(n1428), .A2(n1429), .ZN(n1400) );
  NAND3_X1 U524 ( .A1(n1131), .A2(n1113), .A3(n1430), .ZN(n1429) );
  MUX2_X1 U525 ( .A(n1431), .B(n1253), .S(n1107), .Z(n1428) );
  NAND2_X2 U526 ( .A1(n1141), .A2(n1412), .ZN(n1426) );
  MUX2_X1 U527 ( .A(n1432), .B(n1433), .S(n1152), .Z(n1424) );
  NAND2_X2 U528 ( .A1(n1423), .A2(n1137), .ZN(n1433) );
  NAND2_X2 U529 ( .A1(n1434), .A2(n1137), .ZN(n1432) );
  NAND2_X2 U530 ( .A1(n1435), .A2(n1436), .ZN(B[14]) );
  MUX2_X1 U531 ( .A(n1437), .B(n1438), .S(n1152), .Z(n1436) );
  NAND2_X2 U532 ( .A1(n1141), .A2(n1412), .ZN(n1438) );
  NAND2_X2 U533 ( .A1(n1439), .A2(n1440), .ZN(n1412) );
  NAND3_X1 U534 ( .A1(n1132), .A2(n1113), .A3(n1441), .ZN(n1440) );
  MUX2_X1 U535 ( .A(n1442), .B(n1253), .S(n1107), .Z(n1439) );
  NAND2_X2 U536 ( .A1(n1140), .A2(n1423), .ZN(n1437) );
  MUX2_X1 U537 ( .A(n1443), .B(n1444), .S(n1152), .Z(n1435) );
  NAND2_X2 U538 ( .A1(n1434), .A2(n1137), .ZN(n1444) );
  NAND2_X2 U539 ( .A1(n1446), .A2(n1447), .ZN(B[13]) );
  MUX2_X1 U540 ( .A(n1448), .B(n1449), .S(n1152), .Z(n1447) );
  NAND2_X2 U541 ( .A1(n1140), .A2(n1423), .ZN(n1449) );
  NAND2_X2 U542 ( .A1(n1450), .A2(n1451), .ZN(n1423) );
  NAND3_X1 U543 ( .A1(n1132), .A2(n1113), .A3(n1452), .ZN(n1451) );
  MUX2_X1 U544 ( .A(n1453), .B(n1253), .S(n1107), .Z(n1450) );
  NAND2_X2 U545 ( .A1(n1140), .A2(n1434), .ZN(n1448) );
  MUX2_X1 U546 ( .A(n1454), .B(n1455), .S(n1152), .Z(n1446) );
  NAND2_X2 U547 ( .A1(n1456), .A2(n1138), .ZN(n1454) );
  NAND2_X2 U548 ( .A1(n1457), .A2(n1458), .ZN(B[12]) );
  MUX2_X1 U549 ( .A(n1459), .B(n1460), .S(n1152), .Z(n1458) );
  NAND2_X2 U550 ( .A1(n1140), .A2(n1434), .ZN(n1460) );
  NAND2_X2 U551 ( .A1(n1461), .A2(n1462), .ZN(n1434) );
  NAND3_X1 U552 ( .A1(n1132), .A2(n1114), .A3(n1463), .ZN(n1462) );
  MUX2_X1 U553 ( .A(n1464), .B(n1253), .S(n1107), .Z(n1461) );
  MUX2_X1 U554 ( .A(n1465), .B(n1466), .S(n1152), .Z(n1457) );
  NAND2_X2 U555 ( .A1(n1456), .A2(n1138), .ZN(n1466) );
  NAND2_X2 U556 ( .A1(n1162), .A2(n1138), .ZN(n1465) );
  NAND2_X2 U557 ( .A1(n1467), .A2(n1468), .ZN(B[11]) );
  MUX2_X1 U558 ( .A(n1469), .B(n1470), .S(n1152), .Z(n1468) );
  NAND2_X2 U559 ( .A1(n1471), .A2(n1472), .ZN(n1445) );
  MUX2_X1 U560 ( .A(n1473), .B(n1474), .S(n1108), .Z(n1472) );
  MUX2_X1 U561 ( .A(n1475), .B(n1476), .S(n1108), .Z(n1471) );
  NAND2_X2 U562 ( .A1(n1290), .A2(n1128), .ZN(n1476) );
  NAND2_X2 U563 ( .A1(n1477), .A2(n1128), .ZN(n1475) );
  NAND2_X2 U564 ( .A1(n1139), .A2(n1456), .ZN(n1469) );
  MUX2_X1 U565 ( .A(n1478), .B(n1479), .S(n1153), .Z(n1467) );
  NAND2_X2 U566 ( .A1(n1162), .A2(n1138), .ZN(n1479) );
  NAND2_X2 U567 ( .A1(n1163), .A2(n1138), .ZN(n1478) );
  NAND2_X2 U568 ( .A1(n1480), .A2(n1481), .ZN(B[10]) );
  MUX2_X1 U569 ( .A(n1482), .B(n1483), .S(n1152), .Z(n1481) );
  NAND2_X2 U570 ( .A1(n1139), .A2(n1456), .ZN(n1483) );
  NAND2_X2 U571 ( .A1(n1484), .A2(n1485), .ZN(n1456) );
  MUX2_X1 U572 ( .A(n1486), .B(n1487), .S(n1108), .Z(n1485) );
  MUX2_X1 U573 ( .A(n1488), .B(n1489), .S(n1108), .Z(n1484) );
  NAND2_X2 U574 ( .A1(n1190), .A2(n1127), .ZN(n1489) );
  INV_X2 U575 ( .A(n1490), .ZN(n1190) );
  MUX2_X1 U576 ( .A(n1491), .B(n1253), .S(n1116), .Z(n1490) );
  NAND2_X2 U577 ( .A1(n1191), .A2(n1127), .ZN(n1488) );
  INV_X2 U578 ( .A(n1492), .ZN(n1191) );
  MUX2_X1 U579 ( .A(n1493), .B(n1494), .S(n1116), .Z(n1492) );
  NAND2_X2 U580 ( .A1(n1139), .A2(n1162), .ZN(n1482) );
  NAND2_X2 U581 ( .A1(n1495), .A2(n1496), .ZN(n1162) );
  MUX2_X1 U582 ( .A(n1497), .B(n1498), .S(n1108), .Z(n1496) );
  NAND2_X2 U583 ( .A1(n1119), .A2(n1452), .ZN(n1497) );
  MUX2_X1 U584 ( .A(n1499), .B(n1500), .S(n1108), .Z(n1495) );
  NAND2_X2 U585 ( .A1(n1207), .A2(n1127), .ZN(n1500) );
  INV_X2 U586 ( .A(n1501), .ZN(n1207) );
  MUX2_X1 U587 ( .A(n1502), .B(n1253), .S(n1116), .Z(n1501) );
  NAND2_X2 U588 ( .A1(n1208), .A2(n1127), .ZN(n1499) );
  INV_X2 U589 ( .A(n1503), .ZN(n1208) );
  MUX2_X1 U590 ( .A(n1504), .B(n1505), .S(n1116), .Z(n1503) );
  MUX2_X1 U591 ( .A(n1506), .B(n1507), .S(n1152), .Z(n1480) );
  NAND2_X2 U592 ( .A1(n1163), .A2(n1138), .ZN(n1507) );
  NAND2_X2 U593 ( .A1(n1508), .A2(n1509), .ZN(n1163) );
  MUX2_X1 U594 ( .A(n1510), .B(n1511), .S(n1108), .Z(n1509) );
  INV_X2 U595 ( .A(n1512), .ZN(n1463) );
  MUX2_X1 U596 ( .A(n1513), .B(n1514), .S(n1116), .Z(n1512) );
  MUX2_X1 U597 ( .A(n1515), .B(n1516), .S(n1108), .Z(n1508) );
  NAND2_X2 U598 ( .A1(n1224), .A2(n1126), .ZN(n1516) );
  INV_X2 U599 ( .A(n1517), .ZN(n1224) );
  MUX2_X1 U600 ( .A(n1518), .B(n1253), .S(n1116), .Z(n1517) );
  NAND2_X2 U601 ( .A1(n1225), .A2(n1126), .ZN(n1515) );
  INV_X2 U602 ( .A(n1519), .ZN(n1225) );
  MUX2_X1 U603 ( .A(n1520), .B(n1521), .S(n1116), .Z(n1519) );
  NAND2_X2 U604 ( .A1(n1166), .A2(n1138), .ZN(n1506) );
  NAND2_X2 U605 ( .A1(n1522), .A2(n1523), .ZN(n1166) );
  MUX2_X1 U606 ( .A(n1524), .B(n1525), .S(n1108), .Z(n1523) );
  NAND2_X2 U607 ( .A1(n1119), .A2(n1290), .ZN(n1525) );
  INV_X2 U608 ( .A(n1526), .ZN(n1290) );
  MUX2_X1 U609 ( .A(n1527), .B(n1253), .S(n1116), .Z(n1526) );
  NAND2_X2 U610 ( .A1(n1119), .A2(n1477), .ZN(n1524) );
  INV_X2 U611 ( .A(n1528), .ZN(n1477) );
  MUX2_X1 U612 ( .A(n1529), .B(n1530), .S(n1117), .Z(n1528) );
  MUX2_X1 U613 ( .A(n1531), .B(n1532), .S(n1108), .Z(n1522) );
  NAND2_X2 U614 ( .A1(n1241), .A2(n1126), .ZN(n1532) );
  INV_X2 U615 ( .A(n1533), .ZN(n1241) );
  MUX2_X1 U616 ( .A(n1534), .B(n1253), .S(n1117), .Z(n1533) );
  NAND2_X2 U617 ( .A1(n1242), .A2(n1126), .ZN(n1531) );
  INV_X2 U618 ( .A(n1535), .ZN(n1242) );
  MUX2_X1 U619 ( .A(n1536), .B(n1537), .S(n1117), .Z(n1535) );
  NAND2_X2 U620 ( .A1(n1538), .A2(n1539), .ZN(B[0]) );
  MUX2_X1 U621 ( .A(n1540), .B(n1541), .S(n1152), .Z(n1539) );
  NAND2_X2 U622 ( .A1(n1139), .A2(n1249), .ZN(n1541) );
  NAND2_X2 U623 ( .A1(n1542), .A2(n1543), .ZN(n1249) );
  MUX2_X1 U624 ( .A(n1544), .B(n1545), .S(n1108), .Z(n1543) );
  NAND2_X2 U625 ( .A1(n1119), .A2(n1228), .ZN(n1545) );
  INV_X2 U626 ( .A(n1546), .ZN(n1228) );
  MUX2_X1 U627 ( .A(n1514), .B(n1253), .S(n1117), .Z(n1546) );
  INV_X2 U628 ( .A(A[23]), .ZN(n1514) );
  NAND2_X2 U629 ( .A1(n1119), .A2(n1229), .ZN(n1544) );
  INV_X2 U630 ( .A(n1547), .ZN(n1229) );
  MUX2_X1 U631 ( .A(n1548), .B(n1513), .S(n1117), .Z(n1547) );
  MUX2_X1 U632 ( .A(n1549), .B(n1550), .S(n1108), .Z(n1542) );
  NAND2_X2 U633 ( .A1(n1419), .A2(n1125), .ZN(n1550) );
  INV_X2 U634 ( .A(n1551), .ZN(n1419) );
  MUX2_X1 U635 ( .A(n1521), .B(n1518), .S(n1117), .Z(n1551) );
  NAND2_X2 U636 ( .A1(n1552), .A2(n1125), .ZN(n1549) );
  MUX2_X1 U637 ( .A(A[3]), .B(A[11]), .S(n1117), .Z(n1552) );
  NAND2_X2 U638 ( .A1(n1145), .A2(n1272), .ZN(n1540) );
  NAND2_X2 U639 ( .A1(n1553), .A2(n1554), .ZN(n1272) );
  MUX2_X1 U640 ( .A(n1555), .B(n1556), .S(n1109), .Z(n1554) );
  NAND2_X2 U641 ( .A1(n1119), .A2(n1245), .ZN(n1556) );
  INV_X2 U642 ( .A(n1557), .ZN(n1245) );
  MUX2_X1 U643 ( .A(n1530), .B(n1527), .S(n1117), .Z(n1557) );
  NAND2_X2 U644 ( .A1(n1119), .A2(n1246), .ZN(n1555) );
  INV_X2 U645 ( .A(n1558), .ZN(n1246) );
  MUX2_X1 U646 ( .A(n1559), .B(n1529), .S(n1117), .Z(n1558) );
  MUX2_X1 U647 ( .A(n1560), .B(n1561), .S(n1109), .Z(n1553) );
  NAND2_X2 U648 ( .A1(n1430), .A2(n1125), .ZN(n1561) );
  INV_X2 U649 ( .A(n1562), .ZN(n1430) );
  MUX2_X1 U650 ( .A(n1537), .B(n1534), .S(n1117), .Z(n1562) );
  NAND2_X2 U651 ( .A1(n1563), .A2(n1125), .ZN(n1560) );
  MUX2_X1 U652 ( .A(A[2]), .B(A[10]), .S(n1117), .Z(n1563) );
  MUX2_X1 U653 ( .A(n1564), .B(n1565), .S(n1153), .Z(n1538) );
  NAND2_X2 U654 ( .A1(n1378), .A2(n1138), .ZN(n1565) );
  NAND2_X2 U655 ( .A1(n1566), .A2(n1567), .ZN(n1378) );
  MUX2_X1 U656 ( .A(n1568), .B(n1569), .S(n1109), .Z(n1567) );
  NAND2_X2 U657 ( .A1(n1119), .A2(n1268), .ZN(n1569) );
  INV_X2 U658 ( .A(n1570), .ZN(n1268) );
  MUX2_X1 U659 ( .A(n1494), .B(n1491), .S(n1117), .Z(n1570) );
  NAND2_X2 U660 ( .A1(n1119), .A2(n1269), .ZN(n1568) );
  INV_X2 U661 ( .A(n1571), .ZN(n1269) );
  MUX2_X1 U662 ( .A(n1572), .B(n1493), .S(n1118), .Z(n1571) );
  MUX2_X1 U663 ( .A(n1573), .B(n1574), .S(n1109), .Z(n1566) );
  NAND2_X2 U664 ( .A1(n1441), .A2(n1124), .ZN(n1574) );
  INV_X2 U665 ( .A(n1575), .ZN(n1441) );
  MUX2_X1 U666 ( .A(n1265), .B(n1397), .S(n1118), .Z(n1575) );
  NAND2_X2 U667 ( .A1(n1576), .A2(n1124), .ZN(n1573) );
  MUX2_X1 U668 ( .A(A[1]), .B(A[9]), .S(n1118), .Z(n1576) );
  OAI21_X2 U669 ( .B1(n1577), .B2(n1578), .A(n1138), .ZN(n1564) );
  MUX2_X1 U670 ( .A(n1579), .B(n1580), .S(n1109), .Z(n1578) );
  AND2_X2 U671 ( .A1(n1452), .A2(n1130), .ZN(n1580) );
  INV_X2 U672 ( .A(n1581), .ZN(n1452) );
  MUX2_X1 U673 ( .A(n1371), .B(n1409), .S(n1118), .Z(n1581) );
  AND2_X2 U674 ( .A1(n1582), .A2(n1130), .ZN(n1579) );
  MUX2_X1 U675 ( .A(A[0]), .B(A[8]), .S(n1118), .Z(n1582) );
  MUX2_X1 U676 ( .A(n1583), .B(n1584), .S(n1109), .Z(n1577) );
  AND2_X2 U677 ( .A1(n1122), .A2(n1374), .ZN(n1584) );
  INV_X2 U678 ( .A(n1585), .ZN(n1374) );
  MUX2_X1 U679 ( .A(n1505), .B(n1502), .S(n1118), .Z(n1585) );
  AND2_X2 U680 ( .A1(n1122), .A2(n1375), .ZN(n1583) );
  INV_X2 U681 ( .A(n1586), .ZN(n1375) );
  MUX2_X1 U682 ( .A(n1587), .B(n1504), .S(n1118), .Z(n1586) );
endmodule


module Xi_core_DW_rightsh_1 ( A, SH, B, DATA_TC );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633;

  NAND2_X1 U108 ( .A1(A[24]), .A2(n1178), .ZN(n1420) );
  INV_X1 U109 ( .A(A[24]), .ZN(n1604) );
  INV_X1 U110 ( .A(A[28]), .ZN(n1590) );
  NAND2_X1 U111 ( .A1(A[28]), .A2(n1181), .ZN(n1539) );
  INV_X1 U112 ( .A(A[4]), .ZN(n1620) );
  NAND2_X1 U113 ( .A1(A[27]), .A2(n1180), .ZN(n1536) );
  NAND2_X1 U114 ( .A1(A[29]), .A2(n1180), .ZN(n1535) );
  INV_X1 U115 ( .A(A[1]), .ZN(n1633) );
  NAND2_X1 U116 ( .A1(A[25]), .A2(n1178), .ZN(n1410) );
  INV_X1 U117 ( .A(A[25]), .ZN(n1598) );
  INV_X1 U118 ( .A(A[2]), .ZN(n1626) );
  NAND2_X1 U119 ( .A1(A[30]), .A2(n1179), .ZN(n1530) );
  INV_X1 U120 ( .A(A[30]), .ZN(n1588) );
  INV_X1 U121 ( .A(A[22]), .ZN(n1554) );
  INV_X1 U122 ( .A(A[29]), .ZN(n1584) );
  INV_X1 U123 ( .A(A[27]), .ZN(n1596) );
  INV_X1 U124 ( .A(A[21]), .ZN(n1561) );
  INV_X1 U125 ( .A(A[31]), .ZN(n1582) );
  NAND2_X1 U126 ( .A1(A[31]), .A2(n1179), .ZN(n1528) );
  INV_X1 U127 ( .A(A[6]), .ZN(n1618) );
  INV_X1 U128 ( .A(A[7]), .ZN(n1612) );
  INV_X1 U129 ( .A(A[5]), .ZN(n1614) );
  INV_X1 U130 ( .A(A[19]), .ZN(n1564) );
  INV_X1 U131 ( .A(A[18]), .ZN(n1572) );
  INV_X1 U132 ( .A(A[16]), .ZN(n1385) );
  INV_X1 U133 ( .A(A[13]), .ZN(n1560) );
  INV_X1 U134 ( .A(A[17]), .ZN(n1324) );
  INV_X1 U135 ( .A(A[15]), .ZN(n1548) );
  INV_X1 U136 ( .A(A[14]), .ZN(n1553) );
  INV_X1 U137 ( .A(A[20]), .ZN(n1569) );
  INV_X1 U138 ( .A(A[12]), .ZN(n1568) );
  INV_X1 U139 ( .A(A[9]), .ZN(n1323) );
  INV_X1 U140 ( .A(A[11]), .ZN(n1563) );
  INV_X1 U141 ( .A(A[8]), .ZN(n1384) );
  INV_X1 U142 ( .A(A[10]), .ZN(n1571) );
  INV_X1 U143 ( .A(n1168), .ZN(n1163) );
  INV_X1 U144 ( .A(n1173), .ZN(n1164) );
  INV_X1 U145 ( .A(n1174), .ZN(n1165) );
  INV_X1 U146 ( .A(n1175), .ZN(n1166) );
  CLKBUF_X3 U147 ( .A(SH[4]), .Z(n1167) );
  CLKBUF_X3 U148 ( .A(SH[4]), .Z(n1168) );
  CLKBUF_X3 U149 ( .A(SH[4]), .Z(n1169) );
  CLKBUF_X3 U150 ( .A(SH[4]), .Z(n1170) );
  CLKBUF_X3 U151 ( .A(SH[4]), .Z(n1171) );
  CLKBUF_X3 U152 ( .A(SH[4]), .Z(n1172) );
  CLKBUF_X3 U153 ( .A(SH[4]), .Z(n1173) );
  CLKBUF_X3 U154 ( .A(SH[4]), .Z(n1174) );
  CLKBUF_X3 U155 ( .A(SH[4]), .Z(n1175) );
  INV_X1 U156 ( .A(n1182), .ZN(n1176) );
  INV_X1 U157 ( .A(n1182), .ZN(n1177) );
  INV_X1 U158 ( .A(SH[3]), .ZN(n1178) );
  INV_X1 U159 ( .A(SH[3]), .ZN(n1179) );
  INV_X1 U160 ( .A(SH[3]), .ZN(n1180) );
  INV_X1 U161 ( .A(SH[3]), .ZN(n1181) );
  INV_X1 U162 ( .A(SH[3]), .ZN(n1182) );
  INV_X1 U163 ( .A(n1186), .ZN(n1183) );
  INV_X1 U164 ( .A(n1186), .ZN(n1184) );
  INV_X1 U165 ( .A(n1186), .ZN(n1185) );
  INV_X8 U166 ( .A(SH[2]), .ZN(n1186) );
  INV_X1 U167 ( .A(n1192), .ZN(n1187) );
  INV_X1 U168 ( .A(n1192), .ZN(n1188) );
  INV_X1 U169 ( .A(n1192), .ZN(n1189) );
  INV_X1 U170 ( .A(n1192), .ZN(n1190) );
  INV_X2 U171 ( .A(SH[1]), .ZN(n1191) );
  INV_X2 U172 ( .A(SH[1]), .ZN(n1192) );
  INV_X1 U173 ( .A(n1206), .ZN(n1193) );
  INV_X1 U174 ( .A(n1204), .ZN(n1194) );
  INV_X1 U175 ( .A(n1207), .ZN(n1195) );
  INV_X1 U176 ( .A(n1205), .ZN(n1196) );
  INV_X1 U177 ( .A(n1203), .ZN(n1197) );
  CLKBUF_X3 U178 ( .A(SH[0]), .Z(n1198) );
  CLKBUF_X3 U179 ( .A(SH[0]), .Z(n1199) );
  CLKBUF_X3 U180 ( .A(SH[0]), .Z(n1200) );
  CLKBUF_X3 U181 ( .A(SH[0]), .Z(n1201) );
  CLKBUF_X3 U182 ( .A(SH[0]), .Z(n1202) );
  CLKBUF_X3 U183 ( .A(SH[0]), .Z(n1203) );
  CLKBUF_X3 U184 ( .A(SH[0]), .Z(n1204) );
  CLKBUF_X3 U185 ( .A(SH[0]), .Z(n1205) );
  CLKBUF_X3 U186 ( .A(SH[0]), .Z(n1206) );
  CLKBUF_X3 U187 ( .A(SH[0]), .Z(n1207) );
  CLKBUF_X3 U188 ( .A(SH[0]), .Z(n1208) );
  CLKBUF_X3 U189 ( .A(SH[0]), .Z(n1209) );
  CLKBUF_X3 U190 ( .A(SH[0]), .Z(n1210) );
  CLKBUF_X3 U191 ( .A(SH[0]), .Z(n1211) );
  NAND2_X2 U192 ( .A1(n1212), .A2(n1213), .ZN(B[9]) );
  MUX2_X1 U193 ( .A(n1214), .B(n1215), .S(n1183), .Z(n1213) );
  NAND2_X2 U194 ( .A1(n1174), .A2(n1216), .ZN(n1215) );
  NAND2_X2 U195 ( .A1(n1175), .A2(n1217), .ZN(n1214) );
  MUX2_X1 U196 ( .A(n1218), .B(n1219), .S(n1185), .Z(n1212) );
  NAND2_X2 U197 ( .A1(n1220), .A2(n1163), .ZN(n1219) );
  NAND2_X2 U198 ( .A1(n1221), .A2(n1163), .ZN(n1218) );
  NAND2_X2 U199 ( .A1(n1222), .A2(n1223), .ZN(B[8]) );
  MUX2_X1 U200 ( .A(n1224), .B(n1225), .S(n1185), .Z(n1223) );
  NAND2_X2 U201 ( .A1(n1174), .A2(n1226), .ZN(n1225) );
  NAND2_X2 U202 ( .A1(n1174), .A2(n1227), .ZN(n1224) );
  MUX2_X1 U203 ( .A(n1228), .B(n1229), .S(n1185), .Z(n1222) );
  NAND2_X2 U204 ( .A1(n1230), .A2(n1163), .ZN(n1229) );
  NAND2_X2 U205 ( .A1(n1231), .A2(n1163), .ZN(n1228) );
  NAND2_X2 U206 ( .A1(n1232), .A2(n1233), .ZN(B[7]) );
  MUX2_X1 U207 ( .A(n1234), .B(n1235), .S(n1185), .Z(n1233) );
  NAND2_X2 U208 ( .A1(n1174), .A2(n1236), .ZN(n1235) );
  NAND2_X2 U209 ( .A1(n1173), .A2(n1237), .ZN(n1234) );
  MUX2_X1 U210 ( .A(n1238), .B(n1239), .S(n1185), .Z(n1232) );
  NAND2_X2 U211 ( .A1(n1240), .A2(n1163), .ZN(n1239) );
  NAND2_X2 U212 ( .A1(n1241), .A2(n1163), .ZN(n1238) );
  NAND2_X2 U213 ( .A1(n1242), .A2(n1243), .ZN(B[6]) );
  MUX2_X1 U214 ( .A(n1244), .B(n1245), .S(n1185), .Z(n1243) );
  NAND2_X2 U215 ( .A1(n1173), .A2(n1246), .ZN(n1245) );
  NAND2_X2 U216 ( .A1(n1173), .A2(n1247), .ZN(n1244) );
  MUX2_X1 U217 ( .A(n1248), .B(n1249), .S(n1185), .Z(n1242) );
  NAND2_X2 U218 ( .A1(n1250), .A2(n1163), .ZN(n1249) );
  NAND2_X2 U219 ( .A1(n1251), .A2(n1164), .ZN(n1248) );
  NAND2_X2 U220 ( .A1(n1252), .A2(n1253), .ZN(B[5]) );
  MUX2_X1 U221 ( .A(n1254), .B(n1255), .S(n1185), .Z(n1253) );
  NAND2_X2 U222 ( .A1(n1173), .A2(n1217), .ZN(n1255) );
  NAND2_X2 U223 ( .A1(n1172), .A2(n1256), .ZN(n1254) );
  MUX2_X1 U224 ( .A(n1257), .B(n1258), .S(n1184), .Z(n1252) );
  NAND2_X2 U225 ( .A1(n1221), .A2(n1164), .ZN(n1258) );
  NAND2_X2 U226 ( .A1(n1259), .A2(n1260), .ZN(n1221) );
  MUX2_X1 U227 ( .A(n1261), .B(n1262), .S(n1187), .Z(n1260) );
  NAND2_X2 U228 ( .A1(n1209), .A2(n1263), .ZN(n1262) );
  NAND2_X2 U229 ( .A1(n1210), .A2(n1264), .ZN(n1261) );
  MUX2_X1 U230 ( .A(n1265), .B(n1266), .S(n1190), .Z(n1259) );
  NAND2_X2 U231 ( .A1(n1267), .A2(n1195), .ZN(n1266) );
  NAND2_X2 U232 ( .A1(n1268), .A2(n1193), .ZN(n1265) );
  NAND2_X2 U233 ( .A1(n1269), .A2(n1164), .ZN(n1257) );
  NAND2_X2 U234 ( .A1(n1270), .A2(n1271), .ZN(B[4]) );
  MUX2_X1 U235 ( .A(n1272), .B(n1273), .S(n1184), .Z(n1271) );
  NAND2_X2 U236 ( .A1(n1172), .A2(n1227), .ZN(n1273) );
  NAND2_X2 U237 ( .A1(n1172), .A2(n1274), .ZN(n1272) );
  MUX2_X1 U238 ( .A(n1275), .B(n1276), .S(n1184), .Z(n1270) );
  NAND2_X2 U239 ( .A1(n1231), .A2(n1164), .ZN(n1276) );
  NAND2_X2 U240 ( .A1(n1277), .A2(n1278), .ZN(n1231) );
  MUX2_X1 U241 ( .A(n1279), .B(n1280), .S(n1190), .Z(n1278) );
  NAND2_X2 U242 ( .A1(n1209), .A2(n1267), .ZN(n1280) );
  NAND2_X2 U243 ( .A1(n1210), .A2(n1268), .ZN(n1279) );
  MUX2_X1 U244 ( .A(n1281), .B(n1282), .S(n1190), .Z(n1277) );
  NAND2_X2 U245 ( .A1(n1264), .A2(n1193), .ZN(n1282) );
  NAND2_X2 U246 ( .A1(n1283), .A2(n1193), .ZN(n1281) );
  NAND2_X2 U247 ( .A1(n1284), .A2(n1164), .ZN(n1275) );
  NAND2_X2 U248 ( .A1(n1285), .A2(n1286), .ZN(B[3]) );
  MUX2_X1 U249 ( .A(n1287), .B(n1288), .S(n1184), .Z(n1286) );
  NAND2_X2 U250 ( .A1(n1172), .A2(n1237), .ZN(n1288) );
  NAND2_X2 U251 ( .A1(n1171), .A2(n1289), .ZN(n1287) );
  MUX2_X1 U252 ( .A(n1290), .B(n1291), .S(n1184), .Z(n1285) );
  NAND2_X2 U253 ( .A1(n1241), .A2(n1164), .ZN(n1291) );
  NAND2_X2 U254 ( .A1(n1292), .A2(n1293), .ZN(n1241) );
  MUX2_X1 U255 ( .A(n1294), .B(n1295), .S(n1190), .Z(n1293) );
  NAND2_X2 U256 ( .A1(n1208), .A2(n1264), .ZN(n1295) );
  NAND2_X2 U257 ( .A1(n1209), .A2(n1283), .ZN(n1294) );
  MUX2_X1 U258 ( .A(n1296), .B(n1297), .S(n1190), .Z(n1292) );
  NAND2_X2 U259 ( .A1(n1268), .A2(n1193), .ZN(n1297) );
  NAND2_X2 U260 ( .A1(n1298), .A2(n1193), .ZN(n1296) );
  OAI21_X2 U261 ( .B1(n1299), .B2(n1300), .A(n1164), .ZN(n1290) );
  MUX2_X1 U262 ( .A(n1301), .B(n1302), .S(n1190), .Z(n1300) );
  AND2_X2 U263 ( .A1(n1303), .A2(n1197), .ZN(n1302) );
  AND2_X2 U264 ( .A1(n1304), .A2(n1197), .ZN(n1301) );
  MUX2_X1 U265 ( .A(n1305), .B(n1306), .S(n1190), .Z(n1299) );
  AND2_X2 U266 ( .A1(n1210), .A2(n1307), .ZN(n1306) );
  AND2_X2 U267 ( .A1(n1211), .A2(n1308), .ZN(n1305) );
  AND3_X2 U268 ( .A1(n1186), .A2(n1165), .A3(n1309), .ZN(B[31]) );
  AND3_X2 U269 ( .A1(n1186), .A2(n1165), .A3(n1310), .ZN(B[30]) );
  NAND2_X2 U270 ( .A1(n1311), .A2(n1312), .ZN(B[2]) );
  MUX2_X1 U271 ( .A(n1313), .B(n1314), .S(n1184), .Z(n1312) );
  NAND2_X2 U272 ( .A1(n1171), .A2(n1247), .ZN(n1314) );
  NAND2_X2 U273 ( .A1(n1171), .A2(n1315), .ZN(n1313) );
  MUX2_X1 U274 ( .A(n1316), .B(n1317), .S(n1184), .Z(n1311) );
  NAND2_X2 U275 ( .A1(n1251), .A2(n1164), .ZN(n1317) );
  NAND2_X2 U276 ( .A1(n1318), .A2(n1319), .ZN(n1251) );
  MUX2_X1 U277 ( .A(n1320), .B(n1321), .S(n1190), .Z(n1319) );
  NAND2_X2 U278 ( .A1(n1209), .A2(n1268), .ZN(n1321) );
  INV_X2 U279 ( .A(n1322), .ZN(n1268) );
  MUX2_X1 U280 ( .A(n1323), .B(n1324), .S(n1176), .Z(n1322) );
  NAND2_X2 U281 ( .A1(n1208), .A2(n1298), .ZN(n1320) );
  MUX2_X1 U282 ( .A(n1325), .B(n1326), .S(n1190), .Z(n1318) );
  NAND2_X2 U283 ( .A1(n1283), .A2(n1193), .ZN(n1326) );
  NAND2_X2 U284 ( .A1(n1307), .A2(n1193), .ZN(n1325) );
  OAI21_X2 U285 ( .B1(n1327), .B2(n1328), .A(n1164), .ZN(n1316) );
  MUX2_X1 U286 ( .A(n1329), .B(n1330), .S(n1189), .Z(n1328) );
  AND2_X2 U287 ( .A1(n1308), .A2(n1197), .ZN(n1330) );
  AND2_X2 U288 ( .A1(n1331), .A2(n1197), .ZN(n1329) );
  MUX2_X1 U289 ( .A(n1332), .B(n1333), .S(n1189), .Z(n1327) );
  AND2_X2 U290 ( .A1(n1209), .A2(n1303), .ZN(n1333) );
  AND2_X2 U291 ( .A1(n1210), .A2(n1304), .ZN(n1332) );
  AND3_X2 U292 ( .A1(n1186), .A2(n1165), .A3(n1216), .ZN(B[29]) );
  AND3_X2 U293 ( .A1(n1186), .A2(n1165), .A3(n1226), .ZN(B[28]) );
  MUX2_X1 U294 ( .A(n1334), .B(n1335), .S(n1184), .Z(B[27]) );
  AND2_X2 U295 ( .A1(n1309), .A2(n1165), .ZN(n1335) );
  NOR2_X2 U296 ( .A1(n1169), .A2(n1336), .ZN(n1334) );
  MUX2_X1 U297 ( .A(n1337), .B(n1338), .S(n1184), .Z(B[26]) );
  AND2_X2 U298 ( .A1(n1310), .A2(n1165), .ZN(n1338) );
  NOR2_X2 U299 ( .A1(n1168), .A2(n1339), .ZN(n1337) );
  MUX2_X1 U300 ( .A(n1340), .B(n1341), .S(n1184), .Z(B[25]) );
  AND2_X2 U301 ( .A1(n1216), .A2(n1165), .ZN(n1341) );
  NOR2_X2 U302 ( .A1(n1169), .A2(n1342), .ZN(n1340) );
  MUX2_X1 U303 ( .A(n1343), .B(n1344), .S(n1184), .Z(B[24]) );
  NOR2_X2 U304 ( .A1(n1168), .A2(n1345), .ZN(n1344) );
  INV_X2 U305 ( .A(n1226), .ZN(n1345) );
  NOR2_X2 U306 ( .A1(n1167), .A2(n1346), .ZN(n1343) );
  MUX2_X1 U307 ( .A(n1347), .B(n1348), .S(n1184), .Z(B[23]) );
  NOR2_X2 U308 ( .A1(n1167), .A2(n1336), .ZN(n1348) );
  INV_X2 U309 ( .A(n1236), .ZN(n1336) );
  AND2_X2 U310 ( .A1(n1237), .A2(n1165), .ZN(n1347) );
  MUX2_X1 U311 ( .A(n1349), .B(n1350), .S(n1184), .Z(B[22]) );
  NOR2_X2 U312 ( .A1(n1168), .A2(n1339), .ZN(n1350) );
  INV_X2 U313 ( .A(n1246), .ZN(n1339) );
  AND2_X2 U314 ( .A1(n1247), .A2(n1165), .ZN(n1349) );
  MUX2_X1 U315 ( .A(n1351), .B(n1352), .S(n1184), .Z(B[21]) );
  NOR2_X2 U316 ( .A1(n1167), .A2(n1342), .ZN(n1352) );
  INV_X2 U317 ( .A(n1217), .ZN(n1342) );
  NAND2_X2 U318 ( .A1(n1353), .A2(n1354), .ZN(n1217) );
  MUX2_X1 U319 ( .A(n1355), .B(n1356), .S(n1189), .Z(n1354) );
  NAND2_X2 U320 ( .A1(n1357), .A2(n1198), .ZN(n1356) );
  NAND2_X2 U321 ( .A1(n1358), .A2(n1198), .ZN(n1355) );
  MUX2_X1 U322 ( .A(n1359), .B(n1360), .S(n1189), .Z(n1353) );
  NAND2_X2 U323 ( .A1(n1361), .A2(n1193), .ZN(n1360) );
  NAND2_X2 U324 ( .A1(n1362), .A2(n1193), .ZN(n1359) );
  AND2_X2 U325 ( .A1(n1256), .A2(n1165), .ZN(n1351) );
  MUX2_X1 U326 ( .A(n1363), .B(n1364), .S(n1184), .Z(B[20]) );
  NOR2_X2 U327 ( .A1(n1168), .A2(n1346), .ZN(n1364) );
  INV_X2 U328 ( .A(n1227), .ZN(n1346) );
  NAND2_X2 U329 ( .A1(n1365), .A2(n1366), .ZN(n1227) );
  MUX2_X1 U330 ( .A(n1367), .B(n1368), .S(n1189), .Z(n1366) );
  NAND2_X2 U331 ( .A1(n1361), .A2(n1199), .ZN(n1368) );
  NAND2_X2 U332 ( .A1(n1362), .A2(n1200), .ZN(n1367) );
  MUX2_X1 U333 ( .A(n1369), .B(n1370), .S(n1189), .Z(n1365) );
  NAND2_X2 U334 ( .A1(n1358), .A2(n1193), .ZN(n1370) );
  NAND2_X2 U335 ( .A1(n1371), .A2(n1193), .ZN(n1369) );
  AND2_X2 U336 ( .A1(n1274), .A2(n1165), .ZN(n1363) );
  NAND2_X2 U337 ( .A1(n1372), .A2(n1373), .ZN(B[1]) );
  MUX2_X1 U338 ( .A(n1374), .B(n1375), .S(n1184), .Z(n1373) );
  NAND2_X2 U339 ( .A1(n1170), .A2(n1256), .ZN(n1375) );
  NAND2_X2 U340 ( .A1(n1170), .A2(n1376), .ZN(n1374) );
  MUX2_X1 U341 ( .A(n1377), .B(n1378), .S(n1183), .Z(n1372) );
  NAND2_X2 U342 ( .A1(n1269), .A2(n1164), .ZN(n1378) );
  NAND2_X2 U343 ( .A1(n1379), .A2(n1380), .ZN(n1269) );
  MUX2_X1 U344 ( .A(n1381), .B(n1382), .S(n1189), .Z(n1380) );
  NAND2_X2 U345 ( .A1(n1208), .A2(n1283), .ZN(n1382) );
  INV_X2 U346 ( .A(n1383), .ZN(n1283) );
  MUX2_X1 U347 ( .A(n1384), .B(n1385), .S(n1176), .Z(n1383) );
  NAND2_X2 U348 ( .A1(n1207), .A2(n1307), .ZN(n1381) );
  MUX2_X1 U349 ( .A(n1386), .B(n1387), .S(n1189), .Z(n1379) );
  NAND2_X2 U350 ( .A1(n1298), .A2(n1193), .ZN(n1387) );
  NAND2_X2 U351 ( .A1(n1303), .A2(n1194), .ZN(n1386) );
  OAI21_X2 U352 ( .B1(n1388), .B2(n1389), .A(n1164), .ZN(n1377) );
  MUX2_X1 U353 ( .A(n1390), .B(n1391), .S(n1189), .Z(n1389) );
  AND2_X2 U354 ( .A1(n1304), .A2(n1197), .ZN(n1391) );
  AND2_X2 U355 ( .A1(n1392), .A2(n1197), .ZN(n1390) );
  MUX2_X1 U356 ( .A(n1393), .B(n1394), .S(n1189), .Z(n1388) );
  AND2_X2 U357 ( .A1(n1208), .A2(n1308), .ZN(n1394) );
  AND2_X2 U358 ( .A1(n1210), .A2(n1331), .ZN(n1393) );
  MUX2_X1 U359 ( .A(n1395), .B(n1396), .S(n1183), .Z(B[19]) );
  AND2_X2 U360 ( .A1(n1237), .A2(n1165), .ZN(n1396) );
  NAND2_X2 U361 ( .A1(n1397), .A2(n1398), .ZN(n1237) );
  MUX2_X1 U362 ( .A(n1399), .B(n1400), .S(n1189), .Z(n1398) );
  NAND2_X2 U363 ( .A1(n1358), .A2(n1199), .ZN(n1400) );
  NAND2_X2 U364 ( .A1(n1371), .A2(n1201), .ZN(n1399) );
  MUX2_X1 U365 ( .A(n1401), .B(n1402), .S(n1189), .Z(n1397) );
  NAND2_X2 U366 ( .A1(n1362), .A2(n1194), .ZN(n1402) );
  NAND2_X2 U367 ( .A1(n1403), .A2(n1194), .ZN(n1401) );
  AND2_X2 U368 ( .A1(n1289), .A2(n1165), .ZN(n1395) );
  MUX2_X1 U369 ( .A(n1404), .B(n1405), .S(n1183), .Z(B[18]) );
  AND2_X2 U370 ( .A1(n1247), .A2(n1165), .ZN(n1405) );
  NAND2_X2 U371 ( .A1(n1406), .A2(n1407), .ZN(n1247) );
  MUX2_X1 U372 ( .A(n1408), .B(n1409), .S(n1189), .Z(n1407) );
  NAND2_X2 U373 ( .A1(n1362), .A2(n1198), .ZN(n1409) );
  INV_X2 U374 ( .A(n1410), .ZN(n1362) );
  NAND2_X2 U375 ( .A1(n1208), .A2(n1403), .ZN(n1408) );
  MUX2_X1 U376 ( .A(n1411), .B(n1412), .S(n1189), .Z(n1406) );
  NAND2_X2 U377 ( .A1(n1371), .A2(n1194), .ZN(n1412) );
  NAND2_X2 U378 ( .A1(n1413), .A2(n1194), .ZN(n1411) );
  AND2_X2 U379 ( .A1(n1315), .A2(n1165), .ZN(n1404) );
  MUX2_X1 U380 ( .A(n1414), .B(n1415), .S(n1183), .Z(B[17]) );
  AND2_X2 U381 ( .A1(n1256), .A2(n1165), .ZN(n1415) );
  NAND2_X2 U382 ( .A1(n1416), .A2(n1417), .ZN(n1256) );
  MUX2_X1 U383 ( .A(n1418), .B(n1419), .S(n1189), .Z(n1417) );
  NAND2_X2 U384 ( .A1(n1371), .A2(n1200), .ZN(n1419) );
  INV_X2 U385 ( .A(n1420), .ZN(n1371) );
  NAND2_X2 U386 ( .A1(n1207), .A2(n1413), .ZN(n1418) );
  MUX2_X1 U387 ( .A(n1421), .B(n1422), .S(n1189), .Z(n1416) );
  NAND2_X2 U388 ( .A1(n1403), .A2(n1194), .ZN(n1422) );
  NAND2_X2 U389 ( .A1(n1423), .A2(n1194), .ZN(n1421) );
  AND2_X2 U390 ( .A1(n1376), .A2(n1165), .ZN(n1414) );
  MUX2_X1 U391 ( .A(n1424), .B(n1425), .S(n1183), .Z(B[16]) );
  AND2_X2 U392 ( .A1(n1274), .A2(n1165), .ZN(n1425) );
  AND2_X2 U393 ( .A1(n1426), .A2(n1165), .ZN(n1424) );
  NAND2_X2 U394 ( .A1(n1427), .A2(n1428), .ZN(B[15]) );
  NAND3_X1 U395 ( .A1(n1186), .A2(n1165), .A3(n1429), .ZN(n1428) );
  MUX2_X1 U396 ( .A(n1430), .B(n1431), .S(n1169), .Z(n1427) );
  NAND2_X2 U397 ( .A1(n1309), .A2(n1186), .ZN(n1431) );
  NAND2_X2 U398 ( .A1(n1183), .A2(n1289), .ZN(n1430) );
  NAND2_X2 U399 ( .A1(n1432), .A2(n1433), .ZN(n1289) );
  MUX2_X1 U400 ( .A(n1434), .B(n1435), .S(n1189), .Z(n1433) );
  NAND2_X2 U401 ( .A1(n1207), .A2(n1413), .ZN(n1435) );
  NAND2_X2 U402 ( .A1(n1206), .A2(n1436), .ZN(n1434) );
  MUX2_X1 U403 ( .A(n1437), .B(n1438), .S(n1188), .Z(n1432) );
  NAND2_X2 U404 ( .A1(n1423), .A2(n1194), .ZN(n1438) );
  NAND2_X2 U405 ( .A1(n1439), .A2(n1194), .ZN(n1437) );
  NAND2_X2 U406 ( .A1(n1440), .A2(n1441), .ZN(B[14]) );
  NAND3_X1 U407 ( .A1(n1186), .A2(n1166), .A3(n1442), .ZN(n1441) );
  MUX2_X1 U408 ( .A(n1443), .B(n1444), .S(n1172), .Z(n1440) );
  NAND2_X2 U409 ( .A1(n1310), .A2(n1186), .ZN(n1444) );
  NAND2_X2 U410 ( .A1(n1183), .A2(n1315), .ZN(n1443) );
  NAND2_X2 U411 ( .A1(n1445), .A2(n1446), .ZN(n1315) );
  MUX2_X1 U412 ( .A(n1447), .B(n1448), .S(n1188), .Z(n1446) );
  NAND2_X2 U413 ( .A1(n1207), .A2(n1423), .ZN(n1448) );
  NAND2_X2 U414 ( .A1(n1206), .A2(n1439), .ZN(n1447) );
  MUX2_X1 U415 ( .A(n1449), .B(n1450), .S(n1188), .Z(n1445) );
  NAND2_X2 U416 ( .A1(n1436), .A2(n1194), .ZN(n1450) );
  NAND2_X2 U417 ( .A1(n1451), .A2(n1194), .ZN(n1449) );
  NAND2_X2 U418 ( .A1(n1452), .A2(n1453), .ZN(B[13]) );
  NAND3_X1 U419 ( .A1(n1186), .A2(n1166), .A3(n1220), .ZN(n1453) );
  NAND2_X2 U420 ( .A1(n1454), .A2(n1455), .ZN(n1220) );
  MUX2_X1 U421 ( .A(n1456), .B(n1457), .S(n1188), .Z(n1455) );
  NAND2_X2 U422 ( .A1(n1206), .A2(n1458), .ZN(n1457) );
  NAND2_X2 U423 ( .A1(n1206), .A2(n1459), .ZN(n1456) );
  MUX2_X1 U424 ( .A(n1460), .B(n1461), .S(n1188), .Z(n1454) );
  NAND2_X2 U425 ( .A1(n1462), .A2(n1194), .ZN(n1461) );
  NAND2_X2 U426 ( .A1(n1463), .A2(n1195), .ZN(n1460) );
  MUX2_X1 U427 ( .A(n1464), .B(n1465), .S(n1170), .Z(n1452) );
  NAND2_X2 U428 ( .A1(n1216), .A2(n1186), .ZN(n1465) );
  NAND2_X2 U429 ( .A1(n1466), .A2(n1467), .ZN(n1216) );
  NAND3_X1 U430 ( .A1(n1197), .A2(n1192), .A3(n1468), .ZN(n1467) );
  MUX2_X1 U431 ( .A(n1469), .B(n1470), .S(n1201), .Z(n1466) );
  NAND2_X2 U432 ( .A1(n1471), .A2(n1191), .ZN(n1470) );
  NAND2_X2 U433 ( .A1(n1187), .A2(n1472), .ZN(n1469) );
  NAND2_X2 U434 ( .A1(n1183), .A2(n1376), .ZN(n1464) );
  NAND2_X2 U435 ( .A1(n1473), .A2(n1474), .ZN(n1376) );
  MUX2_X1 U436 ( .A(n1475), .B(n1476), .S(n1188), .Z(n1474) );
  NAND2_X2 U437 ( .A1(n1205), .A2(n1436), .ZN(n1476) );
  NAND2_X2 U438 ( .A1(n1205), .A2(n1451), .ZN(n1475) );
  MUX2_X1 U439 ( .A(n1477), .B(n1478), .S(n1188), .Z(n1473) );
  NAND2_X2 U440 ( .A1(n1439), .A2(n1195), .ZN(n1478) );
  NAND2_X2 U441 ( .A1(n1479), .A2(n1195), .ZN(n1477) );
  NAND2_X2 U442 ( .A1(n1480), .A2(n1481), .ZN(B[12]) );
  NAND3_X1 U443 ( .A1(n1186), .A2(n1166), .A3(n1230), .ZN(n1481) );
  NAND2_X2 U444 ( .A1(n1482), .A2(n1483), .ZN(n1230) );
  MUX2_X1 U445 ( .A(n1484), .B(n1485), .S(n1188), .Z(n1483) );
  NAND2_X2 U446 ( .A1(n1205), .A2(n1462), .ZN(n1485) );
  NAND2_X2 U447 ( .A1(n1204), .A2(n1463), .ZN(n1484) );
  MUX2_X1 U448 ( .A(n1486), .B(n1487), .S(n1188), .Z(n1482) );
  NAND2_X2 U449 ( .A1(n1459), .A2(n1195), .ZN(n1487) );
  NAND2_X2 U450 ( .A1(n1263), .A2(n1195), .ZN(n1486) );
  MUX2_X1 U451 ( .A(n1488), .B(n1489), .S(n1171), .Z(n1480) );
  NAND2_X2 U452 ( .A1(n1226), .A2(n1186), .ZN(n1489) );
  NAND2_X2 U453 ( .A1(n1490), .A2(n1491), .ZN(n1226) );
  MUX2_X1 U454 ( .A(n1492), .B(n1493), .S(n1188), .Z(n1491) );
  NAND2_X2 U455 ( .A1(n1472), .A2(n1199), .ZN(n1493) );
  NAND2_X2 U456 ( .A1(n1468), .A2(n1200), .ZN(n1492) );
  MUX2_X1 U457 ( .A(n1494), .B(n1495), .S(n1188), .Z(n1490) );
  NAND2_X2 U458 ( .A1(n1471), .A2(n1195), .ZN(n1495) );
  NAND2_X2 U459 ( .A1(n1357), .A2(n1195), .ZN(n1494) );
  NAND2_X2 U460 ( .A1(n1183), .A2(n1426), .ZN(n1488) );
  NAND2_X2 U461 ( .A1(n1496), .A2(n1497), .ZN(B[11]) );
  MUX2_X1 U462 ( .A(n1498), .B(n1499), .S(n1183), .Z(n1497) );
  NAND2_X2 U463 ( .A1(n1309), .A2(n1167), .ZN(n1499) );
  INV_X2 U464 ( .A(n1500), .ZN(n1309) );
  NAND3_X1 U465 ( .A1(n1197), .A2(n1192), .A3(n1472), .ZN(n1500) );
  NAND2_X2 U466 ( .A1(n1170), .A2(n1236), .ZN(n1498) );
  NAND2_X2 U467 ( .A1(n1501), .A2(n1502), .ZN(n1236) );
  MUX2_X1 U468 ( .A(n1503), .B(n1504), .S(n1188), .Z(n1502) );
  NAND2_X2 U469 ( .A1(n1205), .A2(n1471), .ZN(n1504) );
  NAND2_X2 U470 ( .A1(n1357), .A2(n1200), .ZN(n1503) );
  MUX2_X1 U471 ( .A(n1505), .B(n1506), .S(n1188), .Z(n1501) );
  NAND2_X2 U472 ( .A1(n1468), .A2(n1195), .ZN(n1506) );
  NAND2_X2 U473 ( .A1(n1361), .A2(n1195), .ZN(n1505) );
  MUX2_X1 U474 ( .A(n1507), .B(n1508), .S(n1183), .Z(n1496) );
  NAND2_X2 U475 ( .A1(n1429), .A2(n1163), .ZN(n1508) );
  NAND2_X2 U476 ( .A1(n1509), .A2(n1510), .ZN(n1429) );
  MUX2_X1 U477 ( .A(n1511), .B(n1512), .S(n1188), .Z(n1510) );
  NAND2_X2 U478 ( .A1(n1204), .A2(n1451), .ZN(n1512) );
  NAND2_X2 U479 ( .A1(n1202), .A2(n1458), .ZN(n1511) );
  MUX2_X1 U480 ( .A(n1513), .B(n1514), .S(n1188), .Z(n1509) );
  NAND2_X2 U481 ( .A1(n1479), .A2(n1196), .ZN(n1514) );
  NAND2_X2 U482 ( .A1(n1462), .A2(n1195), .ZN(n1513) );
  NAND2_X2 U483 ( .A1(n1240), .A2(n1163), .ZN(n1507) );
  NAND2_X2 U484 ( .A1(n1515), .A2(n1516), .ZN(n1240) );
  MUX2_X1 U485 ( .A(n1517), .B(n1518), .S(n1187), .Z(n1516) );
  NAND2_X2 U486 ( .A1(n1204), .A2(n1459), .ZN(n1518) );
  NAND2_X2 U487 ( .A1(n1202), .A2(n1263), .ZN(n1517) );
  MUX2_X1 U488 ( .A(n1519), .B(n1520), .S(n1188), .Z(n1515) );
  NAND2_X2 U489 ( .A1(n1463), .A2(n1196), .ZN(n1520) );
  NAND2_X2 U490 ( .A1(n1267), .A2(n1195), .ZN(n1519) );
  NAND2_X2 U491 ( .A1(n1521), .A2(n1522), .ZN(B[10]) );
  MUX2_X1 U492 ( .A(n1523), .B(n1524), .S(n1183), .Z(n1522) );
  NAND2_X2 U493 ( .A1(n1170), .A2(n1310), .ZN(n1524) );
  MUX2_X1 U494 ( .A(n1525), .B(n1526), .S(n1202), .Z(n1310) );
  INV_X2 U495 ( .A(n1527), .ZN(n1526) );
  NAND2_X2 U496 ( .A1(n1472), .A2(n1191), .ZN(n1527) );
  INV_X2 U497 ( .A(n1528), .ZN(n1472) );
  INV_X2 U498 ( .A(n1529), .ZN(n1525) );
  NAND2_X2 U499 ( .A1(n1471), .A2(n1191), .ZN(n1529) );
  INV_X2 U500 ( .A(n1530), .ZN(n1471) );
  NAND2_X2 U501 ( .A1(n1169), .A2(n1246), .ZN(n1523) );
  NAND2_X2 U502 ( .A1(n1531), .A2(n1532), .ZN(n1246) );
  MUX2_X1 U503 ( .A(n1533), .B(n1534), .S(n1187), .Z(n1532) );
  NAND2_X2 U504 ( .A1(n1468), .A2(n1198), .ZN(n1534) );
  INV_X2 U505 ( .A(n1535), .ZN(n1468) );
  NAND2_X2 U506 ( .A1(n1361), .A2(n1199), .ZN(n1533) );
  INV_X2 U507 ( .A(n1536), .ZN(n1361) );
  MUX2_X1 U508 ( .A(n1537), .B(n1538), .S(n1187), .Z(n1531) );
  NAND2_X2 U509 ( .A1(n1357), .A2(n1196), .ZN(n1538) );
  INV_X2 U510 ( .A(n1539), .ZN(n1357) );
  NAND2_X2 U511 ( .A1(n1358), .A2(n1196), .ZN(n1537) );
  INV_X2 U512 ( .A(n1540), .ZN(n1358) );
  NAND2_X2 U513 ( .A1(A[26]), .A2(n1181), .ZN(n1540) );
  MUX2_X1 U514 ( .A(n1541), .B(n1542), .S(n1183), .Z(n1521) );
  NAND2_X2 U515 ( .A1(n1442), .A2(n1163), .ZN(n1542) );
  NAND2_X2 U516 ( .A1(n1543), .A2(n1544), .ZN(n1442) );
  MUX2_X1 U517 ( .A(n1545), .B(n1546), .S(n1187), .Z(n1544) );
  NAND2_X2 U518 ( .A1(n1204), .A2(n1479), .ZN(n1546) );
  NAND2_X2 U519 ( .A1(n1202), .A2(n1462), .ZN(n1545) );
  INV_X2 U520 ( .A(n1547), .ZN(n1462) );
  MUX2_X1 U521 ( .A(n1548), .B(n1549), .S(n1176), .Z(n1547) );
  MUX2_X1 U522 ( .A(n1550), .B(n1551), .S(n1187), .Z(n1543) );
  NAND2_X2 U523 ( .A1(n1458), .A2(n1196), .ZN(n1551) );
  NAND2_X2 U524 ( .A1(n1459), .A2(n1196), .ZN(n1550) );
  INV_X2 U525 ( .A(n1552), .ZN(n1459) );
  MUX2_X1 U526 ( .A(n1553), .B(n1554), .S(n1176), .Z(n1552) );
  NAND2_X2 U527 ( .A1(n1250), .A2(n1163), .ZN(n1541) );
  NAND2_X2 U528 ( .A1(n1555), .A2(n1556), .ZN(n1250) );
  MUX2_X1 U529 ( .A(n1557), .B(n1558), .S(n1187), .Z(n1556) );
  NAND2_X2 U530 ( .A1(n1203), .A2(n1463), .ZN(n1558) );
  INV_X2 U531 ( .A(n1559), .ZN(n1463) );
  MUX2_X1 U532 ( .A(n1560), .B(n1561), .S(n1176), .Z(n1559) );
  NAND2_X2 U533 ( .A1(n1202), .A2(n1267), .ZN(n1557) );
  INV_X2 U534 ( .A(n1562), .ZN(n1267) );
  MUX2_X1 U535 ( .A(n1563), .B(n1564), .S(n1176), .Z(n1562) );
  MUX2_X1 U536 ( .A(n1565), .B(n1566), .S(n1187), .Z(n1555) );
  NAND2_X2 U537 ( .A1(n1263), .A2(n1196), .ZN(n1566) );
  INV_X2 U538 ( .A(n1567), .ZN(n1263) );
  MUX2_X1 U539 ( .A(n1568), .B(n1569), .S(n1176), .Z(n1567) );
  NAND2_X2 U540 ( .A1(n1264), .A2(n1196), .ZN(n1565) );
  INV_X2 U541 ( .A(n1570), .ZN(n1264) );
  MUX2_X1 U542 ( .A(n1571), .B(n1572), .S(n1176), .Z(n1570) );
  NAND2_X2 U543 ( .A1(n1573), .A2(n1574), .ZN(B[0]) );
  MUX2_X1 U544 ( .A(n1575), .B(n1576), .S(n1183), .Z(n1574) );
  NAND2_X2 U545 ( .A1(n1169), .A2(n1274), .ZN(n1576) );
  NAND2_X2 U546 ( .A1(n1577), .A2(n1578), .ZN(n1274) );
  MUX2_X1 U547 ( .A(n1579), .B(n1580), .S(n1187), .Z(n1578) );
  NAND2_X2 U548 ( .A1(n1203), .A2(n1403), .ZN(n1580) );
  INV_X2 U549 ( .A(n1581), .ZN(n1403) );
  MUX2_X1 U550 ( .A(n1549), .B(n1582), .S(n1176), .Z(n1581) );
  INV_X2 U551 ( .A(A[23]), .ZN(n1549) );
  NAND2_X2 U552 ( .A1(n1201), .A2(n1423), .ZN(n1579) );
  INV_X2 U553 ( .A(n1583), .ZN(n1423) );
  MUX2_X1 U554 ( .A(n1561), .B(n1584), .S(n1176), .Z(n1583) );
  MUX2_X1 U555 ( .A(n1585), .B(n1586), .S(n1187), .Z(n1577) );
  NAND2_X2 U556 ( .A1(n1413), .A2(n1196), .ZN(n1586) );
  INV_X2 U557 ( .A(n1587), .ZN(n1413) );
  MUX2_X1 U558 ( .A(n1554), .B(n1588), .S(n1176), .Z(n1587) );
  NAND2_X2 U559 ( .A1(n1436), .A2(n1196), .ZN(n1585) );
  INV_X2 U560 ( .A(n1589), .ZN(n1436) );
  MUX2_X1 U561 ( .A(n1569), .B(n1590), .S(n1176), .Z(n1589) );
  NAND2_X2 U562 ( .A1(n1171), .A2(n1426), .ZN(n1575) );
  NAND2_X2 U563 ( .A1(n1591), .A2(n1592), .ZN(n1426) );
  MUX2_X1 U564 ( .A(n1593), .B(n1594), .S(n1187), .Z(n1592) );
  NAND2_X2 U565 ( .A1(n1203), .A2(n1439), .ZN(n1594) );
  INV_X2 U566 ( .A(n1595), .ZN(n1439) );
  MUX2_X1 U567 ( .A(n1564), .B(n1596), .S(n1177), .Z(n1595) );
  NAND2_X2 U568 ( .A1(n1201), .A2(n1479), .ZN(n1593) );
  INV_X2 U569 ( .A(n1597), .ZN(n1479) );
  MUX2_X1 U570 ( .A(n1324), .B(n1598), .S(n1177), .Z(n1597) );
  MUX2_X1 U571 ( .A(n1599), .B(n1600), .S(n1187), .Z(n1591) );
  NAND2_X2 U572 ( .A1(n1451), .A2(n1197), .ZN(n1600) );
  INV_X2 U573 ( .A(n1601), .ZN(n1451) );
  MUX2_X1 U574 ( .A(n1572), .B(n1602), .S(n1177), .Z(n1601) );
  INV_X2 U575 ( .A(A[26]), .ZN(n1602) );
  NAND2_X2 U576 ( .A1(n1458), .A2(n1196), .ZN(n1599) );
  INV_X2 U577 ( .A(n1603), .ZN(n1458) );
  MUX2_X1 U578 ( .A(n1385), .B(n1604), .S(n1177), .Z(n1603) );
  MUX2_X1 U579 ( .A(n1605), .B(n1606), .S(n1184), .Z(n1573) );
  NAND2_X2 U580 ( .A1(n1284), .A2(n1163), .ZN(n1606) );
  NAND2_X2 U581 ( .A1(n1607), .A2(n1608), .ZN(n1284) );
  MUX2_X1 U582 ( .A(n1609), .B(n1610), .S(n1187), .Z(n1608) );
  NAND2_X2 U583 ( .A1(n1203), .A2(n1298), .ZN(n1610) );
  INV_X2 U584 ( .A(n1611), .ZN(n1298) );
  MUX2_X1 U585 ( .A(n1612), .B(n1548), .S(n1177), .Z(n1611) );
  NAND2_X2 U586 ( .A1(n1201), .A2(n1303), .ZN(n1609) );
  INV_X2 U587 ( .A(n1613), .ZN(n1303) );
  MUX2_X1 U588 ( .A(n1614), .B(n1560), .S(n1177), .Z(n1613) );
  MUX2_X1 U589 ( .A(n1615), .B(n1616), .S(n1187), .Z(n1607) );
  NAND2_X2 U590 ( .A1(n1307), .A2(n1197), .ZN(n1616) );
  INV_X2 U591 ( .A(n1617), .ZN(n1307) );
  MUX2_X1 U592 ( .A(n1618), .B(n1553), .S(n1177), .Z(n1617) );
  NAND2_X2 U593 ( .A1(n1308), .A2(n1196), .ZN(n1615) );
  INV_X2 U594 ( .A(n1619), .ZN(n1308) );
  MUX2_X1 U595 ( .A(n1620), .B(n1568), .S(n1177), .Z(n1619) );
  OAI21_X2 U596 ( .B1(n1621), .B2(n1622), .A(n1164), .ZN(n1605) );
  MUX2_X1 U597 ( .A(n1623), .B(n1624), .S(n1187), .Z(n1622) );
  AND2_X2 U598 ( .A1(n1331), .A2(n1197), .ZN(n1624) );
  INV_X2 U599 ( .A(n1625), .ZN(n1331) );
  MUX2_X1 U600 ( .A(n1626), .B(n1571), .S(n1177), .Z(n1625) );
  AND2_X2 U601 ( .A1(n1627), .A2(n1197), .ZN(n1623) );
  MUX2_X1 U602 ( .A(A[0]), .B(A[8]), .S(n1177), .Z(n1627) );
  MUX2_X1 U603 ( .A(n1628), .B(n1629), .S(n1188), .Z(n1621) );
  AND2_X2 U604 ( .A1(n1211), .A2(n1304), .ZN(n1629) );
  INV_X2 U605 ( .A(n1630), .ZN(n1304) );
  MUX2_X1 U606 ( .A(n1631), .B(n1563), .S(n1177), .Z(n1630) );
  INV_X2 U607 ( .A(A[3]), .ZN(n1631) );
  AND2_X2 U608 ( .A1(n1210), .A2(n1392), .ZN(n1628) );
  INV_X2 U609 ( .A(n1632), .ZN(n1392) );
  MUX2_X1 U610 ( .A(n1633), .B(n1323), .S(n1177), .Z(n1632) );
endmodule


module Xi_core_DW01_add_3 ( A, B, SUM, CI, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n56, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n105, n106, n107, n108, n110, n111, n112, n113,
         n114, n115, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n130, n131, n132, n133, n134, n135, n138, n139, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157,
         n158, n159, n160, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n191, n192, n193, n194, n195,
         n196, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n213, n214, n215, n216, n217, n218, n219, n220,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n235, n236, n237, n238, n239, n240, n242, n243, n244, n245, n246,
         n247, n248, n249, n252, n253, n254, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n285, n286, n287, n288, n289,
         n290, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n329, n331,
         n332, n333, n334, n335, n336, n340, n342, n343, n345, n347, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n391, n392, n393, n394, n395, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520;

  NAND2_X4 U6 ( .A1(n364), .A2(n38), .ZN(n5) );
  NAND2_X4 U20 ( .A1(n46), .A2(n49), .ZN(n6) );
  AOI21_X4 U35 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NAND2_X4 U38 ( .A1(n61), .A2(n64), .ZN(n7) );
  XNOR2_X2 U42 ( .A(n74), .B(n8), .ZN(SUM[28]) );
  NAND2_X4 U50 ( .A1(n70), .A2(n73), .ZN(n8) );
  XNOR2_X2 U54 ( .A(n87), .B(n9), .ZN(SUM[27]) );
  NAND2_X4 U66 ( .A1(n83), .A2(n86), .ZN(n9) );
  XNOR2_X2 U70 ( .A(n96), .B(n10), .ZN(SUM[26]) );
  NAND2_X4 U78 ( .A1(n369), .A2(n95), .ZN(n10) );
  XNOR2_X2 U82 ( .A(n113), .B(n11), .ZN(SUM[25]) );
  NAND2_X4 U84 ( .A1(n391), .A2(n99), .ZN(n97) );
  AOI21_X4 U85 ( .B1(n347), .B2(n99), .A(n100), .ZN(n98) );
  AOI21_X4 U95 ( .B1(n370), .B2(n119), .A(n110), .ZN(n108) );
  NAND2_X4 U98 ( .A1(n370), .A2(n112), .ZN(n11) );
  XNOR2_X2 U102 ( .A(n122), .B(n12), .ZN(SUM[24]) );
  XNOR2_X2 U114 ( .A(n133), .B(n13), .ZN(SUM[23]) );
  NOR2_X4 U118 ( .A1(n4), .A2(n127), .ZN(n125) );
  NAND2_X4 U124 ( .A1(n372), .A2(n132), .ZN(n13) );
  XNOR2_X2 U128 ( .A(n146), .B(n14), .ZN(SUM[22]) );
  NOR2_X4 U138 ( .A1(n151), .A2(n144), .ZN(n138) );
  NAND2_X4 U140 ( .A1(n373), .A2(n145), .ZN(n14) );
  XNOR2_X2 U144 ( .A(n157), .B(n15), .ZN(SUM[21]) );
  NAND2_X4 U146 ( .A1(n391), .A2(n149), .ZN(n147) );
  AOI21_X4 U147 ( .B1(n347), .B2(n149), .A(n150), .ZN(n148) );
  NAND2_X4 U154 ( .A1(n374), .A2(n156), .ZN(n15) );
  XNOR2_X2 U158 ( .A(n174), .B(n16), .ZN(SUM[20]) );
  NAND2_X4 U174 ( .A1(n375), .A2(n173), .ZN(n16) );
  XNOR2_X2 U178 ( .A(n181), .B(n17), .ZN(SUM[19]) );
  NAND2_X4 U180 ( .A1(n184), .A2(n376), .ZN(n175) );
  AOI21_X4 U181 ( .B1(n185), .B2(n376), .A(n178), .ZN(n176) );
  NAND2_X4 U184 ( .A1(n376), .A2(n180), .ZN(n17) );
  XNOR2_X2 U188 ( .A(n194), .B(n18), .ZN(SUM[18]) );
  NOR2_X4 U192 ( .A1(n4), .A2(n186), .ZN(n184) );
  NAND2_X4 U200 ( .A1(n377), .A2(n193), .ZN(n18) );
  XNOR2_X2 U204 ( .A(n201), .B(n19), .ZN(SUM[17]) );
  NAND2_X4 U206 ( .A1(n204), .A2(n378), .ZN(n195) );
  AOI21_X4 U207 ( .B1(n205), .B2(n378), .A(n198), .ZN(n196) );
  NAND2_X4 U210 ( .A1(n378), .A2(n200), .ZN(n19) );
  XNOR2_X2 U214 ( .A(n218), .B(n20), .ZN(SUM[16]) );
  NOR2_X4 U218 ( .A1(n4), .A2(n206), .ZN(n204) );
  NAND2_X4 U230 ( .A1(n379), .A2(n217), .ZN(n20) );
  XNOR2_X2 U234 ( .A(n225), .B(n21), .ZN(SUM[15]) );
  NAND2_X4 U236 ( .A1(n228), .A2(n380), .ZN(n219) );
  AOI21_X4 U237 ( .B1(n229), .B2(n380), .A(n222), .ZN(n220) );
  NAND2_X4 U240 ( .A1(n380), .A2(n224), .ZN(n21) );
  XNOR2_X2 U244 ( .A(n238), .B(n22), .ZN(SUM[14]) );
  NOR2_X4 U248 ( .A1(n4), .A2(n230), .ZN(n228) );
  NAND2_X4 U256 ( .A1(n381), .A2(n237), .ZN(n22) );
  XNOR2_X2 U260 ( .A(n245), .B(n23), .ZN(SUM[13]) );
  NAND2_X4 U262 ( .A1(n248), .A2(n382), .ZN(n239) );
  AOI21_X4 U263 ( .B1(n249), .B2(n382), .A(n242), .ZN(n240) );
  NAND2_X4 U266 ( .A1(n382), .A2(n244), .ZN(n23) );
  XNOR2_X2 U270 ( .A(n268), .B(n24), .ZN(SUM[12]) );
  NAND2_X4 U292 ( .A1(n383), .A2(n267), .ZN(n24) );
  XNOR2_X2 U296 ( .A(n275), .B(n25), .ZN(SUM[11]) );
  NAND2_X4 U298 ( .A1(n278), .A2(n384), .ZN(n269) );
  AOI21_X4 U299 ( .B1(n279), .B2(n384), .A(n272), .ZN(n270) );
  XNOR2_X2 U306 ( .A(n288), .B(n26), .ZN(SUM[10]) );
  NOR2_X4 U310 ( .A1(n4), .A2(n280), .ZN(n278) );
  NAND2_X4 U318 ( .A1(n385), .A2(n287), .ZN(n26) );
  XNOR2_X2 U322 ( .A(n295), .B(n27), .ZN(SUM[9]) );
  NAND2_X4 U324 ( .A1(n298), .A2(n386), .ZN(n289) );
  AOI21_X4 U325 ( .B1(n299), .B2(n386), .A(n292), .ZN(n290) );
  XNOR2_X2 U332 ( .A(n314), .B(n28), .ZN(SUM[8]) );
  NOR2_X4 U336 ( .A1(n4), .A2(n300), .ZN(n298) );
  NOR2_X4 U344 ( .A1(n308), .A2(n326), .ZN(n302) );
  NAND2_X4 U350 ( .A1(n387), .A2(n313), .ZN(n28) );
  XNOR2_X2 U354 ( .A(n321), .B(n29), .ZN(SUM[7]) );
  NAND2_X4 U356 ( .A1(n324), .A2(n388), .ZN(n315) );
  AOI21_X4 U357 ( .B1(n325), .B2(n388), .A(n318), .ZN(n316) );
  XNOR2_X2 U364 ( .A(n334), .B(n30), .ZN(SUM[6]) );
  NOR2_X4 U368 ( .A1(n4), .A2(n326), .ZN(n324) );
  XNOR2_X2 U380 ( .A(n343), .B(n31), .ZN(SUM[5]) );
  XNOR2_X2 U402 ( .A(n355), .B(n33), .ZN(SUM[3]) );
  AOI21_X4 U403 ( .B1(n351), .B2(n359), .A(n352), .ZN(n2) );
  NOR2_X4 U404 ( .A1(n356), .A2(n353), .ZN(n351) );
  OAI21_X4 U405 ( .B1(n357), .B2(n353), .A(n354), .ZN(n352) );
  NAND2_X4 U406 ( .A1(n392), .A2(n354), .ZN(n33) );
  XOR2_X2 U410 ( .A(n34), .B(n358), .Z(SUM[2]) );
  OAI21_X4 U411 ( .B1(n358), .B2(n356), .A(n357), .ZN(n355) );
  NAND2_X4 U412 ( .A1(n393), .A2(n357), .ZN(n34) );
  XOR2_X2 U416 ( .A(n35), .B(n363), .Z(SUM[1]) );
  OAI21_X4 U418 ( .B1(n360), .B2(n363), .A(n361), .ZN(n359) );
  NAND2_X4 U419 ( .A1(n394), .A2(n361), .ZN(n35) );
  NAND2_X4 U424 ( .A1(n395), .A2(n363), .ZN(n36) );
  NAND2_X1 U431 ( .A1(n391), .A2(n345), .ZN(n32) );
  OAI21_X1 U432 ( .B1(n345), .B2(n127), .A(n128), .ZN(n126) );
  OAI21_X1 U433 ( .B1(n345), .B2(n206), .A(n207), .ZN(n205) );
  OAI21_X1 U434 ( .B1(n345), .B2(n280), .A(n281), .ZN(n279) );
  OAI21_X1 U435 ( .B1(n345), .B2(n230), .A(n231), .ZN(n229) );
  OAI21_X1 U436 ( .B1(n345), .B2(n300), .A(n301), .ZN(n299) );
  OAI21_X1 U437 ( .B1(n345), .B2(n186), .A(n187), .ZN(n185) );
  INV_X1 U438 ( .A(n345), .ZN(n347) );
  AOI21_X1 U439 ( .B1(n163), .B2(n374), .A(n154), .ZN(n152) );
  NOR2_X2 U440 ( .A1(n179), .A2(n172), .ZN(n170) );
  NOR2_X2 U441 ( .A1(n223), .A2(n216), .ZN(n214) );
  NOR2_X2 U442 ( .A1(A[16]), .A2(B[16]), .ZN(n216) );
  NOR2_X1 U443 ( .A1(n236), .A2(n243), .ZN(n498) );
  NOR2_X1 U444 ( .A1(n236), .A2(n243), .ZN(n232) );
  AOI21_X2 U445 ( .B1(n389), .B2(n340), .A(n331), .ZN(n329) );
  INV_X1 U446 ( .A(n223), .ZN(n380) );
  INV_X1 U447 ( .A(n263), .ZN(n261) );
  NAND2_X1 U448 ( .A1(n384), .A2(n274), .ZN(n25) );
  INV_X1 U449 ( .A(n274), .ZN(n272) );
  OAI21_X2 U450 ( .B1(n152), .B2(n144), .A(n145), .ZN(n139) );
  NAND2_X1 U451 ( .A1(n386), .A2(n294), .ZN(n27) );
  OAI21_X2 U452 ( .B1(n286), .B2(n294), .A(n287), .ZN(n285) );
  CLKBUF_X1 U453 ( .A(n82), .Z(n510) );
  NOR2_X2 U454 ( .A1(A[10]), .A2(B[10]), .ZN(n286) );
  INV_X1 U455 ( .A(n167), .ZN(n165) );
  OAI21_X2 U456 ( .B1(n2), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U457 ( .A(n302), .ZN(n300) );
  INV_X1 U458 ( .A(n310), .ZN(n308) );
  NOR2_X2 U459 ( .A1(A[18]), .A2(B[18]), .ZN(n192) );
  INV_X2 U460 ( .A(n332), .ZN(n389) );
  AND2_X2 U461 ( .A1(n347), .A2(n53), .ZN(n499) );
  OR2_X2 U462 ( .A1(A[5]), .A2(B[5]), .ZN(n507) );
  NOR2_X2 U463 ( .A1(n199), .A2(n192), .ZN(n188) );
  NAND2_X1 U464 ( .A1(n391), .A2(n507), .ZN(n335) );
  AOI21_X1 U465 ( .B1(n347), .B2(n507), .A(n340), .ZN(n336) );
  NOR2_X2 U466 ( .A1(n293), .A2(n286), .ZN(n282) );
  INV_X1 U467 ( .A(n79), .ZN(n515) );
  NOR2_X2 U468 ( .A1(A[14]), .A2(B[14]), .ZN(n236) );
  AOI21_X1 U469 ( .B1(n78), .B2(n70), .A(n71), .ZN(n67) );
  NOR2_X1 U470 ( .A1(n499), .A2(n503), .ZN(n52) );
  CLKBUF_X1 U471 ( .A(n266), .Z(n500) );
  XNOR2_X1 U472 ( .A(n65), .B(n7), .ZN(SUM[29]) );
  INV_X1 U473 ( .A(n77), .ZN(n75) );
  NAND2_X1 U474 ( .A1(n77), .A2(n70), .ZN(n66) );
  XNOR2_X1 U475 ( .A(n50), .B(n6), .ZN(SUM[30]) );
  NOR2_X2 U476 ( .A1(A[8]), .A2(B[8]), .ZN(n312) );
  NOR2_X2 U477 ( .A1(A[20]), .A2(B[20]), .ZN(n172) );
  NOR2_X1 U478 ( .A1(A[28]), .A2(B[28]), .ZN(n72) );
  NAND2_X1 U479 ( .A1(A[28]), .A2(B[28]), .ZN(n73) );
  CLKBUF_X1 U480 ( .A(n303), .Z(n501) );
  AOI21_X2 U481 ( .B1(n303), .B2(n260), .A(n261), .ZN(n505) );
  CLKBUF_X1 U482 ( .A(n213), .Z(n502) );
  INV_X1 U483 ( .A(n216), .ZN(n379) );
  CLKBUF_X1 U484 ( .A(n56), .Z(n503) );
  AOI21_X1 U485 ( .B1(n303), .B2(n260), .A(n261), .ZN(n504) );
  AOI21_X1 U486 ( .B1(n56), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X2 U487 ( .B1(n308), .B2(n329), .A(n309), .ZN(n303) );
  OAI21_X2 U488 ( .B1(n82), .B2(n59), .A(n60), .ZN(n56) );
  AOI21_X1 U489 ( .B1(n163), .B2(n374), .A(n154), .ZN(n506) );
  AOI21_X1 U490 ( .B1(n170), .B2(n191), .A(n171), .ZN(n169) );
  OAI21_X1 U491 ( .B1(n192), .B2(n200), .A(n193), .ZN(n191) );
  INV_X1 U492 ( .A(n333), .ZN(n331) );
  NAND2_X1 U493 ( .A1(B[4]), .A2(A[4]), .ZN(n345) );
  NOR2_X4 U494 ( .A1(B[4]), .A2(A[4]), .ZN(n4) );
  NAND2_X1 U495 ( .A1(A[27]), .A2(B[27]), .ZN(n86) );
  NOR2_X1 U496 ( .A1(A[27]), .A2(B[27]), .ZN(n85) );
  NAND2_X1 U497 ( .A1(A[29]), .A2(B[29]), .ZN(n64) );
  NOR2_X1 U498 ( .A1(A[29]), .A2(B[29]), .ZN(n63) );
  OAI21_X1 U499 ( .B1(n172), .B2(n180), .A(n173), .ZN(n171) );
  NAND2_X1 U500 ( .A1(A[24]), .A2(B[24]), .ZN(n121) );
  NAND2_X1 U501 ( .A1(B[1]), .A2(A[1]), .ZN(n361) );
  NOR2_X1 U502 ( .A1(B[1]), .A2(A[1]), .ZN(n360) );
  NOR2_X1 U503 ( .A1(B[0]), .A2(A[0]), .ZN(n362) );
  NAND2_X1 U504 ( .A1(B[0]), .A2(A[0]), .ZN(n363) );
  NOR2_X1 U505 ( .A1(B[2]), .A2(A[2]), .ZN(n356) );
  NAND2_X1 U506 ( .A1(A[30]), .A2(B[30]), .ZN(n49) );
  NOR2_X1 U507 ( .A1(A[30]), .A2(B[30]), .ZN(n48) );
  NAND2_X1 U508 ( .A1(A[22]), .A2(B[22]), .ZN(n145) );
  INV_X1 U509 ( .A(n501), .ZN(n301) );
  NOR2_X1 U510 ( .A1(n319), .A2(n312), .ZN(n310) );
  NOR2_X1 U511 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U512 ( .A1(n520), .A2(n518), .ZN(n79) );
  INV_X2 U513 ( .A(n101), .ZN(n518) );
  CLKBUF_X1 U514 ( .A(n102), .Z(n508) );
  OAI21_X1 U515 ( .B1(n506), .B2(n144), .A(n145), .ZN(n509) );
  NOR2_X1 U516 ( .A1(n4), .A2(n254), .ZN(n248) );
  INV_X1 U517 ( .A(n254), .ZN(n252) );
  NOR2_X2 U518 ( .A1(n164), .A2(n254), .ZN(n160) );
  CLKBUF_X1 U519 ( .A(n93), .Z(n511) );
  INV_X1 U520 ( .A(n500), .ZN(n383) );
  NOR2_X1 U521 ( .A1(n273), .A2(n266), .ZN(n264) );
  OAI21_X1 U522 ( .B1(n266), .B2(n274), .A(n267), .ZN(n265) );
  NOR2_X1 U523 ( .A1(A[12]), .A2(B[12]), .ZN(n266) );
  OAI21_X1 U524 ( .B1(n213), .B2(n168), .A(n169), .ZN(n167) );
  NAND2_X1 U525 ( .A1(B[2]), .A2(A[2]), .ZN(n357) );
  NAND2_X1 U526 ( .A1(A[25]), .A2(B[25]), .ZN(n112) );
  NOR2_X1 U527 ( .A1(A[25]), .A2(B[25]), .ZN(n111) );
  NOR2_X1 U528 ( .A1(A[22]), .A2(B[22]), .ZN(n144) );
  NOR2_X1 U529 ( .A1(A[21]), .A2(B[21]), .ZN(n155) );
  NOR2_X1 U530 ( .A1(n4), .A2(n79), .ZN(n77) );
  NAND2_X1 U531 ( .A1(n302), .A2(n282), .ZN(n280) );
  NAND2_X2 U532 ( .A1(n302), .A2(n260), .ZN(n254) );
  OAI21_X1 U533 ( .B1(n2), .B2(n322), .A(n323), .ZN(n321) );
  OAI21_X1 U534 ( .B1(n2), .B2(n335), .A(n336), .ZN(n334) );
  OAI21_X1 U535 ( .B1(n2), .B2(n4), .A(n345), .ZN(n343) );
  OAI21_X1 U536 ( .B1(n2), .B2(n276), .A(n277), .ZN(n275) );
  OAI21_X1 U537 ( .B1(n2), .B2(n296), .A(n297), .ZN(n295) );
  XOR2_X1 U538 ( .A(n2), .B(n32), .Z(SUM[4]) );
  OAI21_X1 U539 ( .B1(n2), .B2(n315), .A(n316), .ZN(n314) );
  OAI21_X1 U540 ( .B1(n2), .B2(n289), .A(n290), .ZN(n288) );
  OAI21_X1 U541 ( .B1(n2), .B2(n269), .A(n270), .ZN(n268) );
  OAI21_X1 U542 ( .B1(n2), .B2(n75), .A(n76), .ZN(n74) );
  OAI21_X1 U543 ( .B1(n2), .B2(n246), .A(n247), .ZN(n245) );
  OAI21_X1 U544 ( .B1(n2), .B2(n195), .A(n196), .ZN(n194) );
  OAI21_X1 U545 ( .B1(n2), .B2(n88), .A(n89), .ZN(n87) );
  OAI21_X1 U546 ( .B1(n2), .B2(n123), .A(n124), .ZN(n122) );
  OAI21_X1 U547 ( .B1(n2), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X1 U548 ( .B1(n2), .B2(n114), .A(n115), .ZN(n113) );
  OAI21_X1 U549 ( .B1(n2), .B2(n202), .A(n203), .ZN(n201) );
  OAI21_X1 U550 ( .B1(n2), .B2(n97), .A(n98), .ZN(n96) );
  OAI21_X1 U551 ( .B1(n2), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U552 ( .B1(n2), .B2(n219), .A(n220), .ZN(n218) );
  OAI21_X1 U553 ( .B1(n2), .B2(n182), .A(n183), .ZN(n181) );
  OAI21_X1 U554 ( .B1(n2), .B2(n239), .A(n240), .ZN(n238) );
  OAI21_X1 U555 ( .B1(n2), .B2(n226), .A(n227), .ZN(n225) );
  OAI21_X1 U556 ( .B1(n2), .B2(n134), .A(n135), .ZN(n133) );
  OAI21_X1 U557 ( .B1(n2), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U558 ( .B1(n2), .B2(n175), .A(n176), .ZN(n174) );
  NAND2_X1 U559 ( .A1(A[31]), .A2(B[31]), .ZN(n38) );
  NOR2_X1 U560 ( .A1(A[31]), .A2(B[31]), .ZN(n37) );
  NAND2_X1 U561 ( .A1(n388), .A2(n320), .ZN(n29) );
  INV_X1 U562 ( .A(n320), .ZN(n318) );
  INV_X1 U563 ( .A(n506), .ZN(n150) );
  OAI21_X1 U564 ( .B1(n216), .B2(n224), .A(n217), .ZN(n215) );
  INV_X1 U565 ( .A(n192), .ZN(n377) );
  NAND2_X1 U566 ( .A1(n389), .A2(n333), .ZN(n30) );
  NAND2_X2 U567 ( .A1(n507), .A2(n389), .ZN(n326) );
  OAI21_X1 U568 ( .B1(n345), .B2(n326), .A(n329), .ZN(n325) );
  INV_X1 U569 ( .A(n179), .ZN(n376) );
  CLKBUF_X1 U570 ( .A(n163), .Z(n512) );
  NAND2_X1 U571 ( .A1(n513), .A2(n42), .ZN(n514) );
  NAND2_X1 U572 ( .A1(n514), .A2(n41), .ZN(n39) );
  INV_X1 U573 ( .A(n2), .ZN(n513) );
  OAI21_X1 U574 ( .B1(n236), .B2(n244), .A(n237), .ZN(n235) );
  AND2_X1 U575 ( .A1(n46), .A2(n516), .ZN(n517) );
  INV_X1 U576 ( .A(n59), .ZN(n516) );
  AND2_X2 U577 ( .A1(n515), .A2(n516), .ZN(n53) );
  AND2_X2 U578 ( .A1(n83), .A2(n519), .ZN(n520) );
  INV_X1 U579 ( .A(n94), .ZN(n519) );
  AND2_X2 U580 ( .A1(n518), .A2(n519), .ZN(n90) );
  NAND2_X1 U581 ( .A1(n61), .A2(n70), .ZN(n59) );
  OAI21_X1 U582 ( .B1(n345), .B2(n79), .A(n510), .ZN(n78) );
  NAND2_X1 U583 ( .A1(n517), .A2(n515), .ZN(n44) );
  AOI21_X1 U584 ( .B1(n303), .B2(n282), .A(n285), .ZN(n281) );
  OAI21_X1 U585 ( .B1(n345), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X2 U586 ( .B1(n93), .B2(n83), .A(n84), .ZN(n82) );
  OAI21_X1 U587 ( .B1(n107), .B2(n132), .A(n108), .ZN(n106) );
  NOR2_X2 U588 ( .A1(n107), .A2(n131), .ZN(n105) );
  OAI21_X1 U589 ( .B1(n345), .B2(n254), .A(n504), .ZN(n249) );
  INV_X1 U590 ( .A(n505), .ZN(n253) );
  OAI21_X2 U591 ( .B1(n102), .B2(n94), .A(n95), .ZN(n93) );
  OAI21_X2 U592 ( .B1(n505), .B2(n164), .A(n165), .ZN(n163) );
  NOR2_X1 U593 ( .A1(A[26]), .A2(B[26]), .ZN(n94) );
  NAND2_X1 U594 ( .A1(A[26]), .A2(B[26]), .ZN(n95) );
  INV_X1 U595 ( .A(n120), .ZN(n371) );
  NAND2_X1 U596 ( .A1(n370), .A2(n371), .ZN(n107) );
  NAND2_X1 U597 ( .A1(n371), .A2(n121), .ZN(n12) );
  AOI21_X1 U598 ( .B1(n126), .B2(n371), .A(n119), .ZN(n115) );
  NAND2_X1 U599 ( .A1(n125), .A2(n371), .ZN(n114) );
  NOR2_X1 U600 ( .A1(A[24]), .A2(B[24]), .ZN(n120) );
  NOR2_X1 U601 ( .A1(B[3]), .A2(A[3]), .ZN(n353) );
  NAND2_X1 U602 ( .A1(B[3]), .A2(A[3]), .ZN(n354) );
  NAND2_X1 U603 ( .A1(A[23]), .A2(B[23]), .ZN(n132) );
  NOR2_X1 U604 ( .A1(A[23]), .A2(B[23]), .ZN(n131) );
  NAND2_X1 U605 ( .A1(A[21]), .A2(B[21]), .ZN(n156) );
  NAND2_X1 U606 ( .A1(A[6]), .A2(B[6]), .ZN(n333) );
  NAND2_X1 U607 ( .A1(A[7]), .A2(B[7]), .ZN(n320) );
  NOR2_X1 U608 ( .A1(A[7]), .A2(B[7]), .ZN(n319) );
  NAND2_X1 U609 ( .A1(n507), .A2(n342), .ZN(n31) );
  INV_X1 U610 ( .A(n43), .ZN(n41) );
  NOR2_X1 U611 ( .A1(A[19]), .A2(B[19]), .ZN(n179) );
  NAND2_X1 U612 ( .A1(A[19]), .A2(B[19]), .ZN(n180) );
  NAND2_X1 U613 ( .A1(A[18]), .A2(B[18]), .ZN(n193) );
  NAND2_X1 U614 ( .A1(A[16]), .A2(B[16]), .ZN(n217) );
  NOR2_X1 U615 ( .A1(A[13]), .A2(B[13]), .ZN(n243) );
  NAND2_X1 U616 ( .A1(A[13]), .A2(B[13]), .ZN(n244) );
  NOR2_X1 U617 ( .A1(A[17]), .A2(B[17]), .ZN(n199) );
  NAND2_X1 U618 ( .A1(A[17]), .A2(B[17]), .ZN(n200) );
  AOI21_X2 U619 ( .B1(n139), .B2(n105), .A(n106), .ZN(n102) );
  INV_X1 U620 ( .A(n508), .ZN(n100) );
  AOI21_X1 U621 ( .B1(n509), .B2(n372), .A(n130), .ZN(n128) );
  NOR2_X1 U622 ( .A1(A[15]), .A2(B[15]), .ZN(n223) );
  NAND2_X1 U623 ( .A1(A[15]), .A2(B[15]), .ZN(n224) );
  INV_X1 U624 ( .A(n236), .ZN(n381) );
  NAND2_X1 U625 ( .A1(n391), .A2(n53), .ZN(n51) );
  NAND2_X1 U626 ( .A1(A[14]), .A2(B[14]), .ZN(n237) );
  AOI21_X1 U627 ( .B1(n214), .B2(n235), .A(n215), .ZN(n213) );
  NAND2_X1 U628 ( .A1(n232), .A2(n214), .ZN(n210) );
  INV_X1 U629 ( .A(n172), .ZN(n375) );
  NAND2_X1 U630 ( .A1(A[20]), .A2(B[20]), .ZN(n173) );
  NAND2_X1 U631 ( .A1(A[12]), .A2(B[12]), .ZN(n267) );
  NOR2_X1 U632 ( .A1(n254), .A2(n210), .ZN(n208) );
  OAI21_X1 U633 ( .B1(n504), .B2(n210), .A(n502), .ZN(n209) );
  NOR2_X2 U634 ( .A1(n168), .A2(n210), .ZN(n166) );
  NAND2_X1 U635 ( .A1(n208), .A2(n188), .ZN(n186) );
  AOI21_X1 U636 ( .B1(n209), .B2(n188), .A(n191), .ZN(n187) );
  NAND2_X2 U637 ( .A1(n188), .A2(n170), .ZN(n168) );
  NOR2_X1 U638 ( .A1(A[9]), .A2(B[9]), .ZN(n293) );
  NAND2_X1 U639 ( .A1(A[9]), .A2(B[9]), .ZN(n294) );
  NAND2_X1 U640 ( .A1(n282), .A2(n264), .ZN(n262) );
  AOI21_X1 U641 ( .B1(n285), .B2(n264), .A(n265), .ZN(n263) );
  NOR2_X1 U642 ( .A1(A[11]), .A2(B[11]), .ZN(n273) );
  NAND2_X1 U643 ( .A1(A[11]), .A2(B[11]), .ZN(n274) );
  NAND2_X1 U644 ( .A1(n252), .A2(n498), .ZN(n230) );
  AOI21_X1 U645 ( .B1(n253), .B2(n498), .A(n235), .ZN(n231) );
  NOR2_X1 U646 ( .A1(A[6]), .A2(B[6]), .ZN(n332) );
  NAND2_X1 U647 ( .A1(A[5]), .A2(B[5]), .ZN(n342) );
  NAND2_X1 U648 ( .A1(n391), .A2(n160), .ZN(n158) );
  AOI21_X1 U649 ( .B1(n347), .B2(n160), .A(n512), .ZN(n159) );
  NAND2_X2 U650 ( .A1(n160), .A2(n374), .ZN(n151) );
  NAND2_X1 U651 ( .A1(A[8]), .A2(B[8]), .ZN(n313) );
  INV_X1 U652 ( .A(n312), .ZN(n387) );
  NAND2_X1 U653 ( .A1(n391), .A2(n90), .ZN(n88) );
  AOI21_X1 U654 ( .B1(n347), .B2(n90), .A(n511), .ZN(n89) );
  OAI21_X1 U655 ( .B1(n312), .B2(n320), .A(n313), .ZN(n311) );
  INV_X1 U656 ( .A(n286), .ZN(n385) );
  XNOR2_X1 U657 ( .A(n39), .B(n5), .ZN(SUM[31]) );
  NAND2_X1 U658 ( .A1(A[10]), .A2(B[10]), .ZN(n287) );
  NAND2_X1 U659 ( .A1(n391), .A2(n138), .ZN(n134) );
  AOI21_X1 U660 ( .B1(n347), .B2(n138), .A(n509), .ZN(n135) );
  NAND2_X1 U661 ( .A1(n138), .A2(n372), .ZN(n127) );
  NAND2_X2 U662 ( .A1(n138), .A2(n105), .ZN(n101) );
  INV_X2 U663 ( .A(n101), .ZN(n99) );
  INV_X2 U664 ( .A(n86), .ZN(n84) );
  INV_X2 U665 ( .A(n78), .ZN(n76) );
  INV_X2 U666 ( .A(n73), .ZN(n71) );
  INV_X2 U667 ( .A(n64), .ZN(n62) );
  INV_X2 U668 ( .A(n49), .ZN(n47) );
  INV_X2 U669 ( .A(n362), .ZN(n395) );
  INV_X2 U670 ( .A(n360), .ZN(n394) );
  INV_X2 U671 ( .A(n356), .ZN(n393) );
  INV_X2 U672 ( .A(n353), .ZN(n392) );
  INV_X2 U673 ( .A(n144), .ZN(n373) );
  INV_X2 U674 ( .A(n94), .ZN(n369) );
  INV_X2 U675 ( .A(n85), .ZN(n83) );
  INV_X2 U676 ( .A(n72), .ZN(n70) );
  INV_X2 U677 ( .A(n63), .ZN(n61) );
  INV_X2 U678 ( .A(n48), .ZN(n46) );
  INV_X2 U679 ( .A(n37), .ZN(n364) );
  INV_X2 U680 ( .A(n359), .ZN(n358) );
  INV_X2 U681 ( .A(n4), .ZN(n391) );
  INV_X2 U682 ( .A(n342), .ZN(n340) );
  INV_X2 U683 ( .A(n325), .ZN(n323) );
  INV_X2 U684 ( .A(n324), .ZN(n322) );
  INV_X2 U685 ( .A(n319), .ZN(n388) );
  INV_X2 U686 ( .A(n311), .ZN(n309) );
  INV_X2 U687 ( .A(n299), .ZN(n297) );
  INV_X2 U688 ( .A(n298), .ZN(n296) );
  INV_X2 U689 ( .A(n294), .ZN(n292) );
  INV_X2 U690 ( .A(n293), .ZN(n386) );
  INV_X2 U691 ( .A(n279), .ZN(n277) );
  INV_X2 U692 ( .A(n278), .ZN(n276) );
  INV_X2 U693 ( .A(n273), .ZN(n384) );
  INV_X2 U694 ( .A(n262), .ZN(n260) );
  INV_X2 U695 ( .A(n249), .ZN(n247) );
  INV_X2 U696 ( .A(n248), .ZN(n246) );
  INV_X2 U697 ( .A(n244), .ZN(n242) );
  INV_X2 U698 ( .A(n243), .ZN(n382) );
  INV_X2 U699 ( .A(n229), .ZN(n227) );
  INV_X2 U700 ( .A(n228), .ZN(n226) );
  INV_X2 U701 ( .A(n224), .ZN(n222) );
  INV_X2 U702 ( .A(n209), .ZN(n207) );
  INV_X2 U703 ( .A(n208), .ZN(n206) );
  INV_X2 U704 ( .A(n205), .ZN(n203) );
  INV_X2 U705 ( .A(n204), .ZN(n202) );
  INV_X2 U706 ( .A(n200), .ZN(n198) );
  INV_X2 U707 ( .A(n199), .ZN(n378) );
  INV_X2 U708 ( .A(n185), .ZN(n183) );
  INV_X2 U709 ( .A(n184), .ZN(n182) );
  INV_X2 U710 ( .A(n180), .ZN(n178) );
  INV_X2 U711 ( .A(n166), .ZN(n164) );
  INV_X2 U712 ( .A(n156), .ZN(n154) );
  INV_X2 U713 ( .A(n155), .ZN(n374) );
  INV_X2 U714 ( .A(n151), .ZN(n149) );
  INV_X2 U715 ( .A(n132), .ZN(n130) );
  INV_X2 U716 ( .A(n131), .ZN(n372) );
  INV_X2 U717 ( .A(n126), .ZN(n124) );
  INV_X2 U718 ( .A(n125), .ZN(n123) );
  INV_X2 U719 ( .A(n121), .ZN(n119) );
  INV_X2 U720 ( .A(n112), .ZN(n110) );
  INV_X2 U721 ( .A(n111), .ZN(n370) );
  INV_X2 U722 ( .A(n36), .ZN(SUM[0]) );
endmodule


module Xi_core_DW01_sub_1 ( A, B, DIFF, CI, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n123, n124, n126, n127,
         n128, n129, n130, n131, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n146, n148, n149, n150, n151, n152, n153, n154, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n176, n177, n178, n179, n180,
         n181, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n200, n201, n202, n203, n204, n205, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n228, n229, n230, n231, n232,
         n233, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n252, n253, n254, n255, n256, n257, n261,
         n262, n263, n264, n265, n266, n267, n268, n271, n272, n273, n274,
         n277, n278, n279, n280, n281, n282, n284, n285, n286, n287, n288,
         n289, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n308, n309, n310, n311, n312, n313, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n332, n334, n336, n337, n338, n339, n340, n341, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n363, n364, n365, n366, n368, n370, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n388, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  NAND2_X4 U6 ( .A1(n386), .A2(n37), .ZN(n5) );
  NAND2_X4 U20 ( .A1(n45), .A2(n48), .ZN(n6) );
  XNOR2_X2 U24 ( .A(n58), .B(n7), .ZN(DIFF[29]) );
  NAND2_X4 U32 ( .A1(n388), .A2(n57), .ZN(n7) );
  XNOR2_X2 U36 ( .A(n75), .B(n8), .ZN(DIFF[28]) );
  NAND2_X4 U38 ( .A1(n413), .A2(n61), .ZN(n59) );
  AOI21_X4 U39 ( .B1(n370), .B2(n61), .A(n62), .ZN(n60) );
  NOR2_X4 U46 ( .A1(n69), .A2(n93), .ZN(n67) );
  OAI21_X4 U47 ( .B1(n94), .B2(n69), .A(n70), .ZN(n68) );
  NAND2_X4 U48 ( .A1(n80), .A2(n71), .ZN(n69) );
  AOI21_X4 U49 ( .B1(n71), .B2(n81), .A(n72), .ZN(n70) );
  NAND2_X4 U52 ( .A1(n71), .A2(n74), .ZN(n8) );
  XNOR2_X2 U56 ( .A(n84), .B(n9), .ZN(DIFF[27]) );
  NAND2_X4 U58 ( .A1(n87), .A2(n80), .ZN(n76) );
  AOI21_X4 U59 ( .B1(n88), .B2(n80), .A(n81), .ZN(n77) );
  NAND2_X4 U64 ( .A1(n80), .A2(n83), .ZN(n9) );
  NOR2_X4 U72 ( .A1(n4), .A2(n89), .ZN(n87) );
  OAI21_X4 U73 ( .B1(n368), .B2(n89), .A(n90), .ZN(n88) );
  NAND2_X4 U78 ( .A1(n392), .A2(n95), .ZN(n93) );
  AOI21_X4 U79 ( .B1(n95), .B2(n105), .A(n96), .ZN(n94) );
  NAND2_X4 U82 ( .A1(n95), .A2(n98), .ZN(n10) );
  XNOR2_X2 U86 ( .A(n108), .B(n11), .ZN(DIFF[25]) );
  NAND2_X4 U88 ( .A1(n111), .A2(n392), .ZN(n100) );
  AOI21_X4 U89 ( .B1(n112), .B2(n392), .A(n105), .ZN(n101) );
  NAND2_X4 U94 ( .A1(n392), .A2(n107), .ZN(n11) );
  XNOR2_X2 U98 ( .A(n129), .B(n12), .ZN(DIFF[24]) );
  NOR2_X4 U102 ( .A1(n4), .A2(n113), .ZN(n111) );
  OAI21_X4 U103 ( .B1(n368), .B2(n113), .A(n114), .ZN(n112) );
  NAND2_X4 U114 ( .A1(n394), .A2(n393), .ZN(n123) );
  AOI21_X4 U115 ( .B1(n135), .B2(n393), .A(n126), .ZN(n124) );
  NAND2_X4 U118 ( .A1(n393), .A2(n128), .ZN(n12) );
  XNOR2_X2 U122 ( .A(n138), .B(n13), .ZN(DIFF[23]) );
  NAND2_X4 U130 ( .A1(n394), .A2(n137), .ZN(n13) );
  XNOR2_X2 U134 ( .A(n151), .B(n14), .ZN(DIFF[22]) );
  NAND2_X4 U146 ( .A1(n395), .A2(n150), .ZN(n14) );
  XNOR2_X2 U150 ( .A(n160), .B(n15), .ZN(DIFF[21]) );
  NOR2_X4 U156 ( .A1(n165), .A2(n158), .ZN(n154) );
  NAND2_X4 U158 ( .A1(n396), .A2(n159), .ZN(n15) );
  NAND2_X4 U164 ( .A1(n413), .A2(n163), .ZN(n161) );
  AOI21_X4 U165 ( .B1(n370), .B2(n163), .A(n164), .ZN(n162) );
  NOR2_X4 U174 ( .A1(n197), .A2(n173), .ZN(n171) );
  XNOR2_X2 U184 ( .A(n188), .B(n17), .ZN(DIFF[19]) );
  XNOR2_X2 U196 ( .A(n203), .B(n18), .ZN(DIFF[18]) );
  NOR2_X4 U200 ( .A1(n4), .A2(n193), .ZN(n191) );
  OAI21_X4 U201 ( .B1(n368), .B2(n193), .A(n194), .ZN(n192) );
  NAND2_X4 U202 ( .A1(n219), .A2(n195), .ZN(n193) );
  AOI21_X4 U203 ( .B1(n220), .B2(n195), .A(n196), .ZN(n194) );
  XNOR2_X2 U214 ( .A(n212), .B(n19), .ZN(DIFF[17]) );
  XNOR2_X2 U226 ( .A(n231), .B(n20), .ZN(DIFF[16]) );
  NOR2_X4 U230 ( .A1(n4), .A2(n217), .ZN(n215) );
  OAI21_X4 U231 ( .B1(n368), .B2(n217), .A(n218), .ZN(n216) );
  NOR2_X4 U234 ( .A1(n273), .A2(n221), .ZN(n219) );
  OAI21_X4 U235 ( .B1(n274), .B2(n221), .A(n222), .ZN(n220) );
  XNOR2_X2 U248 ( .A(n240), .B(n21), .ZN(DIFF[15]) );
  XNOR2_X2 U260 ( .A(n255), .B(n22), .ZN(DIFF[14]) );
  NOR2_X4 U264 ( .A1(n4), .A2(n245), .ZN(n243) );
  OAI21_X4 U265 ( .B1(n368), .B2(n245), .A(n246), .ZN(n244) );
  XNOR2_X2 U278 ( .A(n264), .B(n23), .ZN(DIFF[13]) );
  NOR2_X4 U294 ( .A1(n4), .A2(n273), .ZN(n267) );
  OAI21_X4 U295 ( .B1(n368), .B2(n273), .A(n274), .ZN(n268) );
  XNOR2_X2 U316 ( .A(n296), .B(n25), .ZN(DIFF[11]) );
  XNOR2_X2 U328 ( .A(n311), .B(n26), .ZN(DIFF[10]) );
  NOR2_X4 U332 ( .A1(n4), .A2(n301), .ZN(n299) );
  OAI21_X4 U333 ( .B1(n368), .B2(n301), .A(n302), .ZN(n300) );
  NAND2_X4 U334 ( .A1(n327), .A2(n303), .ZN(n301) );
  AOI21_X4 U335 ( .B1(n328), .B2(n303), .A(n304), .ZN(n302) );
  XNOR2_X2 U346 ( .A(n320), .B(n27), .ZN(DIFF[9]) );
  XNOR2_X2 U358 ( .A(n339), .B(n28), .ZN(DIFF[8]) );
  NAND2_X4 U376 ( .A1(n409), .A2(n338), .ZN(n28) );
  XNOR2_X2 U380 ( .A(n348), .B(n29), .ZN(DIFF[7]) );
  XNOR2_X2 U392 ( .A(n359), .B(n30), .ZN(DIFF[6]) );
  NOR2_X4 U396 ( .A1(n4), .A2(n353), .ZN(n351) );
  OAI21_X4 U397 ( .B1(n368), .B2(n353), .A(n354), .ZN(n352) );
  NAND2_X4 U402 ( .A1(n411), .A2(n358), .ZN(n30) );
  XNOR2_X2 U406 ( .A(n366), .B(n31), .ZN(DIFF[5]) );
  NAND2_X4 U408 ( .A1(n413), .A2(n412), .ZN(n360) );
  AOI21_X4 U409 ( .B1(n370), .B2(n412), .A(n363), .ZN(n361) );
  NAND2_X4 U422 ( .A1(n413), .A2(n368), .ZN(n32) );
  XNOR2_X2 U426 ( .A(n378), .B(n33), .ZN(DIFF[3]) );
  AOI21_X4 U427 ( .B1(n374), .B2(n382), .A(n375), .ZN(n2) );
  NOR2_X4 U428 ( .A1(n379), .A2(n376), .ZN(n374) );
  NAND2_X4 U430 ( .A1(n414), .A2(n377), .ZN(n33) );
  XOR2_X2 U434 ( .A(n34), .B(n381), .Z(DIFF[2]) );
  OAI21_X4 U435 ( .B1(n381), .B2(n379), .A(n380), .ZN(n378) );
  NAND2_X4 U436 ( .A1(n415), .A2(n380), .ZN(n34) );
  XOR2_X2 U440 ( .A(n35), .B(n385), .Z(DIFF[1]) );
  NAND2_X4 U443 ( .A1(n416), .A2(n384), .ZN(n35) );
  XNOR2_X1 U484 ( .A(n179), .B(n16), .ZN(DIFF[20]) );
  INV_X2 U485 ( .A(n564), .ZN(n274) );
  OR2_X1 U486 ( .A1(n368), .A2(n43), .ZN(n551) );
  NAND2_X1 U487 ( .A1(n551), .A2(n44), .ZN(n42) );
  OAI21_X2 U488 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U489 ( .A(n112), .ZN(n110) );
  CLKBUF_X1 U490 ( .A(n116), .Z(n571) );
  AOI21_X1 U491 ( .B1(n142), .B2(n394), .A(n135), .ZN(n131) );
  INV_X1 U492 ( .A(n142), .ZN(n140) );
  OR2_X1 U493 ( .A1(n2), .A2(n50), .ZN(n552) );
  NAND2_X1 U494 ( .A1(n552), .A2(n51), .ZN(n49) );
  AOI21_X1 U495 ( .B1(n370), .B2(n52), .A(n565), .ZN(n51) );
  AOI21_X2 U496 ( .B1(n224), .B2(n171), .A(n172), .ZN(n170) );
  AOI21_X2 U497 ( .B1(n116), .B2(n67), .A(n68), .ZN(n64) );
  AOI21_X1 U498 ( .B1(n272), .B2(n167), .A(n168), .ZN(n166) );
  OAI21_X1 U499 ( .B1(n146), .B2(n123), .A(n124), .ZN(n116) );
  XNOR2_X1 U500 ( .A(n99), .B(n10), .ZN(DIFF[26]) );
  CLKBUF_X1 U501 ( .A(n55), .Z(n565) );
  INV_X1 U502 ( .A(n211), .ZN(n209) );
  NAND2_X1 U503 ( .A1(n141), .A2(n394), .ZN(n130) );
  INV_X1 U504 ( .A(n141), .ZN(n139) );
  NOR2_X1 U505 ( .A1(A[18]), .A2(n430), .ZN(n201) );
  OAI21_X1 U506 ( .B1(n383), .B2(n385), .A(n384), .ZN(n382) );
  OAI21_X1 U507 ( .B1(n380), .B2(n376), .A(n377), .ZN(n375) );
  INV_X1 U508 ( .A(n285), .ZN(n405) );
  AOI21_X2 U509 ( .B1(n405), .B2(n293), .A(n284), .ZN(n282) );
  AOI21_X2 U510 ( .B1(n403), .B2(n261), .A(n252), .ZN(n250) );
  AOI21_X1 U511 ( .B1(n403), .B2(n558), .A(n252), .ZN(n561) );
  NOR2_X1 U512 ( .A1(n143), .A2(n123), .ZN(n554) );
  NOR2_X1 U513 ( .A1(n143), .A2(n123), .ZN(n553) );
  NOR2_X1 U514 ( .A1(n165), .A2(n158), .ZN(n555) );
  AND2_X1 U515 ( .A1(n555), .A2(n556), .ZN(n115) );
  AND2_X1 U516 ( .A1(n557), .A2(n395), .ZN(n556) );
  INV_X1 U517 ( .A(n123), .ZN(n557) );
  XNOR2_X1 U518 ( .A(n49), .B(n6), .ZN(DIFF[30]) );
  INV_X1 U519 ( .A(n357), .ZN(n411) );
  AOI21_X1 U520 ( .B1(n55), .B2(n45), .A(n46), .ZN(n44) );
  NOR2_X2 U521 ( .A1(n364), .A2(n357), .ZN(n355) );
  XNOR2_X1 U522 ( .A(n287), .B(n24), .ZN(DIFF[12]) );
  NOR2_X1 U523 ( .A1(A[28]), .A2(n420), .ZN(n73) );
  NAND2_X1 U524 ( .A1(A[28]), .A2(n420), .ZN(n74) );
  NOR2_X2 U525 ( .A1(A[6]), .A2(n442), .ZN(n357) );
  NAND2_X4 U526 ( .A1(n574), .A2(A[4]), .ZN(n368) );
  NOR2_X4 U527 ( .A1(n574), .A2(A[4]), .ZN(n4) );
  NAND2_X2 U528 ( .A1(A[27]), .A2(n421), .ZN(n83) );
  NAND2_X1 U529 ( .A1(A[29]), .A2(n419), .ZN(n57) );
  NOR2_X1 U530 ( .A1(A[29]), .A2(n419), .ZN(n56) );
  NOR2_X1 U531 ( .A1(A[24]), .A2(n424), .ZN(n127) );
  NAND2_X1 U532 ( .A1(A[24]), .A2(n424), .ZN(n128) );
  NAND2_X1 U533 ( .A1(n402), .A2(n401), .ZN(n225) );
  NAND2_X1 U534 ( .A1(n403), .A2(n254), .ZN(n22) );
  NAND2_X2 U535 ( .A1(n404), .A2(n403), .ZN(n249) );
  NAND2_X1 U536 ( .A1(n577), .A2(A[1]), .ZN(n384) );
  NOR2_X1 U537 ( .A1(n577), .A2(A[1]), .ZN(n383) );
  XNOR2_X1 U538 ( .A(n578), .B(A[0]), .ZN(DIFF[0]) );
  NAND2_X1 U539 ( .A1(A[25]), .A2(n423), .ZN(n107) );
  NOR2_X4 U540 ( .A1(n576), .A2(A[2]), .ZN(n379) );
  NAND2_X1 U541 ( .A1(A[30]), .A2(n418), .ZN(n48) );
  NOR2_X1 U542 ( .A1(A[30]), .A2(n418), .ZN(n47) );
  OAI21_X1 U543 ( .B1(n326), .B2(n277), .A(n278), .ZN(n272) );
  AOI21_X1 U544 ( .B1(n409), .B2(n345), .A(n336), .ZN(n334) );
  INV_X1 U545 ( .A(n347), .ZN(n345) );
  CLKBUF_X1 U546 ( .A(n261), .Z(n558) );
  INV_X1 U547 ( .A(n328), .ZN(n559) );
  NOR2_X4 U548 ( .A1(n63), .A2(n56), .ZN(n52) );
  NOR2_X2 U549 ( .A1(n249), .A2(n225), .ZN(n223) );
  NAND2_X1 U550 ( .A1(A[15]), .A2(n433), .ZN(n239) );
  INV_X2 U551 ( .A(B[6]), .ZN(n442) );
  NAND2_X1 U552 ( .A1(n405), .A2(n286), .ZN(n24) );
  CLKBUF_X1 U553 ( .A(n168), .Z(n560) );
  NAND2_X1 U554 ( .A1(n407), .A2(n310), .ZN(n26) );
  AOI21_X2 U555 ( .B1(n407), .B2(n317), .A(n308), .ZN(n306) );
  INV_X1 U556 ( .A(n309), .ZN(n407) );
  INV_X1 U557 ( .A(n346), .ZN(n410) );
  AND2_X2 U558 ( .A1(n410), .A2(n409), .ZN(n569) );
  INV_X1 U559 ( .A(n254), .ZN(n252) );
  NAND2_X1 U560 ( .A1(n412), .A2(n365), .ZN(n31) );
  INV_X1 U561 ( .A(n365), .ZN(n363) );
  INV_X1 U562 ( .A(n356), .ZN(n354) );
  INV_X1 U563 ( .A(n63), .ZN(n61) );
  NAND2_X1 U564 ( .A1(n171), .A2(n223), .ZN(n169) );
  INV_X1 U565 ( .A(n223), .ZN(n221) );
  NAND2_X1 U566 ( .A1(n356), .A2(n569), .ZN(n562) );
  INV_X1 U567 ( .A(n332), .ZN(n563) );
  AND2_X2 U568 ( .A1(n562), .A2(n563), .ZN(n326) );
  OAI21_X2 U569 ( .B1(n357), .B2(n365), .A(n358), .ZN(n356) );
  INV_X1 U570 ( .A(n334), .ZN(n332) );
  NAND2_X2 U571 ( .A1(n115), .A2(n67), .ZN(n63) );
  NAND2_X1 U572 ( .A1(A[7]), .A2(n441), .ZN(n347) );
  AOI21_X2 U573 ( .B1(n397), .B2(n185), .A(n176), .ZN(n174) );
  INV_X1 U574 ( .A(n229), .ZN(n401) );
  AOI21_X2 U575 ( .B1(n401), .B2(n237), .A(n228), .ZN(n226) );
  NAND2_X1 U576 ( .A1(n401), .A2(n230), .ZN(n20) );
  NAND2_X1 U577 ( .A1(n267), .A2(n404), .ZN(n256) );
  INV_X1 U578 ( .A(B[17]), .ZN(n431) );
  OAI21_X1 U579 ( .B1(n326), .B2(n277), .A(n278), .ZN(n564) );
  NOR2_X1 U580 ( .A1(n578), .A2(A[0]), .ZN(n385) );
  NAND2_X1 U581 ( .A1(n576), .A2(A[2]), .ZN(n380) );
  NOR2_X1 U582 ( .A1(A[25]), .A2(n423), .ZN(n106) );
  NOR2_X1 U583 ( .A1(A[22]), .A2(n426), .ZN(n149) );
  NAND2_X1 U584 ( .A1(A[22]), .A2(n426), .ZN(n150) );
  NOR2_X1 U585 ( .A1(A[27]), .A2(n421), .ZN(n82) );
  NAND2_X1 U586 ( .A1(A[21]), .A2(n427), .ZN(n159) );
  NOR2_X1 U587 ( .A1(A[21]), .A2(n427), .ZN(n158) );
  NAND2_X1 U588 ( .A1(n410), .A2(n347), .ZN(n29) );
  NAND2_X1 U589 ( .A1(n351), .A2(n410), .ZN(n340) );
  AOI21_X1 U590 ( .B1(n352), .B2(n410), .A(n345), .ZN(n341) );
  NAND2_X1 U591 ( .A1(A[31]), .A2(n417), .ZN(n37) );
  NOR2_X1 U592 ( .A1(A[31]), .A2(n417), .ZN(n36) );
  NAND2_X1 U593 ( .A1(n215), .A2(n400), .ZN(n204) );
  AOI21_X1 U594 ( .B1(n216), .B2(n400), .A(n209), .ZN(n205) );
  NAND2_X1 U595 ( .A1(n400), .A2(n211), .ZN(n19) );
  NAND2_X2 U596 ( .A1(n400), .A2(n399), .ZN(n197) );
  NAND2_X1 U597 ( .A1(A[17]), .A2(n431), .ZN(n211) );
  NOR2_X2 U598 ( .A1(n305), .A2(n281), .ZN(n279) );
  OAI21_X1 U599 ( .B1(n306), .B2(n281), .A(n282), .ZN(n280) );
  INV_X1 U600 ( .A(n279), .ZN(n277) );
  NAND2_X1 U601 ( .A1(n406), .A2(n405), .ZN(n281) );
  AOI21_X1 U602 ( .B1(n564), .B2(n167), .A(n560), .ZN(n566) );
  OAI21_X1 U603 ( .B1(n250), .B2(n225), .A(n226), .ZN(n224) );
  CLKBUF_X1 U604 ( .A(n146), .Z(n567) );
  CLKBUF_X1 U605 ( .A(n157), .Z(n568) );
  NAND2_X1 U606 ( .A1(n299), .A2(n406), .ZN(n288) );
  AOI21_X1 U607 ( .B1(n300), .B2(n406), .A(n293), .ZN(n289) );
  NAND2_X1 U608 ( .A1(n406), .A2(n295), .ZN(n25) );
  OAI21_X1 U609 ( .B1(n166), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U610 ( .A1(n4), .A2(n325), .ZN(n323) );
  INV_X1 U611 ( .A(n325), .ZN(n327) );
  NOR2_X2 U612 ( .A1(n277), .A2(n325), .ZN(n271) );
  INV_X1 U613 ( .A(n170), .ZN(n168) );
  NAND2_X1 U614 ( .A1(n399), .A2(n202), .ZN(n18) );
  INV_X1 U615 ( .A(n202), .ZN(n200) );
  NAND2_X1 U616 ( .A1(n397), .A2(n178), .ZN(n16) );
  INV_X1 U617 ( .A(n178), .ZN(n176) );
  INV_X1 U618 ( .A(n201), .ZN(n399) );
  INV_X1 U619 ( .A(n224), .ZN(n222) );
  AOI21_X2 U620 ( .B1(n399), .B2(n209), .A(n200), .ZN(n198) );
  NAND2_X2 U621 ( .A1(n355), .A2(n569), .ZN(n325) );
  AOI21_X2 U622 ( .B1(n157), .B2(n395), .A(n148), .ZN(n146) );
  NAND2_X1 U623 ( .A1(A[19]), .A2(n429), .ZN(n187) );
  INV_X1 U624 ( .A(n561), .ZN(n248) );
  INV_X1 U625 ( .A(n198), .ZN(n196) );
  OAI21_X1 U626 ( .B1(n198), .B2(n173), .A(n174), .ZN(n172) );
  CLKBUF_X1 U627 ( .A(n64), .Z(n570) );
  NAND2_X1 U628 ( .A1(A[14]), .A2(n434), .ZN(n254) );
  NOR2_X1 U629 ( .A1(A[14]), .A2(n434), .ZN(n253) );
  AOI21_X1 U630 ( .B1(n268), .B2(n404), .A(n558), .ZN(n257) );
  INV_X1 U631 ( .A(B[13]), .ZN(n435) );
  INV_X1 U632 ( .A(B[9]), .ZN(n439) );
  INV_X1 U633 ( .A(B[7]), .ZN(n441) );
  NAND2_X1 U634 ( .A1(n402), .A2(n239), .ZN(n21) );
  NAND2_X1 U635 ( .A1(n243), .A2(n402), .ZN(n232) );
  AOI21_X1 U636 ( .B1(n244), .B2(n402), .A(n237), .ZN(n233) );
  INV_X1 U637 ( .A(B[15]), .ZN(n433) );
  NAND2_X1 U638 ( .A1(n271), .A2(n247), .ZN(n245) );
  INV_X1 U639 ( .A(n271), .ZN(n273) );
  NAND2_X1 U640 ( .A1(A[20]), .A2(n428), .ZN(n178) );
  NAND2_X1 U641 ( .A1(A[18]), .A2(n430), .ZN(n202) );
  NAND2_X1 U642 ( .A1(n52), .A2(n45), .ZN(n43) );
  INV_X1 U643 ( .A(n566), .ZN(n164) );
  AOI21_X1 U644 ( .B1(n564), .B2(n247), .A(n248), .ZN(n246) );
  INV_X1 U645 ( .A(B[11]), .ZN(n437) );
  NOR2_X1 U646 ( .A1(n43), .A2(n4), .ZN(n41) );
  NAND2_X1 U647 ( .A1(n408), .A2(n319), .ZN(n27) );
  AOI21_X1 U648 ( .B1(n324), .B2(n408), .A(n317), .ZN(n313) );
  NAND2_X1 U649 ( .A1(n323), .A2(n408), .ZN(n312) );
  NAND2_X2 U650 ( .A1(n408), .A2(n407), .ZN(n305) );
  NAND2_X2 U651 ( .A1(n154), .A2(n395), .ZN(n143) );
  INV_X1 U652 ( .A(B[5]), .ZN(n443) );
  OAI21_X1 U653 ( .B1(n2), .B2(n340), .A(n341), .ZN(n339) );
  OAI21_X1 U654 ( .B1(n2), .B2(n288), .A(n289), .ZN(n287) );
  OAI21_X1 U655 ( .B1(n2), .B2(n360), .A(n361), .ZN(n359) );
  OAI21_X1 U656 ( .B1(n2), .B2(n349), .A(n350), .ZN(n348) );
  OAI21_X1 U657 ( .B1(n2), .B2(n213), .A(n214), .ZN(n212) );
  OAI21_X1 U658 ( .B1(n2), .B2(n204), .A(n205), .ZN(n203) );
  OAI21_X1 U659 ( .B1(n2), .B2(n297), .A(n298), .ZN(n296) );
  OAI21_X1 U660 ( .B1(n2), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U661 ( .B1(n2), .B2(n321), .A(n322), .ZN(n320) );
  OAI21_X1 U662 ( .B1(n2), .B2(n312), .A(n313), .ZN(n311) );
  OAI21_X1 U663 ( .B1(n2), .B2(n241), .A(n242), .ZN(n240) );
  OAI21_X1 U664 ( .B1(n2), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U665 ( .B1(n2), .B2(n161), .A(n162), .ZN(n160) );
  OAI21_X1 U666 ( .B1(n2), .B2(n85), .A(n86), .ZN(n84) );
  OAI21_X1 U667 ( .B1(n2), .B2(n180), .A(n181), .ZN(n179) );
  OAI21_X1 U668 ( .B1(n2), .B2(n189), .A(n190), .ZN(n188) );
  OAI21_X1 U669 ( .B1(n2), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X1 U670 ( .B1(n2), .B2(n139), .A(n140), .ZN(n138) );
  OAI21_X1 U671 ( .B1(n2), .B2(n232), .A(n233), .ZN(n231) );
  OAI21_X1 U672 ( .B1(n2), .B2(n256), .A(n257), .ZN(n255) );
  OAI21_X1 U673 ( .B1(n2), .B2(n76), .A(n77), .ZN(n75) );
  XOR2_X1 U674 ( .A(n2), .B(n32), .Z(DIFF[4]) );
  OAI21_X1 U675 ( .B1(n2), .B2(n4), .A(n368), .ZN(n366) );
  OAI21_X1 U676 ( .B1(n2), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U677 ( .B1(n2), .B2(n59), .A(n60), .ZN(n58) );
  INV_X4 U678 ( .A(n2), .ZN(n572) );
  INV_X1 U679 ( .A(n326), .ZN(n328) );
  OAI21_X1 U680 ( .B1(n368), .B2(n325), .A(n559), .ZN(n324) );
  AOI21_X1 U681 ( .B1(n571), .B2(n91), .A(n92), .ZN(n90) );
  OAI21_X1 U682 ( .B1(n64), .B2(n56), .A(n57), .ZN(n55) );
  INV_X1 U683 ( .A(B[19]), .ZN(n429) );
  INV_X1 U684 ( .A(B[10]), .ZN(n438) );
  INV_X1 U685 ( .A(B[12]), .ZN(n436) );
  NAND2_X1 U686 ( .A1(n572), .A2(n41), .ZN(n573) );
  NAND2_X1 U687 ( .A1(n40), .A2(n573), .ZN(n38) );
  INV_X1 U688 ( .A(B[14]), .ZN(n434) );
  INV_X1 U689 ( .A(B[20]), .ZN(n428) );
  NOR2_X1 U690 ( .A1(A[26]), .A2(n422), .ZN(n97) );
  NAND2_X1 U691 ( .A1(A[26]), .A2(n422), .ZN(n98) );
  INV_X1 U692 ( .A(B[18]), .ZN(n430) );
  NOR2_X2 U693 ( .A1(n575), .A2(A[3]), .ZN(n376) );
  NAND2_X1 U694 ( .A1(n575), .A2(A[3]), .ZN(n377) );
  NAND2_X1 U695 ( .A1(A[23]), .A2(n425), .ZN(n137) );
  NOR2_X1 U696 ( .A1(A[23]), .A2(n425), .ZN(n136) );
  INV_X1 U697 ( .A(B[8]), .ZN(n440) );
  NAND2_X1 U698 ( .A1(A[6]), .A2(n442), .ZN(n358) );
  NOR2_X1 U699 ( .A1(A[7]), .A2(n441), .ZN(n346) );
  NAND2_X2 U700 ( .A1(n271), .A2(n167), .ZN(n165) );
  NOR2_X1 U701 ( .A1(A[5]), .A2(n443), .ZN(n364) );
  NAND2_X1 U702 ( .A1(A[5]), .A2(n443), .ZN(n365) );
  INV_X1 U703 ( .A(n186), .ZN(n398) );
  NOR2_X1 U704 ( .A1(A[19]), .A2(n429), .ZN(n186) );
  INV_X1 U705 ( .A(n42), .ZN(n40) );
  NOR2_X1 U706 ( .A1(A[16]), .A2(n432), .ZN(n229) );
  INV_X1 U707 ( .A(B[16]), .ZN(n432) );
  NAND2_X1 U708 ( .A1(A[16]), .A2(n432), .ZN(n230) );
  NAND2_X1 U709 ( .A1(n404), .A2(n263), .ZN(n23) );
  INV_X1 U710 ( .A(n263), .ZN(n261) );
  NOR2_X1 U711 ( .A1(A[13]), .A2(n435), .ZN(n262) );
  NAND2_X1 U712 ( .A1(A[13]), .A2(n435), .ZN(n263) );
  NOR2_X1 U713 ( .A1(A[17]), .A2(n431), .ZN(n210) );
  NOR2_X1 U714 ( .A1(A[15]), .A2(n433), .ZN(n238) );
  NAND2_X1 U715 ( .A1(n191), .A2(n398), .ZN(n180) );
  AOI21_X1 U716 ( .B1(n192), .B2(n398), .A(n185), .ZN(n181) );
  NAND2_X1 U717 ( .A1(n398), .A2(n187), .ZN(n17) );
  NOR2_X1 U718 ( .A1(n4), .A2(n143), .ZN(n141) );
  OAI21_X1 U719 ( .B1(n368), .B2(n143), .A(n567), .ZN(n142) );
  NAND2_X2 U720 ( .A1(n398), .A2(n397), .ZN(n173) );
  NOR2_X1 U721 ( .A1(A[20]), .A2(n428), .ZN(n177) );
  INV_X1 U722 ( .A(n571), .ZN(n114) );
  INV_X1 U723 ( .A(n570), .ZN(n62) );
  NAND2_X1 U724 ( .A1(A[12]), .A2(n436), .ZN(n286) );
  NOR2_X1 U725 ( .A1(A[12]), .A2(n436), .ZN(n285) );
  NOR2_X1 U726 ( .A1(A[9]), .A2(n439), .ZN(n318) );
  NAND2_X1 U727 ( .A1(A[9]), .A2(n439), .ZN(n319) );
  NAND2_X1 U728 ( .A1(A[11]), .A2(n437), .ZN(n295) );
  NOR2_X1 U729 ( .A1(A[11]), .A2(n437), .ZN(n294) );
  NAND2_X1 U730 ( .A1(n413), .A2(n154), .ZN(n152) );
  AOI21_X1 U731 ( .B1(n370), .B2(n154), .A(n568), .ZN(n153) );
  INV_X1 U732 ( .A(n553), .ZN(n113) );
  NAND2_X1 U733 ( .A1(n554), .A2(n91), .ZN(n89) );
  NAND2_X1 U734 ( .A1(n413), .A2(n52), .ZN(n50) );
  XNOR2_X1 U735 ( .A(n38), .B(n5), .ZN(DIFF[31]) );
  NAND2_X1 U736 ( .A1(A[8]), .A2(n440), .ZN(n338) );
  NOR2_X1 U737 ( .A1(A[8]), .A2(n440), .ZN(n337) );
  NAND2_X1 U738 ( .A1(A[10]), .A2(n438), .ZN(n310) );
  NOR2_X1 U739 ( .A1(A[10]), .A2(n438), .ZN(n309) );
  INV_X1 U740 ( .A(B[4]), .ZN(n574) );
  INV_X1 U741 ( .A(B[3]), .ZN(n575) );
  INV_X1 U742 ( .A(B[2]), .ZN(n576) );
  INV_X1 U743 ( .A(B[1]), .ZN(n577) );
  INV_X1 U744 ( .A(B[0]), .ZN(n578) );
  INV_X2 U745 ( .A(n98), .ZN(n96) );
  INV_X2 U746 ( .A(n94), .ZN(n92) );
  INV_X2 U747 ( .A(n93), .ZN(n91) );
  INV_X2 U748 ( .A(n88), .ZN(n86) );
  INV_X2 U749 ( .A(n87), .ZN(n85) );
  INV_X2 U750 ( .A(n83), .ZN(n81) );
  INV_X2 U751 ( .A(n74), .ZN(n72) );
  INV_X2 U752 ( .A(n48), .ZN(n46) );
  INV_X2 U753 ( .A(B[21]), .ZN(n427) );
  INV_X2 U754 ( .A(B[22]), .ZN(n426) );
  INV_X2 U755 ( .A(B[23]), .ZN(n425) );
  INV_X2 U756 ( .A(B[24]), .ZN(n424) );
  INV_X2 U757 ( .A(B[25]), .ZN(n423) );
  INV_X2 U758 ( .A(B[26]), .ZN(n422) );
  INV_X2 U759 ( .A(B[27]), .ZN(n421) );
  INV_X2 U760 ( .A(B[28]), .ZN(n420) );
  INV_X2 U761 ( .A(B[29]), .ZN(n419) );
  INV_X2 U762 ( .A(B[30]), .ZN(n418) );
  INV_X2 U763 ( .A(B[31]), .ZN(n417) );
  INV_X2 U764 ( .A(n383), .ZN(n416) );
  INV_X2 U765 ( .A(n379), .ZN(n415) );
  INV_X2 U766 ( .A(n376), .ZN(n414) );
  INV_X2 U767 ( .A(n158), .ZN(n396) );
  INV_X2 U768 ( .A(n97), .ZN(n95) );
  INV_X2 U769 ( .A(n82), .ZN(n80) );
  INV_X2 U770 ( .A(n73), .ZN(n71) );
  INV_X2 U771 ( .A(n56), .ZN(n388) );
  INV_X2 U772 ( .A(n47), .ZN(n45) );
  INV_X2 U773 ( .A(n36), .ZN(n386) );
  INV_X2 U774 ( .A(n382), .ZN(n381) );
  INV_X2 U775 ( .A(n368), .ZN(n370) );
  INV_X2 U776 ( .A(n4), .ZN(n413) );
  INV_X2 U777 ( .A(n364), .ZN(n412) );
  INV_X2 U778 ( .A(n355), .ZN(n353) );
  INV_X2 U779 ( .A(n352), .ZN(n350) );
  INV_X2 U780 ( .A(n351), .ZN(n349) );
  INV_X2 U781 ( .A(n338), .ZN(n336) );
  INV_X2 U782 ( .A(n337), .ZN(n409) );
  INV_X2 U783 ( .A(n324), .ZN(n322) );
  INV_X2 U784 ( .A(n323), .ZN(n321) );
  INV_X2 U785 ( .A(n319), .ZN(n317) );
  INV_X2 U786 ( .A(n318), .ZN(n408) );
  INV_X2 U787 ( .A(n310), .ZN(n308) );
  INV_X2 U788 ( .A(n306), .ZN(n304) );
  INV_X2 U789 ( .A(n305), .ZN(n303) );
  INV_X2 U790 ( .A(n300), .ZN(n298) );
  INV_X2 U791 ( .A(n299), .ZN(n297) );
  INV_X2 U792 ( .A(n295), .ZN(n293) );
  INV_X2 U793 ( .A(n294), .ZN(n406) );
  INV_X2 U794 ( .A(n286), .ZN(n284) );
  INV_X2 U795 ( .A(n280), .ZN(n278) );
  INV_X2 U796 ( .A(n268), .ZN(n266) );
  INV_X2 U797 ( .A(n267), .ZN(n265) );
  INV_X2 U798 ( .A(n262), .ZN(n404) );
  INV_X2 U799 ( .A(n253), .ZN(n403) );
  INV_X2 U800 ( .A(n249), .ZN(n247) );
  INV_X2 U801 ( .A(n244), .ZN(n242) );
  INV_X2 U802 ( .A(n243), .ZN(n241) );
  INV_X2 U803 ( .A(n239), .ZN(n237) );
  INV_X2 U804 ( .A(n238), .ZN(n402) );
  INV_X2 U805 ( .A(n230), .ZN(n228) );
  INV_X2 U806 ( .A(n220), .ZN(n218) );
  INV_X2 U807 ( .A(n219), .ZN(n217) );
  INV_X2 U808 ( .A(n216), .ZN(n214) );
  INV_X2 U809 ( .A(n215), .ZN(n213) );
  INV_X2 U810 ( .A(n210), .ZN(n400) );
  INV_X2 U811 ( .A(n197), .ZN(n195) );
  INV_X2 U812 ( .A(n192), .ZN(n190) );
  INV_X2 U813 ( .A(n191), .ZN(n189) );
  INV_X2 U814 ( .A(n187), .ZN(n185) );
  INV_X2 U815 ( .A(n177), .ZN(n397) );
  INV_X2 U816 ( .A(n169), .ZN(n167) );
  INV_X2 U817 ( .A(n165), .ZN(n163) );
  INV_X2 U818 ( .A(n150), .ZN(n148) );
  INV_X2 U819 ( .A(n149), .ZN(n395) );
  INV_X2 U820 ( .A(n137), .ZN(n135) );
  INV_X2 U821 ( .A(n136), .ZN(n394) );
  INV_X2 U822 ( .A(n128), .ZN(n126) );
  INV_X2 U823 ( .A(n127), .ZN(n393) );
  INV_X2 U824 ( .A(n111), .ZN(n109) );
  INV_X2 U825 ( .A(n107), .ZN(n105) );
  INV_X2 U826 ( .A(n106), .ZN(n392) );
endmodule


module Xi_core_DW01_add_1 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] ;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X2 U1 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X2 U2 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U3 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  AND2_X1 U4 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  XOR2_X1 U5 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  AND2_X1 U6 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U7 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U8 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  XOR2_X1 U9 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  AND2_X1 U10 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  XOR2_X1 U11 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  AND2_X1 U12 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  XOR2_X1 U13 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  AND2_X1 U14 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  XOR2_X1 U15 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  AND2_X1 U16 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  XOR2_X1 U17 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  AND2_X1 U18 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  XOR2_X1 U19 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  AND2_X1 U20 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  XOR2_X1 U21 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  XOR2_X1 U23 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  AND2_X1 U24 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  XOR2_X1 U25 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  AND2_X1 U26 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  XOR2_X1 U27 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  AND2_X1 U28 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  XOR2_X1 U29 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  AND2_X1 U30 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  XOR2_X1 U31 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  AND2_X1 U32 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  XOR2_X1 U33 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  AND2_X1 U34 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  XOR2_X1 U35 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  AND2_X1 U36 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  XOR2_X1 U37 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  AND2_X1 U38 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  XOR2_X1 U39 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  AND2_X1 U40 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  XOR2_X1 U41 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  INV_X1 U42 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module Xi_core_DW01_add_0 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;
  wire   \carry[19] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[2] ,
         \carry[1] , net56331, net56330, net56329, net56383, net57063,
         net57069, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(n53), .CO(\carry[9] ), .S(SUM[8]) );
  XNOR2_X2 syn249 ( .A(A[23]), .B(B[23]), .ZN(n19) );
  NAND2_X2 syn241 ( .A1(n17), .A2(n18), .ZN(n25) );
  NAND2_X2 syn237 ( .A1(n15), .A2(n16), .ZN(n24) );
  NAND2_X2 syn235 ( .A1(A[21]), .A2(B[21]), .ZN(n22) );
  NAND2_X2 syn233 ( .A1(A[22]), .A2(B[22]), .ZN(n23) );
  XNOR2_X2 syn201 ( .A(net57063), .B(n21), .ZN(SUM[22]) );
  XNOR2_X2 syn198 ( .A(A[22]), .B(n18), .ZN(net56383) );
  XNOR2_X2 syn179 ( .A(A[21]), .B(B[21]), .ZN(net57069) );
  NAND3_X1 syn145 ( .A1(net56330), .A2(net56331), .A3(net56329), .ZN(n14) );
  INV_X2 syn21 ( .A(B[22]), .ZN(n18) );
  INV_X2 syn20 ( .A(A[22]), .ZN(n17) );
  INV_X2 syn16 ( .A(A[21]), .ZN(n16) );
  INV_X2 syn15 ( .A(B[21]), .ZN(n15) );
  INV_X1 U1 ( .A(n149), .ZN(n13) );
  NAND2_X1 U2 ( .A1(n14), .A2(n4), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n1), .A2(n2), .ZN(n20) );
  OR2_X1 U4 ( .A1(n3), .A2(n11), .ZN(n2) );
  INV_X1 U5 ( .A(n9), .ZN(n3) );
  AND2_X1 U6 ( .A1(n24), .A2(n9), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n14), .A2(n24), .ZN(n5) );
  NAND2_X1 U8 ( .A1(n50), .A2(B[15]), .ZN(n6) );
  NAND3_X1 U9 ( .A1(net56330), .A2(net56331), .A3(net56329), .ZN(n7) );
  NAND2_X1 U10 ( .A1(n5), .A2(n22), .ZN(n21) );
  NAND2_X1 U11 ( .A1(n34), .A2(B[10]), .ZN(n8) );
  OR2_X1 U12 ( .A1(n10), .A2(n25), .ZN(n9) );
  INV_X1 U13 ( .A(n23), .ZN(n10) );
  AND2_X1 U14 ( .A1(n22), .A2(n23), .ZN(n11) );
  CLKBUF_X1 U15 ( .A(n92), .Z(n12) );
  NAND2_X1 U16 ( .A1(\carry[6] ), .A2(A[6]), .ZN(n92) );
  XNOR2_X1 U17 ( .A(n94), .B(n13), .ZN(SUM[20]) );
  XNOR2_X1 U18 ( .A(n19), .B(n20), .ZN(SUM[23]) );
  NAND2_X1 U19 ( .A1(n128), .A2(A[14]), .ZN(n26) );
  NAND2_X1 U20 ( .A1(n66), .A2(B[6]), .ZN(n91) );
  NAND2_X1 U21 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n27) );
  NAND2_X1 U22 ( .A1(n36), .A2(B[19]), .ZN(n148) );
  NAND3_X1 U23 ( .A1(n148), .A2(n147), .A3(n146), .ZN(n28) );
  CLKBUF_X1 U24 ( .A(B[5]), .Z(n29) );
  NAND2_X1 U25 ( .A1(\carry[15] ), .A2(A[15]), .ZN(n30) );
  NAND2_X1 U26 ( .A1(\carry[15] ), .A2(A[15]), .ZN(n142) );
  CLKBUF_X1 U27 ( .A(n30), .Z(n31) );
  NAND3_X1 U28 ( .A1(n119), .A2(n118), .A3(n117), .ZN(n32) );
  NAND3_X1 U29 ( .A1(n119), .A2(n118), .A3(n117), .ZN(n51) );
  CLKBUF_X1 U30 ( .A(n32), .Z(n33) );
  NAND3_X1 U31 ( .A1(n153), .A2(n152), .A3(n151), .ZN(n34) );
  CLKBUF_X1 U32 ( .A(n148), .Z(n35) );
  NAND3_X1 U33 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n36) );
  NAND2_X1 U34 ( .A1(n51), .A2(A[18]), .ZN(n60) );
  CLKBUF_X1 U35 ( .A(n36), .Z(n37) );
  NAND3_X1 U36 ( .A1(n59), .A2(n60), .A3(n61), .ZN(\carry[19] ) );
  NAND2_X1 U37 ( .A1(n43), .A2(B[16]), .ZN(n38) );
  NAND2_X1 U38 ( .A1(n43), .A2(B[16]), .ZN(n115) );
  NAND2_X1 U39 ( .A1(n110), .A2(A[16]), .ZN(n39) );
  NAND2_X1 U40 ( .A1(n110), .A2(A[16]), .ZN(n114) );
  NAND3_X1 U41 ( .A1(n152), .A2(n153), .A3(n151), .ZN(\carry[10] ) );
  NAND3_X1 U42 ( .A1(n38), .A2(n39), .A3(n113), .ZN(n40) );
  NAND2_X1 U43 ( .A1(\carry[12] ), .A2(A[12]), .ZN(n41) );
  NAND2_X1 U44 ( .A1(\carry[12] ), .A2(A[12]), .ZN(n131) );
  NAND2_X1 U45 ( .A1(n55), .A2(A[13]), .ZN(n42) );
  NAND3_X1 U46 ( .A1(n30), .A2(n143), .A3(n141), .ZN(n43) );
  NAND3_X1 U47 ( .A1(n165), .A2(n163), .A3(n164), .ZN(n44) );
  NAND2_X1 U48 ( .A1(\carry[8] ), .A2(B[8]), .ZN(n45) );
  NAND2_X1 U49 ( .A1(\carry[8] ), .A2(A[8]), .ZN(n46) );
  NAND2_X1 U50 ( .A1(B[8]), .A2(A[8]), .ZN(n47) );
  NAND3_X1 U51 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n56) );
  CLKBUF_X1 U52 ( .A(n27), .Z(n62) );
  NAND3_X1 U53 ( .A1(n109), .A2(n108), .A3(n107), .ZN(\carry[5] ) );
  NAND2_X1 U54 ( .A1(\carry[7] ), .A2(A[7]), .ZN(n48) );
  CLKBUF_X1 U55 ( .A(n39), .Z(n49) );
  NAND3_X1 U56 ( .A1(n26), .A2(n139), .A3(n137), .ZN(n50) );
  CLKBUF_X1 U57 ( .A(\carry[15] ), .Z(n52) );
  NAND3_X1 U58 ( .A1(n71), .A2(n48), .A3(n72), .ZN(n53) );
  NAND3_X1 U59 ( .A1(n138), .A2(n137), .A3(n139), .ZN(\carry[15] ) );
  NAND3_X1 U60 ( .A1(n71), .A2(n48), .A3(n72), .ZN(\carry[8] ) );
  NAND3_X1 U61 ( .A1(n6), .A2(n142), .A3(n141), .ZN(n110) );
  NAND3_X1 U62 ( .A1(n148), .A2(n27), .A3(n146), .ZN(n54) );
  NAND3_X1 U63 ( .A1(n132), .A2(n131), .A3(n130), .ZN(n55) );
  CLKBUF_X1 U64 ( .A(n6), .Z(n57) );
  XOR2_X1 U65 ( .A(B[18]), .B(A[18]), .Z(n58) );
  XOR2_X1 U66 ( .A(n33), .B(n58), .Z(SUM[18]) );
  NAND2_X1 U67 ( .A1(n32), .A2(B[18]), .ZN(n59) );
  NAND2_X1 U68 ( .A1(B[18]), .A2(A[18]), .ZN(n61) );
  CLKBUF_X1 U69 ( .A(n38), .Z(n63) );
  NAND3_X1 U70 ( .A1(n157), .A2(n156), .A3(n155), .ZN(n64) );
  NAND3_X1 U71 ( .A1(n8), .A2(n156), .A3(n155), .ZN(\carry[11] ) );
  CLKBUF_X1 U72 ( .A(n91), .Z(n65) );
  NAND3_X1 U73 ( .A1(n87), .A2(n88), .A3(n89), .ZN(n66) );
  NAND3_X1 U74 ( .A1(n88), .A2(n89), .A3(n87), .ZN(\carry[6] ) );
  CLKBUF_X1 U75 ( .A(n108), .Z(n67) );
  CLKBUF_X1 U76 ( .A(n41), .Z(n68) );
  NAND3_X1 U77 ( .A1(n124), .A2(n125), .A3(n126), .ZN(n69) );
  NAND2_X1 U78 ( .A1(A[3]), .A2(B[3]), .ZN(n103) );
  XOR2_X1 U79 ( .A(B[7]), .B(A[7]), .Z(n70) );
  XOR2_X1 U80 ( .A(n74), .B(n70), .Z(SUM[7]) );
  NAND2_X1 U81 ( .A1(n73), .A2(B[7]), .ZN(n71) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(A[7]), .ZN(n72) );
  NAND3_X1 U83 ( .A1(n65), .A2(n12), .A3(n93), .ZN(n74) );
  NAND3_X1 U84 ( .A1(n91), .A2(n92), .A3(n93), .ZN(n73) );
  CLKBUF_X1 U85 ( .A(B[1]), .Z(n75) );
  CLKBUF_X1 U86 ( .A(\carry[12] ), .Z(n76) );
  NAND3_X1 U87 ( .A1(n124), .A2(n125), .A3(n126), .ZN(\carry[12] ) );
  CLKBUF_X1 U88 ( .A(n128), .Z(n77) );
  CLKBUF_X1 U89 ( .A(n66), .Z(n78) );
  NAND2_X1 U90 ( .A1(n83), .A2(A[4]), .ZN(n108) );
  CLKBUF_X1 U91 ( .A(n34), .Z(n79) );
  CLKBUF_X1 U92 ( .A(n56), .Z(n80) );
  CLKBUF_X1 U93 ( .A(n132), .Z(n81) );
  NAND2_X1 U94 ( .A1(n97), .A2(A[1]), .ZN(n82) );
  NAND2_X1 U95 ( .A1(n97), .A2(A[1]), .ZN(n160) );
  NAND3_X1 U96 ( .A1(n105), .A2(n104), .A3(n103), .ZN(n83) );
  NAND3_X1 U97 ( .A1(n105), .A2(n104), .A3(n103), .ZN(n99) );
  CLKBUF_X1 U98 ( .A(n109), .Z(n84) );
  NAND3_X1 U99 ( .A1(n84), .A2(n67), .A3(n107), .ZN(n85) );
  XOR2_X1 U100 ( .A(n29), .B(A[5]), .Z(n86) );
  XOR2_X1 U101 ( .A(n85), .B(n86), .Z(SUM[5]) );
  NAND2_X1 U102 ( .A1(\carry[5] ), .A2(B[5]), .ZN(n87) );
  NAND2_X1 U103 ( .A1(\carry[5] ), .A2(A[5]), .ZN(n88) );
  NAND2_X1 U104 ( .A1(B[5]), .A2(A[5]), .ZN(n89) );
  XOR2_X1 U105 ( .A(B[6]), .B(A[6]), .Z(n90) );
  XOR2_X1 U106 ( .A(n78), .B(n90), .Z(SUM[6]) );
  NAND2_X1 U107 ( .A1(B[6]), .A2(A[6]), .ZN(n93) );
  NAND3_X1 U108 ( .A1(n91), .A2(n92), .A3(n93), .ZN(\carry[7] ) );
  XNOR2_X1 U109 ( .A(n7), .B(net57069), .ZN(SUM[21]) );
  INV_X32 U110 ( .A(net56383), .ZN(net57063) );
  NAND3_X1 U111 ( .A1(n62), .A2(n146), .A3(n35), .ZN(n94) );
  NAND2_X1 U112 ( .A1(\carry[11] ), .A2(A[11]), .ZN(n125) );
  CLKBUF_X1 U113 ( .A(n64), .Z(n95) );
  NAND3_X1 U114 ( .A1(n165), .A2(n164), .A3(n163), .ZN(n96) );
  AND2_X1 U115 ( .A1(B[0]), .A2(A[0]), .ZN(n97) );
  AND2_X1 U116 ( .A1(B[0]), .A2(A[0]), .ZN(\carry[1] ) );
  CLKBUF_X1 U117 ( .A(n97), .Z(n98) );
  CLKBUF_X1 U118 ( .A(n99), .Z(n100) );
  CLKBUF_X1 U119 ( .A(n44), .Z(n101) );
  XOR2_X1 U120 ( .A(A[3]), .B(B[3]), .Z(n102) );
  XOR2_X1 U121 ( .A(n102), .B(n101), .Z(SUM[3]) );
  NAND2_X1 U122 ( .A1(n96), .A2(A[3]), .ZN(n104) );
  NAND2_X1 U123 ( .A1(n44), .A2(B[3]), .ZN(n105) );
  XOR2_X1 U124 ( .A(A[4]), .B(B[4]), .Z(n106) );
  XOR2_X1 U125 ( .A(n106), .B(n100), .Z(SUM[4]) );
  NAND2_X1 U126 ( .A1(A[4]), .A2(B[4]), .ZN(n107) );
  NAND2_X1 U127 ( .A1(n99), .A2(B[4]), .ZN(n109) );
  NAND3_X1 U128 ( .A1(n57), .A2(n141), .A3(n31), .ZN(\carry[16] ) );
  NAND3_X1 U129 ( .A1(n63), .A2(n113), .A3(n49), .ZN(n111) );
  NAND3_X1 U130 ( .A1(n115), .A2(n114), .A3(n113), .ZN(\carry[17] ) );
  XOR2_X1 U131 ( .A(A[16]), .B(B[16]), .Z(n112) );
  XOR2_X1 U132 ( .A(\carry[16] ), .B(n112), .Z(SUM[16]) );
  NAND2_X1 U133 ( .A1(A[16]), .A2(B[16]), .ZN(n113) );
  XOR2_X1 U134 ( .A(A[17]), .B(B[17]), .Z(n116) );
  XOR2_X1 U135 ( .A(n116), .B(n111), .Z(SUM[17]) );
  NAND2_X1 U136 ( .A1(A[17]), .A2(B[17]), .ZN(n117) );
  NAND2_X1 U137 ( .A1(\carry[17] ), .A2(A[17]), .ZN(n118) );
  NAND2_X1 U138 ( .A1(n40), .A2(B[17]), .ZN(n119) );
  NAND3_X1 U139 ( .A1(n161), .A2(n160), .A3(n159), .ZN(n120) );
  CLKBUF_X1 U140 ( .A(n120), .Z(n121) );
  NAND3_X1 U141 ( .A1(n82), .A2(n161), .A3(n159), .ZN(\carry[2] ) );
  NAND2_X1 U142 ( .A1(B[1]), .A2(A[1]), .ZN(n159) );
  NAND3_X1 U143 ( .A1(n130), .A2(n68), .A3(n81), .ZN(n122) );
  XOR2_X1 U144 ( .A(B[11]), .B(A[11]), .Z(n123) );
  XOR2_X1 U145 ( .A(n95), .B(n123), .Z(SUM[11]) );
  NAND2_X1 U146 ( .A1(n64), .A2(B[11]), .ZN(n124) );
  NAND2_X1 U147 ( .A1(B[11]), .A2(A[11]), .ZN(n126) );
  CLKBUF_X1 U148 ( .A(B[0]), .Z(n127) );
  NAND3_X1 U149 ( .A1(n41), .A2(n132), .A3(n130), .ZN(\carry[13] ) );
  NAND3_X1 U150 ( .A1(n135), .A2(n42), .A3(n134), .ZN(n128) );
  NAND3_X1 U151 ( .A1(n135), .A2(n134), .A3(n42), .ZN(\carry[14] ) );
  XOR2_X1 U152 ( .A(A[12]), .B(B[12]), .Z(n129) );
  XOR2_X1 U153 ( .A(n76), .B(n129), .Z(SUM[12]) );
  NAND2_X2 U154 ( .A1(A[12]), .A2(B[12]), .ZN(n130) );
  NAND2_X1 U155 ( .A1(n69), .A2(B[12]), .ZN(n132) );
  XOR2_X1 U156 ( .A(A[13]), .B(B[13]), .Z(n133) );
  XOR2_X1 U157 ( .A(n133), .B(n122), .Z(SUM[13]) );
  NAND2_X1 U158 ( .A1(A[13]), .A2(B[13]), .ZN(n134) );
  NAND2_X1 U159 ( .A1(\carry[13] ), .A2(B[13]), .ZN(n135) );
  XOR2_X1 U160 ( .A(A[14]), .B(B[14]), .Z(n136) );
  XOR2_X1 U161 ( .A(n77), .B(n136), .Z(SUM[14]) );
  NAND2_X2 U162 ( .A1(A[14]), .A2(B[14]), .ZN(n137) );
  NAND2_X1 U163 ( .A1(n128), .A2(A[14]), .ZN(n138) );
  NAND2_X1 U164 ( .A1(\carry[14] ), .A2(B[14]), .ZN(n139) );
  XOR2_X1 U165 ( .A(A[15]), .B(B[15]), .Z(n140) );
  XOR2_X1 U166 ( .A(n52), .B(n140), .Z(SUM[15]) );
  NAND2_X1 U167 ( .A1(A[15]), .A2(B[15]), .ZN(n141) );
  NAND2_X1 U168 ( .A1(n50), .A2(B[15]), .ZN(n143) );
  CLKBUF_X1 U169 ( .A(B[2]), .Z(n144) );
  XOR2_X1 U170 ( .A(A[19]), .B(B[19]), .Z(n145) );
  XOR2_X1 U171 ( .A(n37), .B(n145), .Z(SUM[19]) );
  NAND2_X1 U172 ( .A1(A[19]), .A2(B[19]), .ZN(n146) );
  NAND2_X1 U173 ( .A1(\carry[19] ), .A2(A[19]), .ZN(n147) );
  XOR2_X1 U174 ( .A(A[20]), .B(B[20]), .Z(n149) );
  NAND2_X1 U175 ( .A1(A[20]), .A2(B[20]), .ZN(net56329) );
  NAND2_X1 U176 ( .A1(n28), .A2(A[20]), .ZN(net56330) );
  NAND2_X1 U177 ( .A1(n54), .A2(B[20]), .ZN(net56331) );
  XOR2_X1 U178 ( .A(A[9]), .B(B[9]), .Z(n150) );
  XOR2_X1 U179 ( .A(n150), .B(n80), .Z(SUM[9]) );
  NAND2_X2 U180 ( .A1(A[9]), .A2(B[9]), .ZN(n151) );
  NAND2_X1 U181 ( .A1(n56), .A2(A[9]), .ZN(n152) );
  NAND2_X1 U182 ( .A1(\carry[9] ), .A2(B[9]), .ZN(n153) );
  XOR2_X1 U183 ( .A(A[10]), .B(B[10]), .Z(n154) );
  XOR2_X1 U184 ( .A(n154), .B(n79), .Z(SUM[10]) );
  NAND2_X1 U185 ( .A1(A[10]), .A2(B[10]), .ZN(n155) );
  NAND2_X1 U186 ( .A1(\carry[10] ), .A2(A[10]), .ZN(n156) );
  NAND2_X1 U187 ( .A1(n34), .A2(B[10]), .ZN(n157) );
  XOR2_X1 U188 ( .A(A[1]), .B(n75), .Z(n158) );
  XOR2_X1 U189 ( .A(n158), .B(n98), .Z(SUM[1]) );
  NAND2_X1 U190 ( .A1(\carry[1] ), .A2(B[1]), .ZN(n161) );
  XOR2_X1 U191 ( .A(A[2]), .B(n144), .Z(n162) );
  XOR2_X1 U192 ( .A(n162), .B(n121), .Z(SUM[2]) );
  NAND2_X1 U193 ( .A1(B[2]), .A2(A[2]), .ZN(n163) );
  NAND2_X1 U194 ( .A1(\carry[2] ), .A2(A[2]), .ZN(n164) );
  NAND2_X1 U195 ( .A1(n120), .A2(B[2]), .ZN(n165) );
  XOR2_X1 U196 ( .A(n127), .B(A[0]), .Z(SUM[0]) );
endmodule


module Xi_core ( CLK, reset, reboot, freeze, I_NREADY, D_NREADY, I_BUSY, 
        D_BUSY, INTERRUPT_VECTOR, I_ADDR_OUTBUS, I_DATA_INBUS, D_ADDR_OUTBUS, 
        D_DATA_INBUS, D_DATA_OUTBUS, mem_read, mem_write, mem_isbyte, 
        mem_ishalf, dbg_enable, ext_bp_request, end_dbg, real_dbg_op, 
        kernel_mode, suspend );
  input [7:0] INTERRUPT_VECTOR;
  output [23:0] I_ADDR_OUTBUS;
  input [31:0] I_DATA_INBUS;
  output [31:0] D_ADDR_OUTBUS;
  input [31:0] D_DATA_INBUS;
  output [31:0] D_DATA_OUTBUS;
  input CLK, reset, reboot, freeze, I_NREADY, D_NREADY, dbg_enable,
         ext_bp_request;
  output I_BUSY, D_BUSY, mem_read, mem_write, mem_isbyte, mem_ishalf, end_dbg,
         real_dbg_op, kernel_mode, suspend;
  wire   n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, serve_exception,
         \x_mem_command[MB] , \x_mem_command[MH] , \x_mem_command[MR] ,
         \x_mem_command[MW] , N5, \exc[ALU_OFLOW1] , \exc[DMEM_MISALIGN] ,
         \Alu_command[OP][5] , \Alu_command[OP][4] , \Alu_command[OP][3] ,
         \Alu_command[OP][2] , \Alu_command[OP][1] , \Alu_command[OP][0] ,
         m_we, \m_mem_command[MR] , \m_mem_command[SIGN] , N80, dcheck_enable,
         N82, N83, \Scc_coproc/N601 , \Scc_coproc/N600 , \Scc_coproc/N599 ,
         \Scc_coproc/N587 , \Scc_coproc/N586 , \Scc_coproc/N585 ,
         \Scc_coproc/N584 , \Scc_coproc/N583 , \Scc_coproc/N582 ,
         \Scc_coproc/N580 , \Scc_coproc/N579 , \Scc_coproc/N578 ,
         \Scc_coproc/N577 , \Scc_coproc/N576 , \Scc_coproc/N575 ,
         \Scc_coproc/N574 , \Scc_coproc/N573 , \Scc_coproc/N572 ,
         \Scc_coproc/N571 , \Scc_coproc/N562 , \Scc_coproc/N553 ,
         \Scc_coproc/N551 , \Scc_coproc/cause[4] , \Scc_coproc/cause[5] ,
         \Scc_coproc/interrupt_active , \Scc_coproc/interrupt[2] ,
         \Scc_coproc/interrupt[3] , \Scc_coproc/interrupt[4] ,
         \Scc_coproc/interrupt[5] , \Scc_coproc/interrupt[6] ,
         \Scc_coproc/interrupt[7] , \Scc_coproc/interrupt[8] ,
         \Scc_coproc/interrupt[9] , \Scc_coproc/x_exc_word[0] ,
         \Scc_coproc/x_exc_word[1] , \Scc_coproc/x_exc_word[2] ,
         \Scc_coproc/x_exc_word[3] , \Scc_coproc/x_exc_word[4] ,
         \Scc_coproc/x_exc_word[5] , \Scc_coproc/x_status[14] ,
         \Scc_coproc/ein_exc_word[0] , \Scc_coproc/ein_exc_word[1] ,
         \Scc_coproc/ein_exc_word[2] , \Scc_coproc/ein_exc_word[3] ,
         \Scc_coproc/ein_exc_word[4] , \Scc_coproc/ein_exc_word[5] ,
         \Scc_coproc/din_exc_word[0] , \Scc_coproc/din_exc_word[4] ,
         \Scc_coproc/din_exc_word[5] , \Scc_coproc/status[2] , \regfile/N456 ,
         \regfile/N455 , \regfile/N444 , \regfile/N438 , \regfile/N433 ,
         \regfile/N432 , \regfile/N427 , \regfile/N426 , \regfile/N421 ,
         \regfile/N420 , \regfile/N415 , \regfile/N414 , \regfile/N409 ,
         \regfile/N402 , \regfile/N397 , \regfile/N396 , \regfile/N391 ,
         \regfile/N390 , \regfile/N385 , \regfile/N384 , \regfile/N379 ,
         \regfile/N378 , \regfile/N372 , \regfile/N367 , \regfile/N366 ,
         \regfile/N360 , \regfile/N359 , \regfile/N358 , \regfile/N353 ,
         \regfile/N347 , \regfile/N342 , \regfile/N341 , \regfile/N336 ,
         \regfile/N335 , \regfile/N329 , \regfile/N324 , \regfile/N323 ,
         \regfile/N318 , \regfile/N317 , \regfile/N315 , \regfile/N311 ,
         \regfile/N310 , \regfile/N304 , \regfile/N299 , \regfile/N298 ,
         \regfile/N293 , \regfile/N292 , \regfile/N290 , \regfile/N286 ,
         \regfile/N285 , \regfile/N279 , \regfile/N273 , \regfile/N272 ,
         \regfile/N269 , \regfile/N267 , \regfile/N266 , \regfile/N265 ,
         \regfile/N264 , \regfile/N262 , \regfile/N261 , \regfile/N260 ,
         \regfile/reg_out[16][0] , \regfile/reg_out[16][1] ,
         \regfile/reg_out[16][2] , \regfile/reg_out[16][3] ,
         \regfile/reg_out[16][4] , \regfile/reg_out[16][5] ,
         \regfile/reg_out[16][6] , \regfile/reg_out[16][7] ,
         \regfile/reg_out[16][8] , \regfile/reg_out[16][9] ,
         \regfile/reg_out[16][10] , \regfile/reg_out[16][11] ,
         \regfile/reg_out[16][12] , \regfile/reg_out[16][13] ,
         \regfile/reg_out[16][14] , \regfile/reg_out[16][15] ,
         \regfile/reg_out[16][16] , \regfile/reg_out[16][17] ,
         \regfile/reg_out[16][18] , \regfile/reg_out[16][19] ,
         \regfile/reg_out[16][20] , \regfile/reg_out[16][21] ,
         \regfile/reg_out[16][22] , \regfile/reg_out[16][23] ,
         \regfile/reg_out[16][24] , \regfile/reg_out[16][25] ,
         \regfile/reg_out[16][26] , \regfile/reg_out[16][27] ,
         \regfile/reg_out[16][28] , \regfile/reg_out[16][29] ,
         \regfile/reg_out[16][30] , \regfile/reg_out[16][31] ,
         \regfile/reg_out[17][0] , \regfile/reg_out[17][1] ,
         \regfile/reg_out[17][2] , \regfile/reg_out[17][3] ,
         \regfile/reg_out[17][4] , \regfile/reg_out[17][5] ,
         \regfile/reg_out[17][6] , \regfile/reg_out[17][7] ,
         \regfile/reg_out[17][8] , \regfile/reg_out[17][9] ,
         \regfile/reg_out[17][10] , \regfile/reg_out[17][11] ,
         \regfile/reg_out[17][12] , \regfile/reg_out[17][13] ,
         \regfile/reg_out[17][14] , \regfile/reg_out[17][15] ,
         \regfile/reg_out[17][16] , \regfile/reg_out[17][17] ,
         \regfile/reg_out[17][18] , \regfile/reg_out[17][19] ,
         \regfile/reg_out[17][20] , \regfile/reg_out[17][21] ,
         \regfile/reg_out[17][22] , \regfile/reg_out[17][23] ,
         \regfile/reg_out[17][24] , \regfile/reg_out[17][25] ,
         \regfile/reg_out[17][26] , \regfile/reg_out[17][27] ,
         \regfile/reg_out[17][28] , \regfile/reg_out[17][29] ,
         \regfile/reg_out[17][30] , \regfile/reg_out[17][31] ,
         \regfile/reg_out[18][0] , \regfile/reg_out[18][1] ,
         \regfile/reg_out[18][2] , \regfile/reg_out[18][3] ,
         \regfile/reg_out[18][4] , \regfile/reg_out[18][5] ,
         \regfile/reg_out[18][6] , \regfile/reg_out[18][7] ,
         \regfile/reg_out[18][8] , \regfile/reg_out[18][9] ,
         \regfile/reg_out[18][10] , \regfile/reg_out[18][11] ,
         \regfile/reg_out[18][12] , \regfile/reg_out[18][13] ,
         \regfile/reg_out[18][14] , \regfile/reg_out[18][15] ,
         \regfile/reg_out[18][16] , \regfile/reg_out[18][17] ,
         \regfile/reg_out[18][18] , \regfile/reg_out[18][19] ,
         \regfile/reg_out[18][20] , \regfile/reg_out[18][21] ,
         \regfile/reg_out[18][22] , \regfile/reg_out[18][23] ,
         \regfile/reg_out[18][24] , \regfile/reg_out[18][25] ,
         \regfile/reg_out[18][26] , \regfile/reg_out[18][27] ,
         \regfile/reg_out[18][28] , \regfile/reg_out[18][29] ,
         \regfile/reg_out[18][30] , \regfile/reg_out[18][31] ,
         \regfile/reg_out[19][0] , \regfile/reg_out[19][1] ,
         \regfile/reg_out[19][2] , \regfile/reg_out[19][3] ,
         \regfile/reg_out[19][4] , \regfile/reg_out[19][5] ,
         \regfile/reg_out[19][6] , \regfile/reg_out[19][7] ,
         \regfile/reg_out[19][8] , \regfile/reg_out[19][9] ,
         \regfile/reg_out[19][10] , \regfile/reg_out[19][11] ,
         \regfile/reg_out[19][12] , \regfile/reg_out[19][13] ,
         \regfile/reg_out[19][14] , \regfile/reg_out[19][15] ,
         \regfile/reg_out[19][16] , \regfile/reg_out[19][17] ,
         \regfile/reg_out[19][18] , \regfile/reg_out[19][19] ,
         \regfile/reg_out[19][20] , \regfile/reg_out[19][21] ,
         \regfile/reg_out[19][22] , \regfile/reg_out[19][23] ,
         \regfile/reg_out[19][24] , \regfile/reg_out[19][25] ,
         \regfile/reg_out[19][26] , \regfile/reg_out[19][27] ,
         \regfile/reg_out[19][28] , \regfile/reg_out[19][29] ,
         \regfile/reg_out[19][30] , \regfile/reg_out[19][31] ,
         \regfile/reg_out[20][0] , \regfile/reg_out[20][1] ,
         \regfile/reg_out[20][2] , \regfile/reg_out[20][3] ,
         \regfile/reg_out[20][4] , \regfile/reg_out[20][5] ,
         \regfile/reg_out[20][6] , \regfile/reg_out[20][7] ,
         \regfile/reg_out[20][8] , \regfile/reg_out[20][9] ,
         \regfile/reg_out[20][10] , \regfile/reg_out[20][11] ,
         \regfile/reg_out[20][12] , \regfile/reg_out[20][13] ,
         \regfile/reg_out[20][14] , \regfile/reg_out[20][15] ,
         \regfile/reg_out[20][16] , \regfile/reg_out[20][17] ,
         \regfile/reg_out[20][18] , \regfile/reg_out[20][19] ,
         \regfile/reg_out[20][20] , \regfile/reg_out[20][21] ,
         \regfile/reg_out[20][22] , \regfile/reg_out[20][23] ,
         \regfile/reg_out[20][24] , \regfile/reg_out[20][25] ,
         \regfile/reg_out[20][26] , \regfile/reg_out[20][27] ,
         \regfile/reg_out[20][28] , \regfile/reg_out[20][29] ,
         \regfile/reg_out[20][30] , \regfile/reg_out[20][31] ,
         \regfile/reg_out[21][0] , \regfile/reg_out[21][1] ,
         \regfile/reg_out[21][2] , \regfile/reg_out[21][3] ,
         \regfile/reg_out[21][4] , \regfile/reg_out[21][5] ,
         \regfile/reg_out[21][6] , \regfile/reg_out[21][7] ,
         \regfile/reg_out[21][8] , \regfile/reg_out[21][9] ,
         \regfile/reg_out[21][10] , \regfile/reg_out[21][11] ,
         \regfile/reg_out[21][12] , \regfile/reg_out[21][13] ,
         \regfile/reg_out[21][14] , \regfile/reg_out[21][15] ,
         \regfile/reg_out[21][16] , \regfile/reg_out[21][17] ,
         \regfile/reg_out[21][18] , \regfile/reg_out[21][19] ,
         \regfile/reg_out[21][20] , \regfile/reg_out[21][21] ,
         \regfile/reg_out[21][22] , \regfile/reg_out[21][23] ,
         \regfile/reg_out[21][24] , \regfile/reg_out[21][25] ,
         \regfile/reg_out[21][26] , \regfile/reg_out[21][27] ,
         \regfile/reg_out[21][28] , \regfile/reg_out[21][29] ,
         \regfile/reg_out[21][30] , \regfile/reg_out[21][31] ,
         \regfile/reg_out[22][0] , \regfile/reg_out[22][1] ,
         \regfile/reg_out[22][2] , \regfile/reg_out[22][3] ,
         \regfile/reg_out[22][4] , \regfile/reg_out[22][5] ,
         \regfile/reg_out[22][6] , \regfile/reg_out[22][7] ,
         \regfile/reg_out[22][8] , \regfile/reg_out[22][9] ,
         \regfile/reg_out[22][10] , \regfile/reg_out[22][11] ,
         \regfile/reg_out[22][12] , \regfile/reg_out[22][13] ,
         \regfile/reg_out[22][14] , \regfile/reg_out[22][15] ,
         \regfile/reg_out[22][16] , \regfile/reg_out[22][17] ,
         \regfile/reg_out[22][18] , \regfile/reg_out[22][19] ,
         \regfile/reg_out[22][20] , \regfile/reg_out[22][21] ,
         \regfile/reg_out[22][22] , \regfile/reg_out[22][23] ,
         \regfile/reg_out[22][24] , \regfile/reg_out[22][25] ,
         \regfile/reg_out[22][26] , \regfile/reg_out[22][27] ,
         \regfile/reg_out[22][28] , \regfile/reg_out[22][29] ,
         \regfile/reg_out[22][30] , \regfile/reg_out[22][31] ,
         \regfile/reg_out[23][0] , \regfile/reg_out[23][1] ,
         \regfile/reg_out[23][2] , \regfile/reg_out[23][3] ,
         \regfile/reg_out[23][4] , \regfile/reg_out[23][5] ,
         \regfile/reg_out[23][6] , \regfile/reg_out[23][7] ,
         \regfile/reg_out[23][8] , \regfile/reg_out[23][9] ,
         \regfile/reg_out[23][10] , \regfile/reg_out[23][11] ,
         \regfile/reg_out[23][12] , \regfile/reg_out[23][13] ,
         \regfile/reg_out[23][14] , \regfile/reg_out[23][15] ,
         \regfile/reg_out[23][16] , \regfile/reg_out[23][17] ,
         \regfile/reg_out[23][18] , \regfile/reg_out[23][19] ,
         \regfile/reg_out[23][20] , \regfile/reg_out[23][21] ,
         \regfile/reg_out[23][22] , \regfile/reg_out[23][23] ,
         \regfile/reg_out[23][24] , \regfile/reg_out[23][25] ,
         \regfile/reg_out[23][26] , \regfile/reg_out[23][27] ,
         \regfile/reg_out[23][28] , \regfile/reg_out[23][29] ,
         \regfile/reg_out[23][30] , \regfile/reg_out[23][31] ,
         \regfile/reg_out[24][0] , \regfile/reg_out[24][1] ,
         \regfile/reg_out[24][2] , \regfile/reg_out[24][3] ,
         \regfile/reg_out[24][4] , \regfile/reg_out[24][5] ,
         \regfile/reg_out[24][6] , \regfile/reg_out[24][7] ,
         \regfile/reg_out[24][8] , \regfile/reg_out[24][9] ,
         \regfile/reg_out[24][10] , \regfile/reg_out[24][11] ,
         \regfile/reg_out[24][12] , \regfile/reg_out[24][13] ,
         \regfile/reg_out[24][14] , \regfile/reg_out[24][15] ,
         \regfile/reg_out[24][16] , \regfile/reg_out[24][17] ,
         \regfile/reg_out[24][18] , \regfile/reg_out[24][19] ,
         \regfile/reg_out[24][20] , \regfile/reg_out[24][21] ,
         \regfile/reg_out[24][22] , \regfile/reg_out[24][23] ,
         \regfile/reg_out[24][24] , \regfile/reg_out[24][25] ,
         \regfile/reg_out[24][26] , \regfile/reg_out[24][27] ,
         \regfile/reg_out[24][28] , \regfile/reg_out[24][29] ,
         \regfile/reg_out[24][30] , \regfile/reg_out[24][31] ,
         \regfile/reg_out[25][0] , \regfile/reg_out[25][1] ,
         \regfile/reg_out[25][2] , \regfile/reg_out[25][3] ,
         \regfile/reg_out[25][4] , \regfile/reg_out[25][5] ,
         \regfile/reg_out[25][6] , \regfile/reg_out[25][7] ,
         \regfile/reg_out[25][8] , \regfile/reg_out[25][9] ,
         \regfile/reg_out[25][10] , \regfile/reg_out[25][11] ,
         \regfile/reg_out[25][12] , \regfile/reg_out[25][13] ,
         \regfile/reg_out[25][14] , \regfile/reg_out[25][15] ,
         \regfile/reg_out[25][16] , \regfile/reg_out[25][17] ,
         \regfile/reg_out[25][18] , \regfile/reg_out[25][19] ,
         \regfile/reg_out[25][20] , \regfile/reg_out[25][21] ,
         \regfile/reg_out[25][22] , \regfile/reg_out[25][23] ,
         \regfile/reg_out[25][24] , \regfile/reg_out[25][25] ,
         \regfile/reg_out[25][26] , \regfile/reg_out[25][27] ,
         \regfile/reg_out[25][28] , \regfile/reg_out[25][29] ,
         \regfile/reg_out[25][30] , \regfile/reg_out[25][31] ,
         \regfile/reg_out[26][0] , \regfile/reg_out[26][1] ,
         \regfile/reg_out[26][2] , \regfile/reg_out[26][3] ,
         \regfile/reg_out[26][4] , \regfile/reg_out[26][5] ,
         \regfile/reg_out[26][6] , \regfile/reg_out[26][7] ,
         \regfile/reg_out[26][8] , \regfile/reg_out[26][9] ,
         \regfile/reg_out[26][10] , \regfile/reg_out[26][11] ,
         \regfile/reg_out[26][12] , \regfile/reg_out[26][13] ,
         \regfile/reg_out[26][14] , \regfile/reg_out[26][15] ,
         \regfile/reg_out[26][16] , \regfile/reg_out[26][17] ,
         \regfile/reg_out[26][18] , \regfile/reg_out[26][19] ,
         \regfile/reg_out[26][20] , \regfile/reg_out[26][21] ,
         \regfile/reg_out[26][22] , \regfile/reg_out[26][23] ,
         \regfile/reg_out[26][24] , \regfile/reg_out[26][25] ,
         \regfile/reg_out[26][26] , \regfile/reg_out[26][27] ,
         \regfile/reg_out[26][28] , \regfile/reg_out[26][29] ,
         \regfile/reg_out[26][30] , \regfile/reg_out[26][31] ,
         \regfile/reg_out[27][0] , \regfile/reg_out[27][1] ,
         \regfile/reg_out[27][2] , \regfile/reg_out[27][3] ,
         \regfile/reg_out[27][4] , \regfile/reg_out[27][5] ,
         \regfile/reg_out[27][6] , \regfile/reg_out[27][7] ,
         \regfile/reg_out[27][8] , \regfile/reg_out[27][9] ,
         \regfile/reg_out[27][10] , \regfile/reg_out[27][11] ,
         \regfile/reg_out[27][12] , \regfile/reg_out[27][13] ,
         \regfile/reg_out[27][14] , \regfile/reg_out[27][15] ,
         \regfile/reg_out[27][16] , \regfile/reg_out[27][17] ,
         \regfile/reg_out[27][18] , \regfile/reg_out[27][19] ,
         \regfile/reg_out[27][20] , \regfile/reg_out[27][21] ,
         \regfile/reg_out[27][22] , \regfile/reg_out[27][23] ,
         \regfile/reg_out[27][24] , \regfile/reg_out[27][25] ,
         \regfile/reg_out[27][26] , \regfile/reg_out[27][27] ,
         \regfile/reg_out[27][28] , \regfile/reg_out[27][29] ,
         \regfile/reg_out[27][30] , \regfile/reg_out[27][31] ,
         \regfile/reg_out[28][0] , \regfile/reg_out[28][1] ,
         \regfile/reg_out[28][2] , \regfile/reg_out[28][3] ,
         \regfile/reg_out[28][4] , \regfile/reg_out[28][5] ,
         \regfile/reg_out[28][6] , \regfile/reg_out[28][7] ,
         \regfile/reg_out[28][8] , \regfile/reg_out[28][9] ,
         \regfile/reg_out[28][10] , \regfile/reg_out[28][11] ,
         \regfile/reg_out[28][12] , \regfile/reg_out[28][13] ,
         \regfile/reg_out[28][14] , \regfile/reg_out[28][15] ,
         \regfile/reg_out[28][16] , \regfile/reg_out[28][17] ,
         \regfile/reg_out[28][18] , \regfile/reg_out[28][19] ,
         \regfile/reg_out[28][20] , \regfile/reg_out[28][21] ,
         \regfile/reg_out[28][22] , \regfile/reg_out[28][23] ,
         \regfile/reg_out[28][24] , \regfile/reg_out[28][25] ,
         \regfile/reg_out[28][26] , \regfile/reg_out[28][27] ,
         \regfile/reg_out[28][28] , \regfile/reg_out[28][29] ,
         \regfile/reg_out[28][30] , \regfile/reg_out[28][31] ,
         \regfile/reg_out[29][0] , \regfile/reg_out[29][1] ,
         \regfile/reg_out[29][2] , \regfile/reg_out[29][3] ,
         \regfile/reg_out[29][4] , \regfile/reg_out[29][5] ,
         \regfile/reg_out[29][6] , \regfile/reg_out[29][7] ,
         \regfile/reg_out[29][8] , \regfile/reg_out[29][9] ,
         \regfile/reg_out[29][10] , \regfile/reg_out[29][11] ,
         \regfile/reg_out[29][12] , \regfile/reg_out[29][13] ,
         \regfile/reg_out[29][14] , \regfile/reg_out[29][15] ,
         \regfile/reg_out[29][16] , \regfile/reg_out[29][17] ,
         \regfile/reg_out[29][18] , \regfile/reg_out[29][19] ,
         \regfile/reg_out[29][20] , \regfile/reg_out[29][21] ,
         \regfile/reg_out[29][22] , \regfile/reg_out[29][23] ,
         \regfile/reg_out[29][24] , \regfile/reg_out[29][25] ,
         \regfile/reg_out[29][26] , \regfile/reg_out[29][27] ,
         \regfile/reg_out[29][28] , \regfile/reg_out[29][29] ,
         \regfile/reg_out[29][30] , \regfile/reg_out[29][31] ,
         \regfile/reg_out[30][0] , \regfile/reg_out[30][1] ,
         \regfile/reg_out[30][2] , \regfile/reg_out[30][3] ,
         \regfile/reg_out[30][4] , \regfile/reg_out[30][5] ,
         \regfile/reg_out[30][6] , \regfile/reg_out[30][7] ,
         \regfile/reg_out[30][8] , \regfile/reg_out[30][9] ,
         \regfile/reg_out[30][10] , \regfile/reg_out[30][11] ,
         \regfile/reg_out[30][12] , \regfile/reg_out[30][13] ,
         \regfile/reg_out[30][14] , \regfile/reg_out[30][15] ,
         \regfile/reg_out[30][16] , \regfile/reg_out[30][17] ,
         \regfile/reg_out[30][18] , \regfile/reg_out[30][19] ,
         \regfile/reg_out[30][20] , \regfile/reg_out[30][21] ,
         \regfile/reg_out[30][22] , \regfile/reg_out[30][23] ,
         \regfile/reg_out[30][24] , \regfile/reg_out[30][25] ,
         \regfile/reg_out[30][26] , \regfile/reg_out[30][27] ,
         \regfile/reg_out[30][28] , \regfile/reg_out[30][29] ,
         \regfile/reg_out[30][30] , \regfile/reg_out[30][31] ,
         \regfile/reg_out[31][0] , \regfile/reg_out[31][1] ,
         \regfile/reg_out[31][2] , \regfile/reg_out[31][3] ,
         \regfile/reg_out[31][4] , \regfile/reg_out[31][5] ,
         \regfile/reg_out[31][6] , \regfile/reg_out[31][7] ,
         \regfile/reg_out[31][8] , \regfile/reg_out[31][9] ,
         \regfile/reg_out[31][10] , \regfile/reg_out[31][11] ,
         \regfile/reg_out[31][12] , \regfile/reg_out[31][13] ,
         \regfile/reg_out[31][14] , \regfile/reg_out[31][15] ,
         \regfile/reg_out[31][16] , \regfile/reg_out[31][17] ,
         \regfile/reg_out[31][18] , \regfile/reg_out[31][19] ,
         \regfile/reg_out[31][20] , \regfile/reg_out[31][21] ,
         \regfile/reg_out[31][22] , \regfile/reg_out[31][23] ,
         \regfile/reg_out[31][24] , \regfile/reg_out[31][25] ,
         \regfile/reg_out[31][26] , \regfile/reg_out[31][27] ,
         \regfile/reg_out[31][28] , \regfile/reg_out[31][29] ,
         \regfile/reg_out[31][30] , \regfile/reg_out[31][31] ,
         \regfile/reg_out[1][0] , \regfile/reg_out[1][1] ,
         \regfile/reg_out[1][2] , \regfile/reg_out[1][3] ,
         \regfile/reg_out[1][4] , \regfile/reg_out[1][5] ,
         \regfile/reg_out[1][6] , \regfile/reg_out[1][7] ,
         \regfile/reg_out[1][8] , \regfile/reg_out[1][9] ,
         \regfile/reg_out[1][10] , \regfile/reg_out[1][11] ,
         \regfile/reg_out[1][12] , \regfile/reg_out[1][13] ,
         \regfile/reg_out[1][14] , \regfile/reg_out[1][15] ,
         \regfile/reg_out[1][16] , \regfile/reg_out[1][17] ,
         \regfile/reg_out[1][18] , \regfile/reg_out[1][19] ,
         \regfile/reg_out[1][20] , \regfile/reg_out[1][21] ,
         \regfile/reg_out[1][22] , \regfile/reg_out[1][23] ,
         \regfile/reg_out[1][24] , \regfile/reg_out[1][25] ,
         \regfile/reg_out[1][26] , \regfile/reg_out[1][27] ,
         \regfile/reg_out[1][28] , \regfile/reg_out[1][29] ,
         \regfile/reg_out[1][30] , \regfile/reg_out[1][31] ,
         \regfile/reg_out[2][0] , \regfile/reg_out[2][1] ,
         \regfile/reg_out[2][2] , \regfile/reg_out[2][3] ,
         \regfile/reg_out[2][4] , \regfile/reg_out[2][5] ,
         \regfile/reg_out[2][6] , \regfile/reg_out[2][7] ,
         \regfile/reg_out[2][8] , \regfile/reg_out[2][9] ,
         \regfile/reg_out[2][10] , \regfile/reg_out[2][11] ,
         \regfile/reg_out[2][12] , \regfile/reg_out[2][13] ,
         \regfile/reg_out[2][14] , \regfile/reg_out[2][15] ,
         \regfile/reg_out[2][16] , \regfile/reg_out[2][17] ,
         \regfile/reg_out[2][18] , \regfile/reg_out[2][19] ,
         \regfile/reg_out[2][20] , \regfile/reg_out[2][21] ,
         \regfile/reg_out[2][22] , \regfile/reg_out[2][23] ,
         \regfile/reg_out[2][24] , \regfile/reg_out[2][25] ,
         \regfile/reg_out[2][26] , \regfile/reg_out[2][27] ,
         \regfile/reg_out[2][28] , \regfile/reg_out[2][29] ,
         \regfile/reg_out[2][30] , \regfile/reg_out[2][31] ,
         \regfile/reg_out[3][0] , \regfile/reg_out[3][1] ,
         \regfile/reg_out[3][2] , \regfile/reg_out[3][3] ,
         \regfile/reg_out[3][4] , \regfile/reg_out[3][5] ,
         \regfile/reg_out[3][6] , \regfile/reg_out[3][7] ,
         \regfile/reg_out[3][8] , \regfile/reg_out[3][9] ,
         \regfile/reg_out[3][10] , \regfile/reg_out[3][11] ,
         \regfile/reg_out[3][12] , \regfile/reg_out[3][13] ,
         \regfile/reg_out[3][14] , \regfile/reg_out[3][15] ,
         \regfile/reg_out[3][16] , \regfile/reg_out[3][17] ,
         \regfile/reg_out[3][18] , \regfile/reg_out[3][19] ,
         \regfile/reg_out[3][20] , \regfile/reg_out[3][21] ,
         \regfile/reg_out[3][22] , \regfile/reg_out[3][23] ,
         \regfile/reg_out[3][24] , \regfile/reg_out[3][25] ,
         \regfile/reg_out[3][26] , \regfile/reg_out[3][27] ,
         \regfile/reg_out[3][28] , \regfile/reg_out[3][29] ,
         \regfile/reg_out[3][30] , \regfile/reg_out[3][31] ,
         \regfile/reg_out[4][0] , \regfile/reg_out[4][1] ,
         \regfile/reg_out[4][2] , \regfile/reg_out[4][3] ,
         \regfile/reg_out[4][4] , \regfile/reg_out[4][5] ,
         \regfile/reg_out[4][6] , \regfile/reg_out[4][7] ,
         \regfile/reg_out[4][8] , \regfile/reg_out[4][9] ,
         \regfile/reg_out[4][10] , \regfile/reg_out[4][11] ,
         \regfile/reg_out[4][12] , \regfile/reg_out[4][13] ,
         \regfile/reg_out[4][14] , \regfile/reg_out[4][15] ,
         \regfile/reg_out[4][16] , \regfile/reg_out[4][17] ,
         \regfile/reg_out[4][18] , \regfile/reg_out[4][19] ,
         \regfile/reg_out[4][20] , \regfile/reg_out[4][21] ,
         \regfile/reg_out[4][22] , \regfile/reg_out[4][23] ,
         \regfile/reg_out[4][24] , \regfile/reg_out[4][25] ,
         \regfile/reg_out[4][26] , \regfile/reg_out[4][27] ,
         \regfile/reg_out[4][28] , \regfile/reg_out[4][29] ,
         \regfile/reg_out[4][30] , \regfile/reg_out[4][31] ,
         \regfile/reg_out[5][0] , \regfile/reg_out[5][1] ,
         \regfile/reg_out[5][2] , \regfile/reg_out[5][3] ,
         \regfile/reg_out[5][4] , \regfile/reg_out[5][5] ,
         \regfile/reg_out[5][6] , \regfile/reg_out[5][7] ,
         \regfile/reg_out[5][8] , \regfile/reg_out[5][9] ,
         \regfile/reg_out[5][10] , \regfile/reg_out[5][11] ,
         \regfile/reg_out[5][12] , \regfile/reg_out[5][13] ,
         \regfile/reg_out[5][14] , \regfile/reg_out[5][15] ,
         \regfile/reg_out[5][16] , \regfile/reg_out[5][17] ,
         \regfile/reg_out[5][18] , \regfile/reg_out[5][19] ,
         \regfile/reg_out[5][20] , \regfile/reg_out[5][21] ,
         \regfile/reg_out[5][22] , \regfile/reg_out[5][23] ,
         \regfile/reg_out[5][24] , \regfile/reg_out[5][25] ,
         \regfile/reg_out[5][26] , \regfile/reg_out[5][27] ,
         \regfile/reg_out[5][28] , \regfile/reg_out[5][29] ,
         \regfile/reg_out[5][30] , \regfile/reg_out[5][31] ,
         \regfile/reg_out[9][0] , \regfile/reg_out[9][1] ,
         \regfile/reg_out[9][2] , \regfile/reg_out[9][3] ,
         \regfile/reg_out[9][4] , \regfile/reg_out[9][5] ,
         \regfile/reg_out[9][6] , \regfile/reg_out[9][7] ,
         \regfile/reg_out[9][8] , \regfile/reg_out[9][9] ,
         \regfile/reg_out[9][10] , \regfile/reg_out[9][11] ,
         \regfile/reg_out[9][12] , \regfile/reg_out[9][13] ,
         \regfile/reg_out[9][14] , \regfile/reg_out[9][15] ,
         \regfile/reg_out[9][16] , \regfile/reg_out[9][17] ,
         \regfile/reg_out[9][18] , \regfile/reg_out[9][19] ,
         \regfile/reg_out[9][20] , \regfile/reg_out[9][21] ,
         \regfile/reg_out[9][22] , \regfile/reg_out[9][23] ,
         \regfile/reg_out[9][24] , \regfile/reg_out[9][25] ,
         \regfile/reg_out[9][26] , \regfile/reg_out[9][27] ,
         \regfile/reg_out[9][28] , \regfile/reg_out[9][29] ,
         \regfile/reg_out[9][30] , \regfile/reg_out[9][31] ,
         \regfile/reg_out[12][0] , \regfile/reg_out[12][1] ,
         \regfile/reg_out[12][2] , \regfile/reg_out[12][3] ,
         \regfile/reg_out[12][4] , \regfile/reg_out[12][5] ,
         \regfile/reg_out[12][6] , \regfile/reg_out[12][7] ,
         \regfile/reg_out[12][8] , \regfile/reg_out[12][9] ,
         \regfile/reg_out[12][10] , \regfile/reg_out[12][11] ,
         \regfile/reg_out[12][12] , \regfile/reg_out[12][13] ,
         \regfile/reg_out[12][14] , \regfile/reg_out[12][15] ,
         \regfile/reg_out[12][16] , \regfile/reg_out[12][17] ,
         \regfile/reg_out[12][18] , \regfile/reg_out[12][19] ,
         \regfile/reg_out[12][20] , \regfile/reg_out[12][21] ,
         \regfile/reg_out[12][22] , \regfile/reg_out[12][23] ,
         \regfile/reg_out[12][24] , \regfile/reg_out[12][25] ,
         \regfile/reg_out[12][26] , \regfile/reg_out[12][27] ,
         \regfile/reg_out[12][28] , \regfile/reg_out[12][29] ,
         \regfile/reg_out[12][30] , \regfile/reg_out[12][31] ,
         \regfile/reg_out[13][0] , \regfile/reg_out[13][1] ,
         \regfile/reg_out[13][2] , \regfile/reg_out[13][3] ,
         \regfile/reg_out[13][4] , \regfile/reg_out[13][5] ,
         \regfile/reg_out[13][6] , \regfile/reg_out[13][7] ,
         \regfile/reg_out[13][8] , \regfile/reg_out[13][9] ,
         \regfile/reg_out[13][10] , \regfile/reg_out[13][11] ,
         \regfile/reg_out[13][12] , \regfile/reg_out[13][13] ,
         \regfile/reg_out[13][14] , \regfile/reg_out[13][15] ,
         \regfile/reg_out[13][16] , \regfile/reg_out[13][17] ,
         \regfile/reg_out[13][18] , \regfile/reg_out[13][19] ,
         \regfile/reg_out[13][20] , \regfile/reg_out[13][21] ,
         \regfile/reg_out[13][22] , \regfile/reg_out[13][23] ,
         \regfile/reg_out[13][24] , \regfile/reg_out[13][25] ,
         \regfile/reg_out[13][26] , \regfile/reg_out[13][27] ,
         \regfile/reg_out[13][28] , \regfile/reg_out[13][29] ,
         \regfile/reg_out[13][30] , \regfile/reg_out[13][31] ,
         \BYP_BRANCH_MUXB/N39 , \BYP_BRANCH_MUXB/N4 , \Mcontrol/N34 ,
         \Mcontrol/N25 , \Mcontrol/N17 ,
         \Mcontrol/x_sampled_dmem_command[SIGN] ,
         \Mcontrol/x_sampled_dmem_command[MW] , \Mcontrol/x_sampled_dwe ,
         \Mcontrol/m_sampled_xrd[0] , \Mcontrol/m_sampled_xrd[1] ,
         \Mcontrol/m_sampled_xrd[2] , \Mcontrol/m_sampled_xrd[3] ,
         \Mcontrol/m_sampled_xrd[4] , \Mcontrol/x_rd[0] , \Mcontrol/x_rd[1] ,
         \Mcontrol/x_rd[2] , \Mcontrol/x_rd[3] , \Mcontrol/x_rd[4] ,
         \Mcontrol/d_jump_type[0] , \Mcontrol/d_jump_type[1] ,
         \Mcontrol/d_jump_type[2] , \Mcontrol/d_jump_type[3] ,
         \Mcontrol/f_currpc[0] , \Mcontrol/f_currpc[1] ,
         \Mcontrol/f_currpc[2] , \Mcontrol/f_currpc[3] ,
         \Mcontrol/f_currpc[4] , \Mcontrol/f_currpc[5] ,
         \Mcontrol/f_currpc[6] , \Mcontrol/f_currpc[7] ,
         \Mcontrol/f_currpc[8] , \Mcontrol/f_currpc[9] ,
         \Mcontrol/f_currpc[10] , \Mcontrol/f_currpc[11] ,
         \Mcontrol/f_currpc[12] , \Mcontrol/f_currpc[13] ,
         \Mcontrol/f_currpc[14] , \Mcontrol/f_currpc[15] ,
         \Mcontrol/f_currpc[16] , \Mcontrol/f_currpc[17] ,
         \Mcontrol/f_currpc[18] , \Mcontrol/f_currpc[19] ,
         \Mcontrol/f_currpc[20] , \Mcontrol/f_currpc[21] ,
         \Mcontrol/f_currpc[22] , \Mcontrol/f_currpc[23] ,
         \Mcontrol/stall_decode , \Mcontrol/int_reset , \Mcontrol/bvgen/N9 ,
         \Mcontrol/bvgen/N8 , \Mcontrol/bvgen/N7 , \Mcontrol/bvgen/N6 ,
         \Mcontrol/bvgen/N4 , \Mcontrol/bvgen/N3 , \Mcontrol/bvgen/N2 ,
         \Mcontrol/bvgen/x_jump_type[0] , \Mcontrol/bvgen/d_curr_pc[0] ,
         \Mcontrol/bvgen/d_curr_pc[1] , \Mcontrol/bvgen/d_curr_pc[2] ,
         \Mcontrol/bvgen/d_curr_pc[3] , \Mcontrol/bvgen/d_curr_pc[4] ,
         \Mcontrol/bvgen/d_curr_pc[5] , \Mcontrol/bvgen/d_curr_pc[6] ,
         \Mcontrol/bvgen/d_curr_pc[7] , \Mcontrol/bvgen/d_curr_pc[8] ,
         \Mcontrol/bvgen/d_curr_pc[9] , \Mcontrol/bvgen/d_curr_pc[10] ,
         \Mcontrol/bvgen/d_curr_pc[11] , \Mcontrol/bvgen/d_curr_pc[12] ,
         \Mcontrol/bvgen/d_curr_pc[13] , \Mcontrol/bvgen/d_curr_pc[14] ,
         \Mcontrol/bvgen/d_curr_pc[15] , \Mcontrol/bvgen/d_curr_pc[16] ,
         \Mcontrol/bvgen/d_curr_pc[17] , \Mcontrol/bvgen/d_curr_pc[18] ,
         \Mcontrol/bvgen/d_curr_pc[19] , \Mcontrol/bvgen/d_curr_pc[20] ,
         \Mcontrol/bvgen/d_curr_pc[21] , \Mcontrol/bvgen/d_curr_pc[22] ,
         \Mcontrol/bvgen/d_curr_pc[23] , \Mcontrol/Operation_decoding32/N2087 ,
         \Mcontrol/Operation_decoding32/N2084 ,
         \Mcontrol/Operation_decoding32/N2071 ,
         \Mcontrol/Operation_decoding32/N2070 ,
         \Mcontrol/Operation_decoding32/N2066 ,
         \Mcontrol/Operation_decoding32/N2064 ,
         \Mcontrol/Operation_decoding32/N2062 ,
         \Mcontrol/Operation_decoding32/N2060 ,
         \Mcontrol/Operation_decoding32/N2056 ,
         \Mcontrol/Operation_decoding32/N2054 ,
         \Mcontrol/Operation_decoding32/N2047 ,
         \Mcontrol/Operation_decoding32/N2046 ,
         \Mcontrol/Operation_decoding32/N2045 ,
         \Mcontrol/Operation_decoding32/N2041 ,
         \Mcontrol/Operation_decoding32/N2037 ,
         \Mcontrol/Operation_decoding32/N2036 ,
         \Mcontrol/Operation_decoding32/N2035 ,
         \Mcontrol/Operation_decoding32/N2030 ,
         \Mcontrol/Operation_decoding32/N2029 ,
         \Mcontrol/Operation_decoding32/N2021 ,
         \Mcontrol/Operation_decoding32/N2017 ,
         \Mcontrol/Operation_decoding32/N2007 ,
         \Mcontrol/Operation_decoding32/N2005 ,
         \Mcontrol/Operation_decoding32/N2003 ,
         \Mcontrol/Operation_decoding32/N2001 ,
         \Mcontrol/Operation_decoding32/N1996 ,
         \Mcontrol/Operation_decoding32/N1990 ,
         \Mcontrol/Operation_decoding32/N1989 ,
         \Mcontrol/Operation_decoding32/N1987 ,
         \Mcontrol/Operation_decoding32/N1984 ,
         \Mcontrol/Operation_decoding32/N1982 ,
         \Mcontrol/Operation_decoding32/N1976 ,
         \Mcontrol/Operation_decoding32/N1975 ,
         \Mcontrol/Operation_decoding32/N1970 ,
         \Mcontrol/Operation_decoding32/N1969 ,
         \Mcontrol/Operation_decoding32/N1968 ,
         \Mcontrol/Operation_decoding32/N1964 ,
         \Mcontrol/Operation_decoding32/N1963 ,
         \Mcontrol/Operation_decoding32/N1958 ,
         \Mcontrol/Operation_decoding32/N1957 ,
         \Mcontrol/Operation_decoding32/N1955 ,
         \Mcontrol/Operation_decoding32/N1952 ,
         \Mcontrol/Operation_decoding32/N1951 ,
         \Mcontrol/Operation_decoding32/N1944 ,
         \Mcontrol/Operation_decoding32/N1939 ,
         \Mcontrol/Operation_decoding32/N1933 ,
         \Mcontrol/Operation_decoding32/N1928 ,
         \Mcontrol/Operation_decoding32/N1924 ,
         \Mcontrol/Operation_decoding32/N1923 ,
         \Mcontrol/Operation_decoding32/N1922 ,
         \Mcontrol/Operation_decoding32/N1921 ,
         \Mcontrol/Operation_decoding32/N1917 ,
         \Mcontrol/Operation_decoding32/N1916 ,
         \Mcontrol/Operation_decoding32/N1915 ,
         \Mcontrol/Operation_decoding32/N1914 ,
         \Mcontrol/Operation_decoding32/N1913 ,
         \Mcontrol/Operation_decoding32/N1912 ,
         \Mcontrol/Operation_decoding32/N1911 ,
         \Mcontrol/Operation_decoding32/N1910 ,
         \Mcontrol/Operation_decoding32/N1909 ,
         \Mcontrol/Operation_decoding32/N1908 ,
         \Mcontrol/Operation_decoding32/N1907 ,
         \Mcontrol/Operation_decoding32/N1906 ,
         \Mcontrol/Operation_decoding32/N1905 ,
         \Mcontrol/Operation_decoding32/N1904 ,
         \Mcontrol/Operation_decoding32/N1903 ,
         \Mcontrol/Operation_decoding32/N1902 ,
         \Mcontrol/Operation_decoding32/N1900 ,
         \Mcontrol/Operation_decoding32/N1899 ,
         \Mcontrol/Operation_decoding32/N1898 ,
         \Mcontrol/Operation_decoding32/N1897 ,
         \Mcontrol/Operation_decoding32/N1896 ,
         \Mcontrol/Operation_decoding32/N1895 ,
         \Mcontrol/Operation_decoding32/N1894 ,
         \Mcontrol/Operation_decoding32/N1893 ,
         \Mcontrol/Operation_decoding32/N1892 ,
         \Mcontrol/Operation_decoding32/N1891 ,
         \Mcontrol/Operation_decoding32/N1890 ,
         \Mcontrol/Operation_decoding32/N1889 ,
         \Mcontrol/Operation_decoding32/N1887 ,
         \Mcontrol/Operation_decoding32/N1886 ,
         \Mcontrol/Operation_decoding32/N1885 ,
         \Mcontrol/Operation_decoding32/N1884 ,
         \Mcontrol/Operation_decoding32/N1883 ,
         \Mcontrol/Operation_decoding32/N1881 ,
         \Mcontrol/Operation_decoding32/N1880 ,
         \Mcontrol/Operation_decoding32/N1873 ,
         \Mcontrol/Operation_decoding32/N1871 ,
         \Mcontrol/Operation_decoding32/N89 ,
         \Mcontrol/Operation_decoding32/N62 , \Mcontrol/Nextpc_decoding/N325 ,
         \Mcontrol/Nextpc_decoding/N324 , \Mcontrol/Nextpc_decoding/N323 ,
         \Mcontrol/Nextpc_decoding/N322 , \Mcontrol/Nextpc_decoding/N321 ,
         \Mcontrol/Nextpc_decoding/N319 , \Mcontrol/Nextpc_decoding/N318 ,
         \Mcontrol/Nextpc_decoding/N317 , \Mcontrol/Nextpc_decoding/N316 ,
         \Mcontrol/Nextpc_decoding/N315 , \Mcontrol/Nextpc_decoding/N313 ,
         \Mcontrol/Nextpc_decoding/N312 , \Mcontrol/Nextpc_decoding/N311 ,
         \Mcontrol/Nextpc_decoding/N310 , \Mcontrol/Nextpc_decoding/N309 ,
         \Mcontrol/Nextpc_decoding/N307 , \Mcontrol/Nextpc_decoding/N306 ,
         \Mcontrol/Nextpc_decoding/N305 , \Mcontrol/Nextpc_decoding/N304 ,
         \Mcontrol/Nextpc_decoding/N303 , \Mcontrol/Nextpc_decoding/N301 ,
         \Mcontrol/Nextpc_decoding/N300 , \Mcontrol/Nextpc_decoding/N299 ,
         \Mcontrol/Nextpc_decoding/N298 , \Mcontrol/Nextpc_decoding/N297 ,
         \Mcontrol/Nextpc_decoding/N295 , \Mcontrol/Nextpc_decoding/N294 ,
         \Mcontrol/Nextpc_decoding/N293 , \Mcontrol/Nextpc_decoding/N292 ,
         \Mcontrol/Nextpc_decoding/N291 , \Mcontrol/Nextpc_decoding/N289 ,
         \Mcontrol/Nextpc_decoding/N288 , \Mcontrol/Nextpc_decoding/N287 ,
         \Mcontrol/Nextpc_decoding/N286 , \Mcontrol/Nextpc_decoding/N285 ,
         \Mcontrol/Nextpc_decoding/N283 , \Mcontrol/Nextpc_decoding/N253 ,
         \Mcontrol/Nextpc_decoding/N252 , \Mcontrol/Nextpc_decoding/N249 ,
         \Mcontrol/Nextpc_decoding/N221 , \Mcontrol/Nextpc_decoding/N219 ,
         \Mcontrol/Nextpc_decoding/N198 , \Mcontrol/Nextpc_decoding/N188 ,
         \Mcontrol/Nextpc_decoding/N182 , \Mcontrol/Nextpc_decoding/N173 ,
         \Mcontrol/Nextpc_decoding/N171 , \Mcontrol/Nextpc_decoding/N170 ,
         \Mcontrol/Nextpc_decoding/N169 , \Mcontrol/Nextpc_decoding/N168 ,
         \Mcontrol/Nextpc_decoding/N36 , \Mcontrol/Nextpc_decoding/N31 ,
         \Mcontrol/Nextpc_decoding/N29 , \Mcontrol/Nextpc_decoding/condition ,
         \Mcontrol/Nextpc_decoding/N26 , \Mcontrol/bp_logicA/N16 ,
         \Mcontrol/bp_logicA/N14 , \Mcontrol/bp_logicA/N13 ,
         \Mcontrol/bp_logicA/N12 , \Mcontrol/bp_logicA/N11 ,
         \Mcontrol/bp_logicA/N10 , \Mcontrol/bp_logicA/N8 ,
         \Mcontrol/bp_logicA/N7 , \Mcontrol/bp_logicA/N6 ,
         \Mcontrol/bp_logicA/N5 , \Mcontrol/bp_logicA/memory_main ,
         \Mcontrol/bp_logicA/N3 , \Mcontrol/bp_logicA/exec_main ,
         \Mcontrol/bp_logicA/N2 , \Mcontrol/bp_logicB/N16 ,
         \Mcontrol/bp_logicB/N15 , \Mcontrol/bp_logicB/N14 ,
         \Mcontrol/bp_logicB/N13 , \Mcontrol/bp_logicB/N12 ,
         \Mcontrol/bp_logicB/N11 , \Mcontrol/bp_logicB/N10 ,
         \Mcontrol/bp_logicB/N9 , \Mcontrol/bp_logicB/N8 ,
         \Mcontrol/bp_logicB/N7 , \Mcontrol/bp_logicB/N6 ,
         \Mcontrol/bp_logicB/N5 , \Mcontrol/bp_logicB/memory_main ,
         \Mcontrol/bp_logicB/N3 , \Mcontrol/bp_logicB/exec_main ,
         \Mcontrol/bp_logicB/N2 , \Mcontrol/st_logic/N120 ,
         \Mcontrol/st_logic/N119 , \Mcontrol/st_logic/N118 ,
         \Mcontrol/st_logic/N117 , \Mcontrol/st_logic/N116 ,
         \Mcontrol/st_logic/N115 , \Mcontrol/st_logic/N114 ,
         \Mcontrol/st_logic/N113 , \Mcontrol/st_logic/N110 ,
         \Mcontrol/st_logic/N109 , \Mcontrol/st_logic/N108 ,
         \Mcontrol/st_logic/N107 , \Mcontrol/st_logic/N106 ,
         \Mcontrol/st_logic/N105 , \Mcontrol/st_logic/N103 ,
         \Mcontrol/st_logic/N102 , \Mcontrol/st_logic/N101 ,
         \Mcontrol/st_logic/N100 , \Mcontrol/st_logic/N99 ,
         \Mcontrol/st_logic/N98 , \Mcontrol/st_logic/N95 ,
         \Mcontrol/st_logic/N94 , \Mcontrol/st_logic/N93 ,
         \Mcontrol/st_logic/N92 , \Mcontrol/st_logic/N90 ,
         \Mcontrol/st_logic/N88 , \Mcontrol/st_logic/N87 ,
         \Mcontrol/st_logic/N86 , \Mcontrol/st_logic/N85 ,
         \Mcontrol/st_logic/N83 , \Mcontrol/st_logic/N82 ,
         \Mcontrol/st_logic/N81 , \Mcontrol/st_logic/N80 ,
         \Mcontrol/st_logic/N79 , \Mcontrol/st_logic/N77 ,
         \Mcontrol/st_logic/N76 , \Mcontrol/st_logic/N75 ,
         \Mcontrol/st_logic/N74 , \Mcontrol/st_logic/N73 ,
         \Mcontrol/st_logic/N71 , \Mcontrol/st_logic/N70 ,
         \Mcontrol/st_logic/N69 , \Mcontrol/st_logic/N68 ,
         \Mcontrol/st_logic/N67 , \Mcontrol/st_logic/N65 ,
         \Mcontrol/st_logic/N64 , \Mcontrol/st_logic/N63 ,
         \Mcontrol/st_logic/N62 , \Mcontrol/st_logic/N61 ,
         \Mcontrol/st_logic/N60 , \Mcontrol/st_logic/N58 ,
         \Mcontrol/st_logic/N57 , \Mcontrol/st_logic/N56 ,
         \Mcontrol/st_logic/N55 , \Mcontrol/st_logic/N54 ,
         \Mcontrol/st_logic/N53 , \Mcontrol/st_logic/N52 ,
         \Mcontrol/st_logic/N51 , \Mcontrol/st_logic/N50 ,
         \Mcontrol/st_logic/N49 , \Mcontrol/st_logic/N47 ,
         \Mcontrol/st_logic/N46 , \Mcontrol/st_logic/N45 ,
         \Mcontrol/st_logic/N44 , \Mcontrol/st_logic/N42 ,
         \Mcontrol/st_logic/N41 , \Mcontrol/st_logic/N40 ,
         \Mcontrol/st_logic/N39 , \Mcontrol/st_logic/N38 ,
         \Mcontrol/st_logic/N37 , \Mcontrol/st_logic/N36 ,
         \Mcontrol/st_logic/N35 , \Mcontrol/st_logic/N34 ,
         \Mcontrol/st_logic/N33 , \Mcontrol/st_logic/N32 ,
         \Mcontrol/st_logic/N31 , \Mcontrol/st_logic/N30 ,
         \Mcontrol/st_logic/N29 , \Mcontrol/st_logic/N28 ,
         \Mcontrol/st_logic/N27 , \Mcontrol/st_logic/N26 ,
         \Mcontrol/st_logic/N25 , \Mcontrol/st_logic/N24 ,
         \Mcontrol/st_logic/N23 , \Mcontrol/st_logic/N22 ,
         \Mcontrol/st_logic/N19 , \Mcontrol/st_logic/N18 ,
         \Mcontrol/st_logic/N15 , \Mcontrol/st_logic/N14 ,
         \Mcontrol/st_logic/N13 , \Mcontrol/st_logic/N12 ,
         \Mcontrol/st_logic/N10 , \Mcontrol/st_logic/branchmul_stall ,
         \Mcontrol/st_logic/N8 ,
         \Mcontrol/st_logic/branch_uses_main_exe_result ,
         \Mcontrol/st_logic/N7 , \Mcontrol/st_logic/branchlw_stall ,
         \Mcontrol/st_logic/N6 ,
         \Mcontrol/st_logic/branch_uses_main_mem_result ,
         \Mcontrol/st_logic/N5 , \Mcontrol/st_logic/branch_uses_regb ,
         \Mcontrol/st_logic/N4 , \Mcontrol/st_logic/branch_uses_rega ,
         \Mcontrol/st_logic/N3 , \Mcontrol/st_logic/load_stall ,
         \Mcontrol/st_logic/N2 , \Mpath/N197 , \Mpath/N196 , \Mpath/N193 ,
         \Mpath/N190 , \Mpath/N189 , \Mpath/N188 , \Mpath/N187 , \Mpath/N186 ,
         \Mpath/N185 , \Mpath/N184 , \Mpath/N183 , \Mpath/N182 , \Mpath/N181 ,
         \Mpath/N180 , \Mpath/N179 , \Mpath/out_jar[0] , \Mpath/out_regB[0] ,
         \Mpath/out_regB[1] , \Mpath/out_regB[2] , \Mpath/out_regB[3] ,
         \Mpath/out_regB[4] , \Mpath/out_regB[5] , \Mpath/out_regB[6] ,
         \Mpath/out_regB[7] , \Mpath/out_regB[8] , \Mpath/out_regB[9] ,
         \Mpath/out_regB[10] , \Mpath/out_regB[11] , \Mpath/out_regB[12] ,
         \Mpath/out_regB[13] , \Mpath/out_regB[14] , \Mpath/out_regB[15] ,
         \Mpath/out_regB[16] , \Mpath/out_regB[17] , \Mpath/out_regB[18] ,
         \Mpath/out_regB[19] , \Mpath/out_regB[20] , \Mpath/out_regB[21] ,
         \Mpath/out_regB[22] , \Mpath/out_regB[23] , \Mpath/out_regB[24] ,
         \Mpath/out_regB[25] , \Mpath/out_regB[26] , \Mpath/out_regB[27] ,
         \Mpath/out_regB[28] , \Mpath/out_regB[29] , \Mpath/out_regB[30] ,
         \Mpath/out_regB[31] , \Mpath/out_regA[0] , \Mpath/out_regA[1] ,
         \Mpath/out_regA[2] , \Mpath/out_regA[3] , \Mpath/out_regA[4] ,
         \Mpath/out_regA[5] , \Mpath/out_regA[6] , \Mpath/out_regA[7] ,
         \Mpath/out_regA[9] , \Mpath/out_regA[10] , \Mpath/out_regA[11] ,
         \Mpath/out_regA[12] , \Mpath/out_regA[13] , \Mpath/out_regA[14] ,
         \Mpath/out_regA[15] , \Mpath/out_regA[16] , \Mpath/out_regA[17] ,
         \Mpath/out_regA[18] , \Mpath/out_regA[19] , \Mpath/out_regA[20] ,
         \Mpath/out_regA[21] , \Mpath/out_regA[22] , \Mpath/out_regA[23] ,
         \Mpath/out_regA[24] , \Mpath/out_regA[25] , \Mpath/out_regA[26] ,
         \Mpath/out_regA[27] , \Mpath/out_regA[28] , \Mpath/out_regA[29] ,
         \Mpath/out_regA[30] , \Mpath/out_regA[31] , \Mpath/the_alu/N526 ,
         \Mpath/the_alu/N525 , \Mpath/the_alu/N524 , \Mpath/the_alu/N523 ,
         \Mpath/the_alu/N520 , \Mpath/the_alu/N519 , \Mpath/the_alu/N518 ,
         \Mpath/the_alu/N517 , \Mpath/the_alu/N515 , \Mpath/the_alu/N514 ,
         \Mpath/the_alu/N513 , \Mpath/the_alu/N512 , \Mpath/the_alu/N511 ,
         \Mpath/the_alu/N509 , \Mpath/the_alu/N508 , \Mpath/the_alu/N507 ,
         \Mpath/the_alu/N506 , \Mpath/the_alu/N505 , \Mpath/the_alu/N503 ,
         \Mpath/the_alu/N502 , \Mpath/the_alu/N501 , \Mpath/the_alu/N500 ,
         \Mpath/the_alu/N499 , \Mpath/the_alu/N498 , \Mpath/the_alu/N497 ,
         \Mpath/the_alu/N496 , \Mpath/the_alu/N495 , \Mpath/the_alu/N494 ,
         \Mpath/the_alu/N493 , \Mpath/the_alu/N492 , \Mpath/the_alu/N491 ,
         \Mpath/the_alu/N490 , \Mpath/the_alu/N489 , \Mpath/the_alu/N488 ,
         \Mpath/the_alu/N487 , \Mpath/the_alu/N486 , \Mpath/the_alu/N485 ,
         \Mpath/the_alu/N484 , \Mpath/the_alu/N483 , \Mpath/the_alu/N482 ,
         \Mpath/the_alu/N481 , \Mpath/the_alu/N480 , \Mpath/the_alu/N479 ,
         \Mpath/the_alu/N478 , \Mpath/the_alu/N477 , \Mpath/the_alu/N476 ,
         \Mpath/the_alu/N475 , \Mpath/the_alu/N474 , \Mpath/the_alu/N473 ,
         \Mpath/the_alu/N472 , \Mpath/the_alu/N471 , \Mpath/the_alu/N470 ,
         \Mpath/the_alu/N469 , \Mpath/the_alu/N468 , \Mpath/the_alu/N467 ,
         \Mpath/the_alu/N466 , \Mpath/the_alu/N465 , \Mpath/the_alu/N464 ,
         \Mpath/the_alu/N463 , \Mpath/the_alu/N462 , \Mpath/the_alu/N461 ,
         \Mpath/the_alu/N460 , \Mpath/the_alu/N457 , \Mpath/the_alu/N456 ,
         \Mpath/the_alu/N455 , \Mpath/the_alu/N454 , \Mpath/the_alu/N453 ,
         \Mpath/the_alu/N448 , \Mpath/the_alu/N221 , \Mpath/the_alu/N219 ,
         \Mpath/the_alu/N218 , \Mpath/the_alu/N217 , \Mpath/the_alu/N216 ,
         \Mpath/the_alu/N215 , \Mpath/the_alu/N214 , \Mpath/the_alu/N213 ,
         \Mpath/the_alu/N212 , \Mpath/the_alu/N211 , \Mpath/the_alu/N210 ,
         \Mpath/the_alu/N209 , \Mpath/the_alu/N208 , \Mpath/the_alu/N207 ,
         \Mpath/the_alu/N206 , \Mpath/the_alu/N205 , \Mpath/the_alu/N204 ,
         \Mpath/the_alu/N203 , \Mpath/the_alu/N202 , \Mpath/the_alu/N201 ,
         \Mpath/the_alu/N200 , \Mpath/the_alu/N199 , \Mpath/the_alu/N198 ,
         \Mpath/the_alu/N189 , \Mpath/the_alu/N187 , \Mpath/the_alu/N186 ,
         \Mpath/the_alu/N185 , \Mpath/the_alu/N184 , \Mpath/the_alu/N183 ,
         \Mpath/the_alu/N182 , \Mpath/the_alu/N181 , \Mpath/the_alu/N180 ,
         \Mpath/the_alu/N179 , \Mpath/the_alu/N178 , \Mpath/the_alu/N177 ,
         \Mpath/the_alu/N176 , \Mpath/the_alu/N175 , \Mpath/the_alu/N174 ,
         \Mpath/the_alu/N173 , \Mpath/the_alu/N172 , \Mpath/the_alu/N171 ,
         \Mpath/the_alu/N170 , \Mpath/the_alu/N169 , \Mpath/the_alu/N168 ,
         \Mpath/the_alu/N167 , \Mpath/the_alu/N166 , \Mpath/the_alu/N157 ,
         \Mpath/the_alu/N155 , \Mpath/the_alu/N154 , \Mpath/the_alu/N153 ,
         \Mpath/the_alu/N152 , \Mpath/the_alu/N151 , \Mpath/the_alu/N150 ,
         \Mpath/the_alu/N149 , \Mpath/the_alu/N148 , \Mpath/the_alu/N147 ,
         \Mpath/the_alu/N146 , \Mpath/the_alu/N145 , \Mpath/the_alu/N144 ,
         \Mpath/the_alu/N143 , \Mpath/the_alu/N142 , \Mpath/the_alu/N141 ,
         \Mpath/the_alu/N140 , \Mpath/the_alu/N139 , \Mpath/the_alu/N138 ,
         \Mpath/the_alu/N137 , \Mpath/the_alu/N136 , \Mpath/the_alu/N135 ,
         \Mpath/the_alu/N134 , \Mpath/the_alu/N125 , \Mpath/the_alu/N123 ,
         \Mpath/the_alu/N122 , \Mpath/the_alu/N121 , \Mpath/the_alu/N120 ,
         \Mpath/the_alu/N119 , \Mpath/the_alu/N118 , \Mpath/the_alu/N117 ,
         \Mpath/the_alu/N116 , \Mpath/the_alu/N115 , \Mpath/the_alu/N114 ,
         \Mpath/the_alu/N113 , \Mpath/the_alu/N112 , \Mpath/the_alu/N111 ,
         \Mpath/the_alu/N110 , \Mpath/the_alu/N109 , \Mpath/the_alu/N108 ,
         \Mpath/the_alu/N107 , \Mpath/the_alu/N106 , \Mpath/the_alu/N105 ,
         \Mpath/the_alu/N104 , \Mpath/the_alu/N103 , \Mpath/the_alu/N102 ,
         \Mpath/the_alu/N93 , \Mpath/the_alu/N91 , \Mpath/the_alu/diff[0] ,
         \Mpath/the_alu/diff[1] , \Mpath/the_alu/diff[2] ,
         \Mpath/the_alu/diff[3] , \Mpath/the_alu/diff[4] ,
         \Mpath/the_alu/diff[5] , \Mpath/the_alu/diff[6] ,
         \Mpath/the_alu/diff[7] , \Mpath/the_alu/diff[8] ,
         \Mpath/the_alu/diff[9] , \Mpath/the_alu/diff[10] ,
         \Mpath/the_alu/diff[11] , \Mpath/the_alu/diff[12] ,
         \Mpath/the_alu/diff[13] , \Mpath/the_alu/diff[14] ,
         \Mpath/the_alu/diff[15] , \Mpath/the_alu/diff[16] ,
         \Mpath/the_alu/diff[17] , \Mpath/the_alu/diff[18] ,
         \Mpath/the_alu/diff[19] , \Mpath/the_alu/diff[20] ,
         \Mpath/the_alu/diff[21] , \Mpath/the_alu/diff[22] ,
         \Mpath/the_alu/diff[23] , \Mpath/the_alu/diff[24] ,
         \Mpath/the_alu/diff[25] , \Mpath/the_alu/diff[26] ,
         \Mpath/the_alu/diff[27] , \Mpath/the_alu/diff[28] ,
         \Mpath/the_alu/diff[29] , \Mpath/the_alu/diff[30] ,
         \Mpath/the_alu/diff[31] , \Mpath/the_alu/sum[0] ,
         \Mpath/the_alu/sum[1] , \Mpath/the_alu/sum[2] ,
         \Mpath/the_alu/sum[3] , \Mpath/the_alu/sum[4] ,
         \Mpath/the_alu/sum[5] , \Mpath/the_alu/sum[6] ,
         \Mpath/the_alu/sum[7] , \Mpath/the_alu/sum[8] ,
         \Mpath/the_alu/sum[9] , \Mpath/the_alu/sum[10] ,
         \Mpath/the_alu/sum[11] , \Mpath/the_alu/sum[12] ,
         \Mpath/the_alu/sum[13] , \Mpath/the_alu/sum[14] ,
         \Mpath/the_alu/sum[15] , \Mpath/the_alu/sum[16] ,
         \Mpath/the_alu/sum[17] , \Mpath/the_alu/sum[18] ,
         \Mpath/the_alu/sum[19] , \Mpath/the_alu/sum[20] ,
         \Mpath/the_alu/sum[21] , \Mpath/the_alu/sum[22] ,
         \Mpath/the_alu/sum[23] , \Mpath/the_alu/sum[24] ,
         \Mpath/the_alu/sum[25] , \Mpath/the_alu/sum[26] ,
         \Mpath/the_alu/sum[27] , \Mpath/the_alu/sum[28] ,
         \Mpath/the_alu/sum[29] , \Mpath/the_alu/sum[30] ,
         \Mpath/the_alu/sum[31] , \Mpath/the_alu/N84 , \Mpath/the_alu/N83 ,
         \Mpath/the_alu/N82 , \Mpath/the_alu/N81 , \Mpath/the_alu/N80 ,
         \Mpath/the_alu/N79 , \Mpath/the_alu/N78 , \Mpath/the_alu/N77 ,
         \Mpath/the_alu/N76 , \Mpath/the_alu/N75 , \Mpath/the_alu/N74 ,
         \Mpath/the_alu/N73 , \Mpath/the_alu/N72 , \Mpath/the_alu/N71 ,
         \Mpath/the_alu/N70 , \Mpath/the_alu/N69 , \Mpath/the_alu/N68 ,
         \Mpath/the_alu/N66 , \Mpath/the_alu/N65 , \Mpath/the_alu/N64 ,
         \Mpath/the_alu/N63 , \Mpath/the_alu/N62 , \Mpath/the_alu/N61 ,
         \Mpath/the_alu/N60 , \Mpath/the_alu/N59 , \Mpath/the_alu/N58 ,
         \Mpath/the_alu/N57 , \Mpath/the_alu/N56 , \Mpath/the_alu/N55 ,
         \Mpath/the_alu/N54 , \Mpath/the_alu/N53 , \Mpath/the_alu/N52 ,
         \Mpath/the_alu/N51 , \Mpath/the_alu/N50 , \Mpath/the_alu/N49 ,
         \Mpath/the_alu/N48 , \Mpath/the_alu/N47 , \Mpath/the_alu/N46 ,
         \Mpath/the_alu/N45 , \Mpath/the_alu/N44 , \Mpath/the_alu/N43 ,
         \Mpath/the_alu/N42 , \Mpath/the_alu/N41 , \Mpath/the_alu/N40 ,
         \Mpath/the_alu/N39 , \Mpath/the_alu/N38 , \Mpath/the_alu/N37 ,
         \Mpath/the_alu/N36 , \Mpath/the_alu/N35 , \Mpath/the_alu/N34 ,
         \Mpath/the_alu/N33 , \Mpath/the_alu/N32 , \Mpath/the_alu/N31 ,
         \Mpath/the_alu/N30 , \Mpath/the_alu/N29 , \Mpath/the_alu/N28 ,
         \Mpath/the_alu/N27 , \Mpath/the_alu/N26 , \Mpath/the_alu/N25 ,
         \Mpath/the_alu/N24 , \Mpath/the_alu/N23 , \Mpath/the_alu/N22 ,
         \Mpath/the_alu/N21 , \Mpath/the_alu/N1 , \Mpath/the_shift/N118 ,
         \Mpath/the_shift/N117 , \Mpath/the_shift/N116 ,
         \Mpath/the_shift/N115 , \Mpath/the_shift/N114 ,
         \Mpath/the_shift/N113 , \Mpath/the_shift/N112 ,
         \Mpath/the_shift/N111 , \Mpath/the_shift/N110 ,
         \Mpath/the_shift/N109 , \Mpath/the_shift/N107 ,
         \Mpath/the_shift/N106 , \Mpath/the_shift/N105 ,
         \Mpath/the_shift/N104 , \Mpath/the_memhandle/N244 ,
         \Mpath/the_memhandle/N243 , \Mpath/the_memhandle/N242 ,
         \Mpath/the_memhandle/N241 , \Mpath/the_memhandle/N240 ,
         \Mpath/the_memhandle/N239 , \Mpath/the_memhandle/N238 ,
         \Mpath/the_memhandle/N236 , \Mpath/the_memhandle/N235 ,
         \Mpath/the_memhandle/N120 , \Mpath/the_memhandle/N86 ,
         \Mpath/the_memhandle/N77 , \Mpath/the_memhandle/N76 ,
         \Mpath/the_memhandle/N74 , \Mpath/the_memhandle/N72 ,
         \Mpath/the_memhandle/N39 , \Mpath/the_memhandle/N38 ,
         \Mpath/the_memhandle/N37 , \Mpath/the_memhandle/N36 ,
         \Mpath/the_memhandle/N34 , \Mpath/the_memhandle/smdr_out[8] ,
         \Mpath/the_memhandle/smdr_out[9] , \Mpath/the_memhandle/smdr_out[10] ,
         \Mpath/the_memhandle/smdr_out[11] ,
         \Mpath/the_memhandle/smdr_out[12] ,
         \Mpath/the_memhandle/smdr_out[13] ,
         \Mpath/the_memhandle/smdr_out[14] ,
         \Mpath/the_memhandle/smdr_out[15] ,
         \Mpath/the_memhandle/smdr_out[16] ,
         \Mpath/the_memhandle/smdr_out[17] ,
         \Mpath/the_memhandle/smdr_out[18] ,
         \Mpath/the_memhandle/smdr_out[19] ,
         \Mpath/the_memhandle/smdr_out[20] ,
         \Mpath/the_memhandle/smdr_out[21] ,
         \Mpath/the_memhandle/smdr_out[22] ,
         \Mpath/the_memhandle/smdr_out[23] ,
         \Mpath/the_memhandle/smdr_out[24] ,
         \Mpath/the_memhandle/smdr_out[25] ,
         \Mpath/the_memhandle/smdr_out[26] ,
         \Mpath/the_memhandle/smdr_out[27] ,
         \Mpath/the_memhandle/smdr_out[28] ,
         \Mpath/the_memhandle/smdr_out[29] ,
         \Mpath/the_memhandle/smdr_out[30] ,
         \Mpath/the_memhandle/smdr_out[31] , \d_chk/N13 , \d_chk/N12 ,
         \d_chk/N11 , \d_chk/N10 , \d_chk/N7 , n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n235, n236, n237, n238, n239,
         n240, n241, n243, n244, n246, n247, n248, n249, n250, n251, n252,
         n253, n255, n256, n257, n258, n259, n260, n261, n262, n263, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n278, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n302, n303, n304, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n317, n318, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1436, n1437, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1512, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1849, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n3028, n3039, n3041, n3043, n3045, n3049, n3051, n3052,
         n3054, n3056, n3072, n3083, n3085, n3086, n3087, n3102, n3103, n3104,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4506, n4507, n4508, n4509, n4510,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6057, n6058, n6059, n6060,
         n6063, n6065, n6066, n6067, n6068, n6069, n6073, n6074, n6075, n6076,
         n6077, n6078, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6196, n6197, n6198, n6199,
         n6200, n6201, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6379,
         n6380, n6381, n6383, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6393, n6394, n6395, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6416, n6417, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, net55918, net55916, net55914, net55912, net55910,
         net55908, net55906, net55904, net55902, net55900, net55898, net55896,
         net55894, net55892, net55890, net55888, net55886, net55884, net55882,
         net55880, net55878, net55876, net55874, net55872, net55870, net55868,
         net55866, net55864, net55862, net55860, net55858, net55856, net55854,
         net55852, net55850, net55848, net55846, net55844, net55842, net55840,
         net55838, net55836, net55834, net55832, net55830, net55828, net55826,
         net55824, net55822, net55921, net56216, net56319, net56316, net56595,
         net56605, net56617, net56668, net56678, net56765, net56784, net56846,
         net56922, net56977, net56982, net56996, net57039, net57038, net57184,
         net57236, net57253, net57255, net57268, net57297, net57313, net57323,
         net57331, net57341, net57346, net57366, net57368, net57379, net57386,
         net57388, net57460, net57465, net57474, net57683, net57730, net57757,
         net57810, net57843, net57942, net57954, net58000, net58101, net58300,
         net58533, net58543, net58542, net58547, net58594, net58625, net58826,
         net59543, net59767, net59757, net59736, net59734, net59732, net59612,
         n6100, n6079, n2462, n2461, n1482, \Mcontrol/d_instr[6] ,
         \Mcontrol/d_instr[0] , \Mcontrol/Operation_decoding32/N1901 , n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6890, n6891, n6892, n6893, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7284,
         n7285, n7286, n7287, n7288, n7289, n7291, n7292, n7293, n7294, n7295,
         n7296, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870;
  wire   [7:0] serve_proc_addr;
  wire   [31:0] daddr_out;
  wire   [31:0] break_code;
  wire   [23:0] epc;
  wire   [4:0] rs1_addr;
  wire   [4:0] rs2_addr;
  wire   [4:0] rd_addr;
  wire   [2:0] byp_controlA;
  wire   [2:0] byp_controlB;
  wire   [31:0] branch_rega;
  wire   [31:0] branch_regb;
  wire   [23:0] jar_in;
  wire   [2:0] shift_op;
  wire   [2:0] exe_outsel;
  wire   [5:0] \Scc_coproc/mem_cop_op ;
  wire   [5:0] \Mcontrol/x_mul_command ;
  wire   [31:0] \Mcontrol/d_instr ;
  wire   [31:0] \Mcontrol/d_sampled_finstr ;
  wire   [23:0] \Mcontrol/bvgen/x_curr_pc ;
  wire   [23:0] \Mcontrol/Nextpc_decoding/Bta ;
  wire   [1:0] \Mpath/mem_baddr ;
  wire   [31:0] \Mpath/the_shift/sh_sll ;
  wire   [31:0] \Mpath/the_shift/sh_srl ;
  wire   [31:0] \Mpath/the_shift/sh_sra ;
  wire   [31:0] \Mpath/the_shift/sh_ror ;
  wire   [31:0] \Mpath/the_shift/sh_rol ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign real_dbg_op = 1'b0;
  assign end_dbg = 1'b0;
  assign I_ADDR_OUTBUS[0] = 1'b0;
  assign I_ADDR_OUTBUS[1] = 1'b0;
  assign suspend = 1'b1;
  assign I_ADDR_OUTBUS[23] = net56216;
  assign I_ADDR_OUTBUS[22] = net57039;

  INV_X2 \d_chk/I_0  ( .A(\x_mem_command[MB] ), .ZN(\d_chk/N10 ) );
  INV_X2 \d_chk/I_1  ( .A(\x_mem_command[MH] ), .ZN(\d_chk/N11 ) );
  INV_X2 \d_chk/I_4  ( .A(dcheck_enable), .ZN(\d_chk/N13 ) );
  AND2_X2 \Mpath/the_memhandle/C342  ( .A1(\Mpath/the_memhandle/N235 ), .A2(
        \Mpath/the_memhandle/N236 ), .ZN(\Mpath/the_memhandle/N34 ) );
  AND2_X2 \Mpath/the_memhandle/C344  ( .A1(\Mpath/the_memhandle/N239 ), .A2(
        \Mpath/the_memhandle/N240 ), .ZN(\Mpath/the_memhandle/N36 ) );
  INV_X2 \Mpath/the_memhandle/I_8  ( .A(\Mpath/the_memhandle/N241 ), .ZN(
        \Mpath/the_memhandle/N37 ) );
  OR2_X2 \Mpath/the_memhandle/C348  ( .A1(\Mpath/mem_baddr [1]), .A2(
        \Mpath/the_memhandle/N240 ), .ZN(\Mpath/the_memhandle/N241 ) );
  INV_X2 \Mpath/the_memhandle/I_9  ( .A(\Mpath/the_memhandle/N242 ), .ZN(
        \Mpath/the_memhandle/N38 ) );
  OR2_X2 \Mpath/the_memhandle/C351  ( .A1(\Mpath/the_memhandle/N239 ), .A2(
        \Mpath/mem_baddr [0]), .ZN(\Mpath/the_memhandle/N242 ) );
  AND2_X2 \Mpath/the_memhandle/C353  ( .A1(\Mpath/mem_baddr [1]), .A2(
        \Mpath/mem_baddr [0]), .ZN(\Mpath/the_memhandle/N39 ) );
  AND2_X2 \Mpath/the_memhandle/C354  ( .A1(\m_mem_command[SIGN] ), .A2(
        \Mpath/the_memhandle/N236 ), .ZN(\Mpath/the_memhandle/N72 ) );
  AND2_X2 \Mpath/the_memhandle/C356  ( .A1(\Mpath/the_memhandle/N239 ), .A2(
        \Mpath/the_memhandle/N240 ), .ZN(\Mpath/the_memhandle/N74 ) );
  OR2_X2 \Mpath/the_memhandle/C360  ( .A1(\Mpath/mem_baddr [1]), .A2(
        \Mpath/the_memhandle/N240 ), .ZN(\Mpath/the_memhandle/N243 ) );
  INV_X2 \Mpath/the_memhandle/I_12  ( .A(\Mpath/the_memhandle/N244 ), .ZN(
        \Mpath/the_memhandle/N76 ) );
  OR2_X2 \Mpath/the_memhandle/C363  ( .A1(\Mpath/the_memhandle/N239 ), .A2(
        \Mpath/mem_baddr [0]), .ZN(\Mpath/the_memhandle/N244 ) );
  AND2_X2 \Mpath/the_memhandle/C365  ( .A1(\Mpath/mem_baddr [1]), .A2(
        \Mpath/mem_baddr [0]), .ZN(\Mpath/the_memhandle/N77 ) );
  AND2_X2 \Mpath/the_memhandle/C366  ( .A1(\Mpath/the_memhandle/N235 ), .A2(
        \Mpath/the_memhandle/N238 ), .ZN(\Mpath/the_memhandle/N86 ) );
  AND2_X2 \Mpath/the_memhandle/C369  ( .A1(\m_mem_command[SIGN] ), .A2(
        \Mpath/the_memhandle/N238 ), .ZN(\Mpath/the_memhandle/N120 ) );
  OR2_X2 \Mpath/the_shift/C151  ( .A1(shift_op[1]), .A2(\Mpath/the_shift/N104 ), .ZN(\Mpath/the_shift/N106 ) );
  OR2_X2 \Mpath/the_shift/C152  ( .A1(\Mpath/the_shift/N105 ), .A2(
        \Mpath/the_shift/N106 ), .ZN(\Mpath/the_shift/N107 ) );
  OR2_X2 \Mpath/the_shift/C155  ( .A1(shift_op[1]), .A2(\Mpath/the_shift/N104 ), .ZN(\Mpath/the_shift/N109 ) );
  OR2_X2 \Mpath/the_shift/C156  ( .A1(shift_op[0]), .A2(\Mpath/the_shift/N109 ), .ZN(\Mpath/the_shift/N110 ) );
  INV_X2 \Mpath/the_shift/I_3  ( .A(\Mpath/the_shift/N110 ), .ZN(
        \Mpath/the_shift/N111 ) );
  OR2_X2 \Mpath/the_shift/C159  ( .A1(\Mpath/the_shift/N112 ), .A2(shift_op[2]), .ZN(\Mpath/the_shift/N113 ) );
  OR2_X2 \Mpath/the_shift/C160  ( .A1(shift_op[0]), .A2(\Mpath/the_shift/N113 ), .ZN(\Mpath/the_shift/N114 ) );
  INV_X2 \Mpath/the_shift/I_5  ( .A(\Mpath/the_shift/N114 ), .ZN(
        \Mpath/the_shift/N115 ) );
  OR2_X2 \Mpath/the_shift/C163  ( .A1(shift_op[1]), .A2(shift_op[2]), .ZN(
        \Mpath/the_shift/N116 ) );
  OR2_X2 \Mpath/the_shift/C164  ( .A1(\Mpath/the_shift/N105 ), .A2(
        \Mpath/the_shift/N116 ), .ZN(\Mpath/the_shift/N117 ) );
  INV_X2 \Mpath/the_shift/I_6  ( .A(\Mpath/the_shift/N117 ), .ZN(
        \Mpath/the_shift/N118 ) );
  OR2_X2 \Mpath/the_alu/C462  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N455 ), .ZN(\Mpath/the_alu/N456 ) );
  OR2_X2 \Mpath/the_alu/C463  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N456 ), .ZN(\Mpath/the_alu/N457 ) );
  OR2_X2 \Mpath/the_alu/C468  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N461 ), .ZN(\Mpath/the_alu/N462 ) );
  OR2_X2 \Mpath/the_alu/C469  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N462 ), .ZN(\Mpath/the_alu/N463 ) );
  OR2_X2 \Mpath/the_alu/C470  ( .A1(\Alu_command[OP][0] ), .A2(
        \Mpath/the_alu/N463 ), .ZN(\Mpath/the_alu/N464 ) );
  INV_X2 \Mpath/the_alu/I_5  ( .A(\Mpath/the_alu/N464 ), .ZN(
        \Mpath/the_alu/N465 ) );
  OR2_X2 \Mpath/the_alu/C478  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N470 ), .ZN(\Mpath/the_alu/N471 ) );
  OR2_X2 \Mpath/the_alu/C479  ( .A1(\Mpath/the_alu/N467 ), .A2(
        \Mpath/the_alu/N471 ), .ZN(\Mpath/the_alu/N472 ) );
  OR2_X2 \Mpath/the_alu/C480  ( .A1(\Mpath/the_alu/N468 ), .A2(
        \Mpath/the_alu/N472 ), .ZN(\Mpath/the_alu/N473 ) );
  OR2_X2 \Mpath/the_alu/C487  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N476 ), .ZN(\Mpath/the_alu/N477 ) );
  OR2_X2 \Mpath/the_alu/C488  ( .A1(\Mpath/the_alu/N467 ), .A2(
        \Mpath/the_alu/N477 ), .ZN(\Mpath/the_alu/N478 ) );
  OR2_X2 \Mpath/the_alu/C489  ( .A1(\Alu_command[OP][0] ), .A2(
        \Mpath/the_alu/N478 ), .ZN(\Mpath/the_alu/N479 ) );
  INV_X2 \Mpath/the_alu/I_10  ( .A(\Mpath/the_alu/N479 ), .ZN(
        \Mpath/the_alu/N480 ) );
  OR2_X2 \Mpath/the_alu/C496  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N482 ), .ZN(\Mpath/the_alu/N483 ) );
  OR2_X2 \Mpath/the_alu/C497  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N483 ), .ZN(\Mpath/the_alu/N484 ) );
  OR2_X2 \Mpath/the_alu/C498  ( .A1(\Mpath/the_alu/N468 ), .A2(
        \Mpath/the_alu/N484 ), .ZN(\Mpath/the_alu/N485 ) );
  INV_X2 \Mpath/the_alu/I_11  ( .A(\Mpath/the_alu/N485 ), .ZN(
        \Mpath/the_alu/N486 ) );
  OR2_X2 \Mpath/the_alu/C504  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N488 ), .ZN(\Mpath/the_alu/N489 ) );
  OR2_X2 \Mpath/the_alu/C505  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N489 ), .ZN(\Mpath/the_alu/N490 ) );
  OR2_X2 \Mpath/the_alu/C506  ( .A1(\Alu_command[OP][0] ), .A2(
        \Mpath/the_alu/N490 ), .ZN(\Mpath/the_alu/N491 ) );
  OR2_X2 \Mpath/the_alu/C510  ( .A1(\Alu_command[OP][4] ), .A2(
        \Mpath/the_alu/N466 ), .ZN(\Mpath/the_alu/N493 ) );
  OR2_X2 \Mpath/the_alu/C512  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N494 ), .ZN(\Mpath/the_alu/N495 ) );
  OR2_X2 \Mpath/the_alu/C513  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N495 ), .ZN(\Mpath/the_alu/N496 ) );
  OR2_X2 \Mpath/the_alu/C514  ( .A1(\Mpath/the_alu/N468 ), .A2(
        \Mpath/the_alu/N496 ), .ZN(\Mpath/the_alu/N497 ) );
  INV_X2 \Mpath/the_alu/I_13  ( .A(\Mpath/the_alu/N497 ), .ZN(
        \Mpath/the_alu/N498 ) );
  OR2_X2 \Mpath/the_alu/C517  ( .A1(\Alu_command[OP][4] ), .A2(
        \Mpath/the_alu/N466 ), .ZN(\Mpath/the_alu/N499 ) );
  OR2_X2 \Mpath/the_alu/C519  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N500 ), .ZN(\Mpath/the_alu/N501 ) );
  OR2_X2 \Mpath/the_alu/C520  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N501 ), .ZN(\Mpath/the_alu/N502 ) );
  OR2_X2 \Mpath/the_alu/C521  ( .A1(\Alu_command[OP][0] ), .A2(
        \Mpath/the_alu/N502 ), .ZN(\Mpath/the_alu/N503 ) );
  OR2_X2 \Mpath/the_alu/C526  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N506 ), .ZN(\Mpath/the_alu/N507 ) );
  OR2_X2 \Mpath/the_alu/C527  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N507 ), .ZN(\Mpath/the_alu/N508 ) );
  OR2_X2 \Mpath/the_alu/C528  ( .A1(\Alu_command[OP][0] ), .A2(
        \Mpath/the_alu/N508 ), .ZN(\Mpath/the_alu/N509 ) );
  OR2_X2 \Mpath/the_alu/C534  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N512 ), .ZN(\Mpath/the_alu/N513 ) );
  OR2_X2 \Mpath/the_alu/C535  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N513 ), .ZN(\Mpath/the_alu/N514 ) );
  OR2_X2 \Mpath/the_alu/C536  ( .A1(\Mpath/the_alu/N468 ), .A2(
        \Mpath/the_alu/N514 ), .ZN(\Mpath/the_alu/N515 ) );
  OR2_X2 \Mpath/the_alu/C540  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N518 ), .ZN(\Mpath/the_alu/N519 ) );
  OR2_X2 \Mpath/the_alu/C541  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N519 ), .ZN(\Mpath/the_alu/N520 ) );
  OR2_X2 \Mpath/the_alu/C545  ( .A1(\Alu_command[OP][4] ), .A2(
        \Alu_command[OP][5] ), .ZN(\Mpath/the_alu/N523 ) );
  OR2_X2 \Mpath/the_alu/C546  ( .A1(\Alu_command[OP][3] ), .A2(
        \Mpath/the_alu/N523 ), .ZN(\Mpath/the_alu/N524 ) );
  OR2_X2 \Mpath/the_alu/C547  ( .A1(\Alu_command[OP][2] ), .A2(
        \Mpath/the_alu/N524 ), .ZN(\Mpath/the_alu/N525 ) );
  OR2_X2 \Mpath/the_alu/C548  ( .A1(\Alu_command[OP][1] ), .A2(
        \Mpath/the_alu/N525 ), .ZN(\Mpath/the_alu/N526 ) );
  AND2_X2 \Mpath/the_alu/C583  ( .A1(\Mpath/out_regA[23] ), .A2(
        \Mpath/out_regB[23] ), .ZN(\Mpath/the_alu/N102 ) );
  AND2_X2 \Mpath/the_alu/C585  ( .A1(\Mpath/out_regA[21] ), .A2(
        \Mpath/out_regB[21] ), .ZN(\Mpath/the_alu/N104 ) );
  AND2_X2 \Mpath/the_alu/C603  ( .A1(\Mpath/out_regA[3] ), .A2(n7708), .ZN(
        \Mpath/the_alu/N122 ) );
  OR2_X2 \Mpath/the_alu/C616  ( .A1(\Mpath/out_regA[23] ), .A2(
        \Mpath/out_regB[23] ), .ZN(\Mpath/the_alu/N134 ) );
  OR2_X2 \Mpath/the_alu/C636  ( .A1(\Mpath/out_regA[3] ), .A2(n7708), .ZN(
        \Mpath/the_alu/N154 ) );
  XOR2_X1 \Mpath/the_alu/C649  ( .A(\Mpath/out_regA[23] ), .B(
        \Mpath/out_regB[23] ), .Z(\Mpath/the_alu/N166 ) );
  XOR2_X1 \Mpath/the_alu/C650  ( .A(\Mpath/out_regA[22] ), .B(
        \Mpath/out_regB[22] ), .Z(\Mpath/the_alu/N167 ) );
  XOR2_X1 \Mpath/the_alu/C651  ( .A(\Mpath/out_regA[21] ), .B(
        \Mpath/out_regB[21] ), .Z(\Mpath/the_alu/N168 ) );
  XOR2_X1 \Mpath/the_alu/C652  ( .A(\Mpath/out_regA[20] ), .B(n7476), .Z(
        \Mpath/the_alu/N169 ) );
  XOR2_X1 \Mpath/the_alu/C653  ( .A(\Mpath/out_regA[19] ), .B(n7333), .Z(
        \Mpath/the_alu/N170 ) );
  XOR2_X1 \Mpath/the_alu/C654  ( .A(\Mpath/out_regA[18] ), .B(n7361), .Z(
        \Mpath/the_alu/N171 ) );
  XOR2_X1 \Mpath/the_alu/C655  ( .A(\Mpath/out_regA[17] ), .B(n7344), .Z(
        \Mpath/the_alu/N172 ) );
  XOR2_X1 \Mpath/the_alu/C656  ( .A(\Mpath/out_regA[16] ), .B(n7388), .Z(
        \Mpath/the_alu/N173 ) );
  XOR2_X1 \Mpath/the_alu/C657  ( .A(\Mpath/out_regA[15] ), .B(n7323), .Z(
        \Mpath/the_alu/N174 ) );
  XOR2_X1 \Mpath/the_alu/C658  ( .A(\Mpath/out_regA[14] ), .B(n7395), .Z(
        \Mpath/the_alu/N175 ) );
  XOR2_X1 \Mpath/the_alu/C659  ( .A(\Mpath/out_regA[13] ), .B(n7106), .Z(
        \Mpath/the_alu/N176 ) );
  XOR2_X1 \Mpath/the_alu/C660  ( .A(n7182), .B(\Mpath/out_regB[12] ), .Z(
        \Mpath/the_alu/N177 ) );
  XOR2_X1 \Mpath/the_alu/C661  ( .A(\Mpath/out_regA[11] ), .B(
        \Mpath/out_regB[11] ), .Z(\Mpath/the_alu/N178 ) );
  XOR2_X1 \Mpath/the_alu/C662  ( .A(\Mpath/out_regA[10] ), .B(n7192), .Z(
        \Mpath/the_alu/N179 ) );
  XOR2_X1 \Mpath/the_alu/C663  ( .A(\Mpath/out_regA[9] ), .B(
        \Mpath/out_regB[9] ), .Z(\Mpath/the_alu/N180 ) );
  XOR2_X1 \Mpath/the_alu/C664  ( .A(n7185), .B(n7616), .Z(\Mpath/the_alu/N181 ) );
  XOR2_X1 \Mpath/the_alu/C665  ( .A(\Mpath/out_regA[7] ), .B(
        \Mpath/out_regB[7] ), .Z(\Mpath/the_alu/N182 ) );
  XOR2_X1 \Mpath/the_alu/C666  ( .A(\Mpath/out_regA[6] ), .B(
        \Mpath/out_regB[6] ), .Z(\Mpath/the_alu/N183 ) );
  XOR2_X1 \Mpath/the_alu/C667  ( .A(\Mpath/out_regA[5] ), .B(
        \Mpath/out_regB[5] ), .Z(\Mpath/the_alu/N184 ) );
  XOR2_X1 \Mpath/the_alu/C668  ( .A(\Mpath/out_regA[4] ), .B(n7707), .Z(
        \Mpath/the_alu/N185 ) );
  XOR2_X1 \Mpath/the_alu/C669  ( .A(\Mpath/out_regA[3] ), .B(n7708), .Z(
        \Mpath/the_alu/N186 ) );
  XOR2_X1 \Mpath/the_alu/C670  ( .A(\Mpath/out_regA[2] ), .B(n7711), .Z(
        \Mpath/the_alu/N187 ) );
  XOR2_X1 \Mpath/the_alu/C672  ( .A(\Mpath/out_regA[0] ), .B(n7715), .Z(
        \Mpath/the_alu/N189 ) );
  AND2_X2 \Mpath/the_alu/C682  ( .A1(\Mpath/the_alu/N37 ), .A2(
        \Mpath/the_alu/N38 ), .ZN(\Mpath/the_alu/N198 ) );
  AND2_X2 \Mpath/the_alu/C683  ( .A1(\Mpath/the_alu/N39 ), .A2(
        \Mpath/the_alu/N40 ), .ZN(\Mpath/the_alu/N199 ) );
  AND2_X2 \Mpath/the_alu/C684  ( .A1(\Mpath/the_alu/N41 ), .A2(
        \Mpath/the_alu/N42 ), .ZN(\Mpath/the_alu/N200 ) );
  AND2_X2 \Mpath/the_alu/C685  ( .A1(\Mpath/the_alu/N43 ), .A2(
        \Mpath/the_alu/N44 ), .ZN(\Mpath/the_alu/N201 ) );
  AND2_X2 \Mpath/the_alu/C686  ( .A1(\Mpath/the_alu/N45 ), .A2(
        \Mpath/the_alu/N46 ), .ZN(\Mpath/the_alu/N202 ) );
  AND2_X2 \Mpath/the_alu/C687  ( .A1(\Mpath/the_alu/N47 ), .A2(
        \Mpath/the_alu/N48 ), .ZN(\Mpath/the_alu/N203 ) );
  AND2_X2 \Mpath/the_alu/C688  ( .A1(\Mpath/the_alu/N49 ), .A2(
        \Mpath/the_alu/N50 ), .ZN(\Mpath/the_alu/N204 ) );
  AND2_X2 \Mpath/the_alu/C689  ( .A1(\Mpath/the_alu/N51 ), .A2(
        \Mpath/the_alu/N52 ), .ZN(\Mpath/the_alu/N205 ) );
  AND2_X2 \Mpath/the_alu/C690  ( .A1(\Mpath/the_alu/N53 ), .A2(
        \Mpath/the_alu/N54 ), .ZN(\Mpath/the_alu/N206 ) );
  AND2_X2 \Mpath/the_alu/C691  ( .A1(\Mpath/the_alu/N55 ), .A2(
        \Mpath/the_alu/N56 ), .ZN(\Mpath/the_alu/N207 ) );
  AND2_X2 \Mpath/the_alu/C692  ( .A1(\Mpath/the_alu/N57 ), .A2(
        \Mpath/the_alu/N58 ), .ZN(\Mpath/the_alu/N208 ) );
  AND2_X2 \Mpath/the_alu/C693  ( .A1(\Mpath/the_alu/N59 ), .A2(
        \Mpath/the_alu/N60 ), .ZN(\Mpath/the_alu/N209 ) );
  AND2_X2 \Mpath/the_alu/C694  ( .A1(\Mpath/the_alu/N61 ), .A2(
        \Mpath/the_alu/N62 ), .ZN(\Mpath/the_alu/N210 ) );
  AND2_X2 \Mpath/the_alu/C695  ( .A1(\Mpath/the_alu/N63 ), .A2(
        \Mpath/the_alu/N64 ), .ZN(\Mpath/the_alu/N211 ) );
  AND2_X2 \Mpath/the_alu/C696  ( .A1(\Mpath/the_alu/N65 ), .A2(
        \Mpath/the_alu/N66 ), .ZN(\Mpath/the_alu/N212 ) );
  AND2_X2 \Mpath/the_alu/C697  ( .A1(n7184), .A2(\Mpath/the_alu/N68 ), .ZN(
        \Mpath/the_alu/N213 ) );
  AND2_X2 \Mpath/the_alu/C698  ( .A1(\Mpath/the_alu/N69 ), .A2(
        \Mpath/the_alu/N70 ), .ZN(\Mpath/the_alu/N214 ) );
  AND2_X2 \Mpath/the_alu/C699  ( .A1(\Mpath/the_alu/N71 ), .A2(
        \Mpath/the_alu/N72 ), .ZN(\Mpath/the_alu/N215 ) );
  AND2_X2 \Mpath/the_alu/C700  ( .A1(\Mpath/the_alu/N73 ), .A2(
        \Mpath/the_alu/N74 ), .ZN(\Mpath/the_alu/N216 ) );
  AND2_X2 \Mpath/the_alu/C701  ( .A1(\Mpath/the_alu/N75 ), .A2(
        \Mpath/the_alu/N76 ), .ZN(\Mpath/the_alu/N217 ) );
  AND2_X2 \Mpath/the_alu/C702  ( .A1(\Mpath/the_alu/N77 ), .A2(
        \Mpath/the_alu/N78 ), .ZN(\Mpath/the_alu/N218 ) );
  AND2_X2 \Mpath/the_alu/C703  ( .A1(\Mpath/the_alu/N79 ), .A2(
        \Mpath/the_alu/N80 ), .ZN(\Mpath/the_alu/N219 ) );
  AND2_X2 \Mpath/the_alu/C705  ( .A1(\Mpath/the_alu/N83 ), .A2(
        \Mpath/the_alu/N84 ), .ZN(\Mpath/the_alu/N221 ) );
  OR2_X2 \Mpath/C335  ( .A1(exe_outsel[1]), .A2(\Mpath/N179 ), .ZN(
        \Mpath/N181 ) );
  OR2_X2 \Mpath/C336  ( .A1(\Mpath/N180 ), .A2(\Mpath/N181 ), .ZN(\Mpath/N182 ) );
  INV_X2 \Mpath/I_3  ( .A(\Mpath/N182 ), .ZN(\Mpath/N183 ) );
  OR2_X2 \Mpath/C340  ( .A1(exe_outsel[1]), .A2(\Mpath/N179 ), .ZN(
        \Mpath/N184 ) );
  OR2_X2 \Mpath/C341  ( .A1(\Mpath/N180 ), .A2(\Mpath/N184 ), .ZN(\Mpath/N185 ) );
  INV_X2 \Mpath/I_4  ( .A(\Mpath/N185 ), .ZN(\Mpath/N186 ) );
  OR2_X2 \Mpath/C344  ( .A1(\Mpath/N187 ), .A2(exe_outsel[2]), .ZN(
        \Mpath/N188 ) );
  OR2_X2 \Mpath/C345  ( .A1(exe_outsel[0]), .A2(\Mpath/N188 ), .ZN(
        \Mpath/N189 ) );
  INV_X2 \Mpath/I_6  ( .A(\Mpath/N189 ), .ZN(\Mpath/N190 ) );
  OR2_X2 \Mpath/C355  ( .A1(exe_outsel[1]), .A2(\Mpath/N179 ), .ZN(
        \Mpath/N196 ) );
  OR2_X2 \Mpath/C356  ( .A1(\Mpath/N180 ), .A2(\Mpath/N196 ), .ZN(\Mpath/N197 ) );
  INV_X2 \Mcontrol/st_logic/I_0  ( .A(\Mcontrol/st_logic/load_stall ), .ZN(
        \Mcontrol/st_logic/N12 ) );
  INV_X2 \Mcontrol/st_logic/I_2  ( .A(\Mcontrol/st_logic/branchmul_stall ), 
        .ZN(\Mcontrol/st_logic/N14 ) );
  INV_X2 \Mcontrol/st_logic/I_3  ( .A(\x_mem_command[MR] ), .ZN(
        \Mcontrol/st_logic/N15 ) );
  INV_X2 \Mcontrol/st_logic/I_5  ( .A(\Mcontrol/st_logic/N18 ), .ZN(
        \Mcontrol/st_logic/N19 ) );
  INV_X2 \Mcontrol/st_logic/I_6  ( .A(byp_controlB[2]), .ZN(
        \Mcontrol/st_logic/N52 ) );
  OR2_X2 \Mcontrol/st_logic/C79  ( .A1(byp_controlB[0]), .A2(
        \Mcontrol/st_logic/N52 ), .ZN(\Mcontrol/st_logic/N22 ) );
  INV_X2 \Mcontrol/st_logic/I_7  ( .A(\Mcontrol/st_logic/N22 ), .ZN(
        \Mcontrol/st_logic/N23 ) );
  INV_X2 \Mcontrol/st_logic/I_8  ( .A(\m_mem_command[MR] ), .ZN(
        \Mcontrol/st_logic/N24 ) );
  OR2_X2 \Mcontrol/st_logic/C85  ( .A1(\Mcontrol/x_mul_command [4]), .A2(
        \Mcontrol/x_mul_command [5]), .ZN(\Mcontrol/st_logic/N28 ) );
  OR2_X2 \Mcontrol/st_logic/C86  ( .A1(\Mcontrol/x_mul_command [3]), .A2(
        \Mcontrol/st_logic/N28 ), .ZN(\Mcontrol/st_logic/N29 ) );
  OR2_X2 \Mcontrol/st_logic/C87  ( .A1(\Mcontrol/st_logic/N26 ), .A2(
        \Mcontrol/st_logic/N29 ), .ZN(\Mcontrol/st_logic/N30 ) );
  OR2_X2 \Mcontrol/st_logic/C88  ( .A1(\Mcontrol/st_logic/N27 ), .A2(
        \Mcontrol/st_logic/N30 ), .ZN(\Mcontrol/st_logic/N31 ) );
  OR2_X2 \Mcontrol/st_logic/C89  ( .A1(\Mcontrol/x_mul_command [0]), .A2(
        \Mcontrol/st_logic/N31 ), .ZN(\Mcontrol/st_logic/N32 ) );
  INV_X2 \Mcontrol/st_logic/I_12  ( .A(\Mcontrol/st_logic/N32 ), .ZN(
        \Mcontrol/st_logic/N33 ) );
  OR2_X2 \Mcontrol/st_logic/C94  ( .A1(\Mcontrol/x_mul_command [4]), .A2(
        \Mcontrol/x_mul_command [5]), .ZN(\Mcontrol/st_logic/N35 ) );
  OR2_X2 \Mcontrol/st_logic/C95  ( .A1(\Mcontrol/x_mul_command [3]), .A2(
        \Mcontrol/st_logic/N35 ), .ZN(\Mcontrol/st_logic/N36 ) );
  OR2_X2 \Mcontrol/st_logic/C96  ( .A1(\Mcontrol/st_logic/N26 ), .A2(
        \Mcontrol/st_logic/N36 ), .ZN(\Mcontrol/st_logic/N37 ) );
  OR2_X2 \Mcontrol/st_logic/C97  ( .A1(\Mcontrol/st_logic/N27 ), .A2(
        \Mcontrol/st_logic/N37 ), .ZN(\Mcontrol/st_logic/N38 ) );
  OR2_X2 \Mcontrol/st_logic/C98  ( .A1(\Mcontrol/st_logic/N34 ), .A2(
        \Mcontrol/st_logic/N38 ), .ZN(\Mcontrol/st_logic/N39 ) );
  INV_X2 \Mcontrol/st_logic/I_14  ( .A(\Mcontrol/st_logic/N39 ), .ZN(
        \Mcontrol/st_logic/N40 ) );
  INV_X2 \Mcontrol/st_logic/I_15  ( .A(
        \Mcontrol/st_logic/branch_uses_main_exe_result ), .ZN(
        \Mcontrol/st_logic/N41 ) );
  OR2_X2 \Mcontrol/st_logic/C104  ( .A1(\Mcontrol/st_logic/N42 ), .A2(
        \Mcontrol/st_logic/N52 ), .ZN(\Mcontrol/st_logic/N44 ) );
  INV_X2 \Mcontrol/st_logic/I_17  ( .A(\Mcontrol/st_logic/N44 ), .ZN(
        \Mcontrol/st_logic/N45 ) );
  INV_X2 \Mcontrol/st_logic/I_18  ( .A(\Mcontrol/st_logic/branch_uses_regb ), 
        .ZN(\Mcontrol/st_logic/N46 ) );
  INV_X2 \Mcontrol/st_logic/I_20  ( .A(\Mcontrol/st_logic/N49 ), .ZN(
        \Mcontrol/st_logic/N50 ) );
  OR2_X2 \Mcontrol/st_logic/C115  ( .A1(byp_controlB[0]), .A2(
        \Mcontrol/st_logic/N52 ), .ZN(\Mcontrol/st_logic/N53 ) );
  INV_X2 \Mcontrol/st_logic/I_22  ( .A(\Mcontrol/st_logic/N53 ), .ZN(
        \Mcontrol/st_logic/N54 ) );
  INV_X2 \Mcontrol/st_logic/I_23  ( .A(\Mcontrol/st_logic/N56 ), .ZN(
        \Mcontrol/st_logic/N57 ) );
  INV_X2 \Mcontrol/st_logic/I_24  ( .A(\Mcontrol/d_jump_type[2] ), .ZN(
        \Mcontrol/st_logic/N58 ) );
  OR2_X2 \Mcontrol/st_logic/C126  ( .A1(\Mcontrol/st_logic/N58 ), .A2(
        \Mcontrol/st_logic/N60 ), .ZN(\Mcontrol/st_logic/N61 ) );
  OR2_X2 \Mcontrol/st_logic/C127  ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/st_logic/N61 ), .ZN(\Mcontrol/st_logic/N62 ) );
  INV_X2 \Mcontrol/st_logic/I_25  ( .A(\Mcontrol/st_logic/N63 ), .ZN(
        \Mcontrol/st_logic/N64 ) );
  OR2_X2 \Mcontrol/st_logic/C134  ( .A1(\Mcontrol/st_logic/N58 ), .A2(
        \Mcontrol/st_logic/N67 ), .ZN(\Mcontrol/st_logic/N68 ) );
  OR2_X2 \Mcontrol/st_logic/C135  ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/st_logic/N68 ), .ZN(\Mcontrol/st_logic/N69 ) );
  INV_X2 \Mcontrol/st_logic/I_27  ( .A(\Mcontrol/st_logic/N70 ), .ZN(
        \Mcontrol/st_logic/N71 ) );
  INV_X2 \Mcontrol/st_logic/I_28  ( .A(\Mcontrol/st_logic/N76 ), .ZN(
        \Mcontrol/st_logic/N77 ) );
  OR2_X2 \Mcontrol/st_logic/C149  ( .A1(\Mcontrol/st_logic/N58 ), .A2(
        \Mcontrol/st_logic/N79 ), .ZN(\Mcontrol/st_logic/N80 ) );
  OR2_X2 \Mcontrol/st_logic/C150  ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/st_logic/N80 ), .ZN(\Mcontrol/st_logic/N81 ) );
  OR2_X2 \Mcontrol/st_logic/C151  ( .A1(\Mcontrol/st_logic/N65 ), .A2(
        \Mcontrol/st_logic/N81 ), .ZN(\Mcontrol/st_logic/N82 ) );
  OR2_X2 \Mcontrol/st_logic/C155  ( .A1(\Mcontrol/d_jump_type[2] ), .A2(
        \Mcontrol/st_logic/N85 ), .ZN(\Mcontrol/st_logic/N86 ) );
  OR2_X2 \Mcontrol/st_logic/C156  ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/st_logic/N86 ), .ZN(\Mcontrol/st_logic/N87 ) );
  INV_X2 \Mcontrol/st_logic/I_31  ( .A(\Mcontrol/d_jump_type[1] ), .ZN(
        \Mcontrol/st_logic/N90 ) );
  OR2_X2 \Mcontrol/st_logic/C163  ( .A1(\Mcontrol/d_jump_type[2] ), .A2(
        \Mcontrol/st_logic/N92 ), .ZN(\Mcontrol/st_logic/N93 ) );
  OR2_X2 \Mcontrol/st_logic/C164  ( .A1(\Mcontrol/st_logic/N90 ), .A2(
        \Mcontrol/st_logic/N93 ), .ZN(\Mcontrol/st_logic/N94 ) );
  OR2_X2 \Mcontrol/st_logic/C171  ( .A1(\Mcontrol/st_logic/N58 ), .A2(
        \Mcontrol/st_logic/N98 ), .ZN(\Mcontrol/st_logic/N99 ) );
  OR2_X2 \Mcontrol/st_logic/C172  ( .A1(\Mcontrol/st_logic/N90 ), .A2(
        \Mcontrol/st_logic/N99 ), .ZN(\Mcontrol/st_logic/N100 ) );
  INV_X2 \Mcontrol/st_logic/I_33  ( .A(\Mcontrol/st_logic/N101 ), .ZN(
        \Mcontrol/st_logic/N102 ) );
  OR2_X2 \Mcontrol/st_logic/C179  ( .A1(\Mcontrol/d_jump_type[2] ), .A2(
        \Mcontrol/st_logic/N105 ), .ZN(\Mcontrol/st_logic/N106 ) );
  OR2_X2 \Mcontrol/st_logic/C180  ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/st_logic/N106 ), .ZN(\Mcontrol/st_logic/N107 ) );
  INV_X2 \Mcontrol/st_logic/I_35  ( .A(\Mcontrol/st_logic/N108 ), .ZN(
        \Mcontrol/st_logic/N109 ) );
  AND2_X2 \Mcontrol/st_logic/C193  ( .A1(\Mcontrol/st_logic/N15 ), .A2(
        \Mcontrol/st_logic/N110 ), .ZN(\Mcontrol/st_logic/N2 ) );
  OR2_X2 \Mcontrol/st_logic/C194  ( .A1(\Mcontrol/st_logic/N19 ), .A2(
        \Mcontrol/st_logic/N23 ), .ZN(\Mcontrol/st_logic/N110 ) );
  OR2_X2 \Mcontrol/st_logic/C195  ( .A1(\Mcontrol/st_logic/N114 ), .A2(
        \Mcontrol/st_logic/N109 ), .ZN(\Mcontrol/st_logic/N3 ) );
  OR2_X2 \Mcontrol/st_logic/C196  ( .A1(\Mcontrol/st_logic/N113 ), .A2(
        \Mcontrol/st_logic/N102 ), .ZN(\Mcontrol/st_logic/N114 ) );
  OR2_X2 \Mcontrol/st_logic/C200  ( .A1(\Mcontrol/st_logic/N64 ), .A2(
        \Mcontrol/st_logic/N71 ), .ZN(\Mcontrol/st_logic/N4 ) );
  OR2_X2 \Mcontrol/st_logic/C201  ( .A1(\Mcontrol/st_logic/N115 ), .A2(
        \Mcontrol/st_logic/N116 ), .ZN(\Mcontrol/st_logic/N5 ) );
  AND2_X2 \Mcontrol/st_logic/C202  ( .A1(\Mcontrol/st_logic/N45 ), .A2(
        \Mcontrol/st_logic/N46 ), .ZN(\Mcontrol/st_logic/N115 ) );
  AND2_X2 \Mcontrol/st_logic/C203  ( .A1(\Mcontrol/st_logic/N50 ), .A2(
        \Mcontrol/st_logic/N51 ), .ZN(\Mcontrol/st_logic/N116 ) );
  AND2_X2 \Mcontrol/st_logic/C204  ( .A1(\Mcontrol/st_logic/N24 ), .A2(
        \Mcontrol/st_logic/N25 ), .ZN(\Mcontrol/st_logic/N6 ) );
  OR2_X2 \Mcontrol/st_logic/C205  ( .A1(\Mcontrol/st_logic/N117 ), .A2(
        \Mcontrol/st_logic/N118 ), .ZN(\Mcontrol/st_logic/N7 ) );
  AND2_X2 \Mcontrol/st_logic/C206  ( .A1(\Mcontrol/st_logic/N54 ), .A2(
        \Mcontrol/st_logic/N46 ), .ZN(\Mcontrol/st_logic/N117 ) );
  AND2_X2 \Mcontrol/st_logic/C208  ( .A1(\Mcontrol/st_logic/N119 ), .A2(
        \Mcontrol/st_logic/N41 ), .ZN(\Mcontrol/st_logic/N8 ) );
  OR2_X2 \Mcontrol/st_logic/C209  ( .A1(\Mcontrol/st_logic/N33 ), .A2(
        \Mcontrol/st_logic/N40 ), .ZN(\Mcontrol/st_logic/N119 ) );
  OR2_X2 \Mcontrol/st_logic/C211  ( .A1(\Mcontrol/st_logic/N120 ), .A2(
        \Mcontrol/st_logic/N14 ), .ZN(\Mcontrol/st_logic/N10 ) );
  OR2_X2 \Mcontrol/st_logic/C212  ( .A1(\Mcontrol/st_logic/N12 ), .A2(
        \Mcontrol/st_logic/N13 ), .ZN(\Mcontrol/st_logic/N120 ) );
  OR2_X2 \Mcontrol/bp_logicB/C19  ( .A1(\Mcontrol/x_rd[3] ), .A2(
        \Mcontrol/x_rd[4] ), .ZN(\Mcontrol/bp_logicB/N5 ) );
  OR2_X2 \Mcontrol/bp_logicB/C20  ( .A1(\Mcontrol/x_rd[2] ), .A2(
        \Mcontrol/bp_logicB/N5 ), .ZN(\Mcontrol/bp_logicB/N6 ) );
  OR2_X2 \Mcontrol/bp_logicB/C21  ( .A1(\Mcontrol/x_rd[1] ), .A2(
        \Mcontrol/bp_logicB/N6 ), .ZN(\Mcontrol/bp_logicB/N7 ) );
  OR2_X2 \Mcontrol/bp_logicB/C22  ( .A1(\Mcontrol/x_rd[0] ), .A2(
        \Mcontrol/bp_logicB/N7 ), .ZN(\Mcontrol/bp_logicB/N8 ) );
  INV_X2 \Mcontrol/bp_logicB/I_1  ( .A(\Mcontrol/x_sampled_dwe ), .ZN(
        \Mcontrol/bp_logicB/N9 ) );
  OR2_X2 \Mcontrol/bp_logicB/C26  ( .A1(\Mcontrol/m_sampled_xrd[3] ), .A2(
        \Mcontrol/m_sampled_xrd[4] ), .ZN(\Mcontrol/bp_logicB/N10 ) );
  OR2_X2 \Mcontrol/bp_logicB/C27  ( .A1(\Mcontrol/m_sampled_xrd[2] ), .A2(
        \Mcontrol/bp_logicB/N10 ), .ZN(\Mcontrol/bp_logicB/N11 ) );
  OR2_X2 \Mcontrol/bp_logicB/C28  ( .A1(\Mcontrol/m_sampled_xrd[1] ), .A2(
        \Mcontrol/bp_logicB/N11 ), .ZN(\Mcontrol/bp_logicB/N12 ) );
  OR2_X2 \Mcontrol/bp_logicB/C29  ( .A1(\Mcontrol/m_sampled_xrd[0] ), .A2(
        \Mcontrol/bp_logicB/N12 ), .ZN(\Mcontrol/bp_logicB/N13 ) );
  INV_X2 \Mcontrol/bp_logicB/I_3  ( .A(m_we), .ZN(\Mcontrol/bp_logicB/N14 ) );
  AND2_X2 \Mcontrol/bp_logicB/C36  ( .A1(\Mcontrol/bp_logicB/N15 ), .A2(
        \Mcontrol/bp_logicB/N9 ), .ZN(\Mcontrol/bp_logicB/exec_main ) );
  AND2_X2 \Mcontrol/bp_logicB/C38  ( .A1(\Mcontrol/bp_logicB/N16 ), .A2(
        \Mcontrol/bp_logicB/N14 ), .ZN(\Mcontrol/bp_logicB/memory_main ) );
  OR2_X2 \Mcontrol/bp_logicA/C19  ( .A1(\Mcontrol/x_rd[3] ), .A2(
        \Mcontrol/x_rd[4] ), .ZN(\Mcontrol/bp_logicA/N5 ) );
  OR2_X2 \Mcontrol/bp_logicA/C20  ( .A1(\Mcontrol/x_rd[2] ), .A2(
        \Mcontrol/bp_logicA/N5 ), .ZN(\Mcontrol/bp_logicA/N6 ) );
  OR2_X2 \Mcontrol/bp_logicA/C21  ( .A1(\Mcontrol/x_rd[1] ), .A2(
        \Mcontrol/bp_logicA/N6 ), .ZN(\Mcontrol/bp_logicA/N7 ) );
  OR2_X2 \Mcontrol/bp_logicA/C22  ( .A1(\Mcontrol/x_rd[0] ), .A2(
        \Mcontrol/bp_logicA/N7 ), .ZN(\Mcontrol/bp_logicA/N8 ) );
  OR2_X2 \Mcontrol/bp_logicA/C26  ( .A1(\Mcontrol/m_sampled_xrd[3] ), .A2(
        \Mcontrol/m_sampled_xrd[4] ), .ZN(\Mcontrol/bp_logicA/N10 ) );
  OR2_X2 \Mcontrol/bp_logicA/C27  ( .A1(\Mcontrol/m_sampled_xrd[2] ), .A2(
        \Mcontrol/bp_logicA/N10 ), .ZN(\Mcontrol/bp_logicA/N11 ) );
  OR2_X2 \Mcontrol/bp_logicA/C28  ( .A1(\Mcontrol/m_sampled_xrd[1] ), .A2(
        \Mcontrol/bp_logicA/N11 ), .ZN(\Mcontrol/bp_logicA/N12 ) );
  OR2_X2 \Mcontrol/bp_logicA/C29  ( .A1(\Mcontrol/m_sampled_xrd[0] ), .A2(
        \Mcontrol/bp_logicA/N12 ), .ZN(\Mcontrol/bp_logicA/N13 ) );
  AND2_X2 \Mcontrol/bp_logicA/C38  ( .A1(\Mcontrol/bp_logicA/N16 ), .A2(
        \Mcontrol/bp_logicA/N14 ), .ZN(\Mcontrol/bp_logicA/memory_main ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C254  ( .A1(\Mcontrol/d_jump_type[2] ), 
        .A2(\Mcontrol/Nextpc_decoding/N182 ), .ZN(
        \Mcontrol/Nextpc_decoding/N168 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C255  ( .A1(\Mcontrol/d_jump_type[1] ), 
        .A2(\Mcontrol/Nextpc_decoding/N168 ), .ZN(
        \Mcontrol/Nextpc_decoding/N169 ) );
  INV_X2 \Mcontrol/Nextpc_decoding/I_2  ( .A(\Mcontrol/Nextpc_decoding/N170 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N171 ) );
  INV_X2 \Mcontrol/Nextpc_decoding/I_13  ( .A(\Mcontrol/d_jump_type[2] ), .ZN(
        \Mcontrol/Nextpc_decoding/N283 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C382  ( .A1(\Mcontrol/Nextpc_decoding/N283 ), .A2(\Mcontrol/Nextpc_decoding/N285 ), .ZN(\Mcontrol/Nextpc_decoding/N286 )
         );
  INV_X2 \Mcontrol/Nextpc_decoding/I_14  ( .A(\Mcontrol/Nextpc_decoding/N288 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N289 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C390  ( .A1(\Mcontrol/d_jump_type[2] ), 
        .A2(\Mcontrol/Nextpc_decoding/N291 ), .ZN(
        \Mcontrol/Nextpc_decoding/N292 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C392  ( .A1(\Mcontrol/Nextpc_decoding/N173 ), .A2(\Mcontrol/Nextpc_decoding/N293 ), .ZN(\Mcontrol/Nextpc_decoding/N294 )
         );
  OR2_X2 \Mcontrol/Nextpc_decoding/C397  ( .A1(\Mcontrol/d_jump_type[2] ), 
        .A2(\Mcontrol/Nextpc_decoding/N297 ), .ZN(
        \Mcontrol/Nextpc_decoding/N298 ) );
  INV_X2 \Mcontrol/Nextpc_decoding/I_16  ( .A(\Mcontrol/Nextpc_decoding/N300 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N301 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C404  ( .A1(\Mcontrol/d_jump_type[2] ), 
        .A2(\Mcontrol/Nextpc_decoding/N303 ), .ZN(
        \Mcontrol/Nextpc_decoding/N304 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C405  ( .A1(n6953), .A2(
        \Mcontrol/Nextpc_decoding/N304 ), .ZN(\Mcontrol/Nextpc_decoding/N305 )
         );
  OR2_X2 \Mcontrol/Nextpc_decoding/C406  ( .A1(\Mcontrol/Nextpc_decoding/N173 ), .A2(\Mcontrol/Nextpc_decoding/N305 ), .ZN(\Mcontrol/Nextpc_decoding/N306 )
         );
  INV_X2 \Mcontrol/Nextpc_decoding/I_17  ( .A(\Mcontrol/Nextpc_decoding/N306 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N307 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C410  ( .A1(\Mcontrol/d_jump_type[2] ), 
        .A2(\Mcontrol/Nextpc_decoding/N309 ), .ZN(
        \Mcontrol/Nextpc_decoding/N310 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C411  ( .A1(n6953), .A2(
        \Mcontrol/Nextpc_decoding/N310 ), .ZN(\Mcontrol/Nextpc_decoding/N311 )
         );
  INV_X2 \Mcontrol/Nextpc_decoding/I_18  ( .A(\Mcontrol/Nextpc_decoding/N312 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N313 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C418  ( .A1(\Mcontrol/Nextpc_decoding/N283 ), .A2(\Mcontrol/Nextpc_decoding/N315 ), .ZN(\Mcontrol/Nextpc_decoding/N316 )
         );
  OR2_X2 \Mcontrol/Nextpc_decoding/C419  ( .A1(n6953), .A2(
        \Mcontrol/Nextpc_decoding/N316 ), .ZN(\Mcontrol/Nextpc_decoding/N317 )
         );
  OR2_X2 \Mcontrol/Nextpc_decoding/C420  ( .A1(\Mcontrol/Nextpc_decoding/N173 ), .A2(\Mcontrol/Nextpc_decoding/N317 ), .ZN(\Mcontrol/Nextpc_decoding/N318 )
         );
  INV_X2 \Mcontrol/Nextpc_decoding/I_19  ( .A(\Mcontrol/Nextpc_decoding/N318 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N319 ) );
  OR2_X2 \Mcontrol/Nextpc_decoding/C425  ( .A1(\Mcontrol/Nextpc_decoding/N283 ), .A2(\Mcontrol/Nextpc_decoding/N321 ), .ZN(\Mcontrol/Nextpc_decoding/N322 )
         );
  OR2_X2 \Mcontrol/Nextpc_decoding/C426  ( .A1(n6953), .A2(
        \Mcontrol/Nextpc_decoding/N322 ), .ZN(\Mcontrol/Nextpc_decoding/N323 )
         );
  AND2_X2 \Mcontrol/Operation_decoding32/C2059  ( .A1(\Mcontrol/d_instr [3]), 
        .A2(\Mcontrol/Operation_decoding32/N1883 ), .ZN(
        \Mcontrol/Operation_decoding32/N1884 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2060  ( .A1(\Mcontrol/d_instr [2]), 
        .A2(\Mcontrol/Operation_decoding32/N1884 ), .ZN(
        \Mcontrol/Operation_decoding32/N1885 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2061  ( .A1(\Mcontrol/d_instr [1]), 
        .A2(\Mcontrol/Operation_decoding32/N1885 ), .ZN(
        \Mcontrol/Operation_decoding32/N1886 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2071  ( .A1(net56765), .A2(
        \Mcontrol/Operation_decoding32/N1892 ), .ZN(
        \Mcontrol/Operation_decoding32/N1893 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2076  ( .A1(\Mcontrol/d_instr [2]), 
        .A2(\Mcontrol/Operation_decoding32/N1895 ), .ZN(
        \Mcontrol/Operation_decoding32/N1896 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2077  ( .A1(\Mcontrol/d_instr [1]), 
        .A2(\Mcontrol/Operation_decoding32/N1896 ), .ZN(
        \Mcontrol/Operation_decoding32/N1897 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2084  ( .A1(\Mcontrol/d_instr [2]), 
        .A2(\Mcontrol/Operation_decoding32/N1903 ), .ZN(
        \Mcontrol/Operation_decoding32/N1904 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2085  ( .A1(\Mcontrol/d_instr [1]), 
        .A2(\Mcontrol/Operation_decoding32/N1904 ), .ZN(
        \Mcontrol/Operation_decoding32/N1905 ) );
  INV_X2 \Mcontrol/Operation_decoding32/I_9  ( .A(
        \Mcontrol/Operation_decoding32/N1906 ), .ZN(
        \Mcontrol/Operation_decoding32/N1907 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2090  ( .A1(\Mcontrol/d_instr [2]), 
        .A2(\Mcontrol/Operation_decoding32/N1909 ), .ZN(
        \Mcontrol/Operation_decoding32/N1910 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2091  ( .A1(\Mcontrol/d_instr [1]), 
        .A2(\Mcontrol/Operation_decoding32/N1910 ), .ZN(
        \Mcontrol/Operation_decoding32/N1911 ) );
  INV_X2 \Mcontrol/Operation_decoding32/I_10  ( .A(
        \Mcontrol/Operation_decoding32/N1912 ), .ZN(
        \Mcontrol/Operation_decoding32/N1913 ) );
  INV_X2 \Mcontrol/Operation_decoding32/I_11  ( .A(
        \Mcontrol/Operation_decoding32/N1914 ), .ZN(
        \Mcontrol/Operation_decoding32/N1915 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2606  ( .A1(
        \Mcontrol/Operation_decoding32/N1913 ), .A2(
        \Mcontrol/Operation_decoding32/N1915 ), .ZN(
        \Mcontrol/Operation_decoding32/N62 ) );
  OR2_X2 \Mcontrol/bvgen/C39  ( .A1(\Mcontrol/bvgen/N2 ), .A2(
        \Mcontrol/bvgen/N6 ), .ZN(\Mcontrol/bvgen/N7 ) );
  OR2_X2 \Mcontrol/bvgen/C40  ( .A1(\Mcontrol/bvgen/N3 ), .A2(
        \Mcontrol/bvgen/N7 ), .ZN(\Mcontrol/bvgen/N8 ) );
  OR2_X2 \Mcontrol/bvgen/C41  ( .A1(\Mcontrol/bvgen/N4 ), .A2(
        \Mcontrol/bvgen/N8 ), .ZN(\Mcontrol/bvgen/N9 ) );
  OR2_X2 \regfile/C1395  ( .A1(rs2_addr[2]), .A2(\regfile/N265 ), .ZN(
        \regfile/N266 ) );
  OR2_X2 \regfile/C1424  ( .A1(\regfile/N290 ), .A2(\regfile/N292 ), .ZN(
        \regfile/N293 ) );
  OR2_X2 \regfile/C1432  ( .A1(\regfile/N290 ), .A2(\regfile/N298 ), .ZN(
        \regfile/N299 ) );
  OR2_X2 \regfile/C1449  ( .A1(\regfile/N290 ), .A2(\regfile/N310 ), .ZN(
        \regfile/N311 ) );
  INV_X2 \regfile/I_12  ( .A(rd_addr[3]), .ZN(\regfile/N315 ) );
  OR2_X2 \regfile/C1489  ( .A1(\regfile/N290 ), .A2(\regfile/N341 ), .ZN(
        \regfile/N342 ) );
  OR2_X2 \regfile/C1517  ( .A1(\regfile/N290 ), .A2(\regfile/N359 ), .ZN(
        \regfile/N360 ) );
  OR2_X2 \regfile/C1557  ( .A1(\regfile/N290 ), .A2(\regfile/N390 ), .ZN(
        \regfile/N391 ) );
  OR2_X2 \regfile/C1566  ( .A1(\regfile/N290 ), .A2(\regfile/N396 ), .ZN(
        \regfile/N397 ) );
  OR2_X2 \regfile/C1585  ( .A1(\regfile/N290 ), .A2(\regfile/N402 ), .ZN(
        \regfile/N409 ) );
  INV_X2 \Scc_coproc/I_16  ( .A(\Scc_coproc/interrupt_active ), .ZN(
        \Scc_coproc/N551 ) );
  AND2_X2 \Scc_coproc/C954  ( .A1(\Scc_coproc/din_exc_word[4] ), .A2(
        \Scc_coproc/din_exc_word[5] ), .ZN(\Scc_coproc/N562 ) );
  AND2_X2 \Scc_coproc/C964  ( .A1(\Scc_coproc/ein_exc_word[4] ), .A2(
        \Scc_coproc/ein_exc_word[5] ), .ZN(\Scc_coproc/N571 ) );
  AND2_X2 \Scc_coproc/C965  ( .A1(\Scc_coproc/ein_exc_word[3] ), .A2(
        \Scc_coproc/N571 ), .ZN(\Scc_coproc/N572 ) );
  AND2_X2 \Scc_coproc/C966  ( .A1(\Scc_coproc/ein_exc_word[2] ), .A2(
        \Scc_coproc/N572 ), .ZN(\Scc_coproc/N573 ) );
  AND2_X2 \Scc_coproc/C967  ( .A1(\Scc_coproc/ein_exc_word[1] ), .A2(
        \Scc_coproc/N573 ), .ZN(\Scc_coproc/N574 ) );
  AND2_X2 \Scc_coproc/C968  ( .A1(\Scc_coproc/ein_exc_word[0] ), .A2(
        \Scc_coproc/N574 ), .ZN(\Scc_coproc/N575 ) );
  AND2_X2 \Scc_coproc/C970  ( .A1(\Scc_coproc/x_exc_word[3] ), .A2(
        \Scc_coproc/N576 ), .ZN(\Scc_coproc/N577 ) );
  AND2_X2 \Scc_coproc/C971  ( .A1(\Scc_coproc/x_exc_word[2] ), .A2(
        \Scc_coproc/N577 ), .ZN(\Scc_coproc/N578 ) );
  AND2_X2 \Scc_coproc/C972  ( .A1(\Scc_coproc/x_exc_word[1] ), .A2(
        \Scc_coproc/N578 ), .ZN(\Scc_coproc/N579 ) );
  OR2_X2 \Scc_coproc/C975  ( .A1(\Scc_coproc/interrupt[8] ), .A2(
        \Scc_coproc/interrupt[9] ), .ZN(\Scc_coproc/N582 ) );
  OR2_X2 \Scc_coproc/C976  ( .A1(\Scc_coproc/interrupt[7] ), .A2(
        \Scc_coproc/N582 ), .ZN(\Scc_coproc/N583 ) );
  OR2_X2 \Scc_coproc/C977  ( .A1(\Scc_coproc/interrupt[6] ), .A2(
        \Scc_coproc/N583 ), .ZN(\Scc_coproc/N584 ) );
  OR2_X2 \Scc_coproc/C978  ( .A1(\Scc_coproc/interrupt[5] ), .A2(
        \Scc_coproc/N584 ), .ZN(\Scc_coproc/N585 ) );
  OR2_X2 \Scc_coproc/C979  ( .A1(\Scc_coproc/interrupt[4] ), .A2(
        \Scc_coproc/N585 ), .ZN(\Scc_coproc/N586 ) );
  OR2_X2 \Scc_coproc/C980  ( .A1(\Scc_coproc/interrupt[3] ), .A2(
        \Scc_coproc/N586 ), .ZN(\Scc_coproc/N587 ) );
  OR2_X2 \Scc_coproc/C995  ( .A1(\Scc_coproc/mem_cop_op [1]), .A2(
        \Scc_coproc/N599 ), .ZN(\Scc_coproc/N600 ) );
  OR2_X2 \Scc_coproc/C996  ( .A1(\Scc_coproc/mem_cop_op [0]), .A2(
        \Scc_coproc/N600 ), .ZN(\Scc_coproc/N601 ) );
  AND2_X2 \Scc_coproc/C1247  ( .A1(INTERRUPT_VECTOR[0]), .A2(
        \Scc_coproc/status[2] ), .ZN(\Scc_coproc/interrupt[2] ) );
  OR2_X2 C209 ( .A1(N82), .A2(N83), .ZN(N80) );
  OR2_X2 C205 ( .A1(N82), .A2(N83), .ZN(N5) );
  INV_X2 I_5 ( .A(\x_mem_command[MW] ), .ZN(N83) );
  INV_X2 I_4 ( .A(\x_mem_command[MR] ), .ZN(N82) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_e/data_out_reg[0]  ( .D(n4504), .CK(CLK), 
        .SN(n7825), .QN(n3107) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_m/data_out_reg[0]  ( .D(n4501), .CK(CLK), 
        .SN(n7825), .Q(\Scc_coproc/mem_cop_op [0]), .QN(n3104) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_m/data_out_reg[1]  ( .D(n4500), .CK(CLK), 
        .SN(n7825), .Q(\Scc_coproc/mem_cop_op [1]), .QN(n3103) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_m/data_out_reg[2]  ( .D(n4499), .CK(CLK), 
        .SN(n7825), .Q(\Scc_coproc/N599 ), .QN(n3102) );
  DFFR_X1 \Mpath/regMaddr/data_out_reg[1]  ( .D(n4498), .CK(CLK), .RN(n7750), 
        .Q(\Mpath/mem_baddr [1]), .QN(\Mpath/the_memhandle/N239 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[0]  ( .D(n4497), .CK(CLK), .RN(n7745), .Q(
        \Mpath/out_regB[0] ), .QN(\Mpath/the_alu/N84 ) );
  DFFR_X1 \Mpath/regMaddr/data_out_reg[0]  ( .D(n4496), .CK(CLK), .RN(n7751), 
        .Q(\Mpath/mem_baddr [0]), .QN(\Mpath/the_memhandle/N240 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[0]  ( .D(n4495), .CK(CLK), .RN(n7751), .QN(
        n5620) );
  DFFR_X1 \Mpath/regM/data_out_reg[31]  ( .D(n4493), .CK(CLK), .RN(n7753), 
        .QN(n5548) );
  DFFR_X1 \Mpath/regB/data_out_reg[31]  ( .D(n4492), .CK(CLK), .RN(n7769), .Q(
        \Mpath/out_regB[31] ), .QN(\Mpath/the_alu/N22 ) );
  DFFR_X1 \Scc_coproc/CAUSE_REG/data_out_reg[0]  ( .D(n4491), .CK(CLK), .RN(
        n7784), .QN(n6489) );
  DFFR_X1 \Mpath/JAR/data_out_reg[1]  ( .D(n4487), .CK(CLK), .RN(n7753), .QN(
        n6087) );
  DFFR_X1 \Mpath/JAR/data_out_reg[2]  ( .D(n4486), .CK(CLK), .RN(n7753), .QN(
        n6209) );
  DFFR_X1 \Mpath/JAR/data_out_reg[3]  ( .D(n4485), .CK(CLK), .RN(n7720), .QN(
        n6194) );
  DFFR_X1 \Mpath/JAR/data_out_reg[4]  ( .D(n4484), .CK(CLK), .RN(n7720), .QN(
        n6180) );
  DFFR_X1 \Mpath/JAR/data_out_reg[5]  ( .D(n4483), .CK(CLK), .RN(n7741), .QN(
        n6163) );
  DFFR_X1 \Mpath/JAR/data_out_reg[6]  ( .D(n4482), .CK(CLK), .RN(n7740), .QN(
        n6151) );
  DFFR_X1 \Mpath/JAR/data_out_reg[7]  ( .D(n4481), .CK(CLK), .RN(n7741), .QN(
        n6139) );
  DFFR_X1 \Mpath/JAR/data_out_reg[8]  ( .D(n4480), .CK(CLK), .RN(n7752), .QN(
        n6127) );
  DFFR_X1 \Mpath/JAR/data_out_reg[9]  ( .D(n4479), .CK(CLK), .RN(n7812), .QN(
        n6114) );
  DFFR_X1 \Mpath/JAR/data_out_reg[10]  ( .D(n4478), .CK(CLK), .RN(n7782), .QN(
        n6391) );
  DFFR_X1 \Mpath/JAR/data_out_reg[11]  ( .D(n4477), .CK(CLK), .RN(n7737), .QN(
        n6377) );
  DFFR_X1 \Mpath/JAR/data_out_reg[12]  ( .D(n4476), .CK(CLK), .RN(n7782), .QN(
        n6365) );
  DFFR_X1 \Mpath/JAR/data_out_reg[13]  ( .D(n4475), .CK(CLK), .RN(n7752), .QN(
        n6353) );
  DFFR_X1 \Mpath/JAR/data_out_reg[14]  ( .D(n4474), .CK(CLK), .RN(n7772), .QN(
        n6341) );
  DFFR_X1 \Mpath/JAR/data_out_reg[15]  ( .D(n4473), .CK(CLK), .RN(n7779), .QN(
        n6329) );
  DFFR_X1 \Mpath/JAR/data_out_reg[16]  ( .D(n4472), .CK(CLK), .RN(n7773), .QN(
        n6317) );
  DFFR_X1 \Mpath/JAR/data_out_reg[17]  ( .D(n4471), .CK(CLK), .RN(n7752), .QN(
        n6305) );
  DFFR_X1 \Mpath/JAR/data_out_reg[18]  ( .D(n4470), .CK(CLK), .RN(n7773), .QN(
        n6291) );
  DFFR_X1 \Mpath/JAR/data_out_reg[19]  ( .D(n4469), .CK(CLK), .RN(n7734), .QN(
        n6276) );
  DFFR_X1 \Mpath/JAR/data_out_reg[20]  ( .D(n4468), .CK(CLK), .RN(n7773), .QN(
        n6263) );
  DFFR_X1 \Mpath/JAR/data_out_reg[21]  ( .D(n4467), .CK(CLK), .RN(n7751), .QN(
        n6247) );
  DFFR_X1 \Mpath/JAR/data_out_reg[22]  ( .D(n4466), .CK(CLK), .RN(n7773), .QN(
        n6235) );
  DFFR_X1 \Mpath/JAR/data_out_reg[23]  ( .D(n4465), .CK(CLK), .RN(n7754), .QN(
        n6223) );
  DFFR_X1 \Mpath/regM/data_out_reg[23]  ( .D(n4464), .CK(CLK), .RN(n7754), 
        .QN(n5575) );
  DFFR_X1 \Mpath/regB/data_out_reg[23]  ( .D(n4463), .CK(CLK), .RN(n7766), .Q(
        \Mpath/out_regB[23] ), .QN(\Mpath/the_alu/N38 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[30]  ( .D(n4462), .CK(CLK), .RN(n7751), 
        .QN(n5551) );
  DFFR_X1 \Mpath/regM/data_out_reg[29]  ( .D(n4460), .CK(CLK), .RN(n7717), 
        .QN(n5557) );
  DFFR_X1 \Mpath/regM/data_out_reg[28]  ( .D(n4458), .CK(CLK), .RN(n7806), 
        .QN(n5560) );
  DFFR_X1 \Mpath/regM/data_out_reg[27]  ( .D(n4456), .CK(CLK), .RN(n7809), 
        .QN(n5563) );
  DFFR_X1 \Mpath/regM/data_out_reg[26]  ( .D(n4454), .CK(CLK), .RN(n7817), 
        .QN(n5566) );
  DFFR_X1 \Mpath/regM/data_out_reg[14]  ( .D(n4452), .CK(CLK), .RN(n7772), 
        .QN(n5605) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[14]  ( .D(n4451), .CK(CLK), .RN(
        n7756), .QN(n5739) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[14]  ( .D(n4450), .CK(CLK), .SN(
        n7825), .QN(n5740) );
  DFFR_X1 \Mpath/regM/data_out_reg[8]  ( .D(n4448), .CK(CLK), .RN(n7752), .QN(
        n5530) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[8]  ( .D(n4447), .CK(CLK), .RN(
        n7755), .QN(n5724) );
  DFFR_X1 \Scc_coproc/STATUS_REG/data_out_reg[8]  ( .D(n4446), .CK(CLK), .RN(
        n7755), .QN(n5723) );
  DFFR_X1 \Mpath/regM/data_out_reg[4]  ( .D(n4443), .CK(CLK), .RN(n7720), .QN(
        n5542) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[4]  ( .D(n4442), .CK(CLK), .RN(
        n7755), .QN(n5732) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[4]  ( .D(n4441), .CK(CLK), .SN(
        n7825), .QN(n5731) );
  DFFR_X1 \Scc_coproc/CAUSE_REG/data_out_reg[3]  ( .D(n4439), .CK(CLK), .RN(
        n7784), .QN(n6482) );
  DFFR_X1 \Mpath/regM/data_out_reg[3]  ( .D(n4438), .CK(CLK), .RN(n7803), .QN(
        n5545) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[3]  ( .D(n4437), .CK(CLK), .RN(
        n7755), .QN(n5734) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[3]  ( .D(n4436), .CK(CLK), .SN(
        n7824), .QN(n5733) );
  DFFR_X1 \Scc_coproc/CAUSE_REG/data_out_reg[2]  ( .D(n4434), .CK(CLK), .RN(
        n7783), .QN(n6484) );
  DFFR_X1 \Mpath/regM/data_out_reg[2]  ( .D(n4433), .CK(CLK), .RN(n7753), .QN(
        n5554) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[2]  ( .D(n4432), .CK(CLK), .RN(
        n7755), .QN(n5736) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[2]  ( .D(n4431), .CK(CLK), .SN(
        n7824), .Q(\Scc_coproc/status[2] ), .QN(n5735) );
  DFFR_X1 \Mpath/regM/data_out_reg[1]  ( .D(n4429), .CK(CLK), .RN(n7723), .QN(
        n5587) );
  DFFR_X1 \Mpath/regB/data_out_reg[1]  ( .D(n4428), .CK(CLK), .RN(n7720), .Q(
        \Mpath/out_regB[1] ), .QN(\Mpath/the_alu/N82 ) );
  DFFS_X1 \Mcontrol/ir_xm/out_rf_we_reg  ( .D(n4422), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(m_we), .QN(\Mcontrol/bp_logicA/N14 ) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[31]  ( .D(n4421), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [31]), .QN(n7653)
         );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[30]  ( .D(n4420), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [30]), .QN(n7150)
         );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[29]  ( .D(n4419), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [29]), .QN(n7631)
         );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[28]  ( .D(n4418), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .QN(n3087) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[27]  ( .D(n4417), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [27]), .QN(n3086)
         );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[26]  ( .D(n4416), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [26]), .QN(n3085)
         );
  DFFS_X1 \Mcontrol/ir_xm/out_mem_command_reg[SIGN]  ( .D(n4414), .CK(CLK), 
        .SN(\Mcontrol/int_reset ), .Q(\m_mem_command[SIGN] ), .QN(
        \Mpath/the_memhandle/N235 ) );
  DFFS_X1 \Mcontrol/ir_xm/out_mem_command_reg[MH]  ( .D(n4409), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(\Mpath/the_memhandle/N238 ) );
  DFFS_X1 \Mcontrol/ir_xm/out_mem_command_reg[MB]  ( .D(n4407), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(\Mpath/the_memhandle/N236 ) );
  DFFS_X1 \Mcontrol/ir_xm/out_alu_command_reg[HRDWIT]  ( .D(n4405), .CK(CLK), 
        .SN(\Mcontrol/int_reset ), .QN(\Mcontrol/N17 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_exe_outsel1_reg[2]  ( .D(n4404), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(exe_outsel[2]), .QN(\Mpath/N179 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_exe_outsel1_reg[1]  ( .D(n4403), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(exe_outsel[1]), .QN(\Mpath/N187 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_exe_outsel1_reg[0]  ( .D(n4402), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(exe_outsel[0]), .QN(\Mpath/N180 ) );
  DFFR_X1 \Mcontrol/bvgen/jtype_reg1/data_out_reg[4]  ( .D(n4395), .CK(CLK), 
        .RN(n7754), .Q(\Mcontrol/bvgen/N6 ), .QN(n3072) );
  DFFR_X1 \Mcontrol/bvgen/jtype_reg1/data_out_reg[3]  ( .D(n4393), .CK(CLK), 
        .RN(n7754), .QN(\Mcontrol/bvgen/N2 ) );
  DFFR_X1 \Mcontrol/bvgen/jtype_reg1/data_out_reg[1]  ( .D(n4390), .CK(CLK), 
        .RN(n7754), .QN(\Mcontrol/bvgen/N4 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_mul_command_reg[5]  ( .D(n4377), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_mul_command [5]), .QN(n3056) );
  DFFR_X1 \Mcontrol/ir_dx/out_alu_command_reg[OP][5]  ( .D(n4376), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][5] ), .QN(
        \Mpath/the_alu/N466 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_mul_command_reg[4]  ( .D(n4374), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_mul_command [4]), .QN(n3054) );
  DFFR_X1 \Mcontrol/ir_dx/out_alu_command_reg[OP][4]  ( .D(n4373), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][4] ), .QN(
        \Mpath/the_alu/N453 ) );
  DFFS_X1 \Mcontrol/ir_dx/out_mul_command_reg[2]  ( .D(n4368), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(\Mcontrol/st_logic/N26 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_shift_op1_reg[2]  ( .D(n4367), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(shift_op[2]), .QN(\Mpath/the_shift/N104 ) );
  DFFS_X1 \Mcontrol/ir_dx/out_mul_command_reg[1]  ( .D(n4364), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(\Mcontrol/st_logic/N27 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_shift_op1_reg[1]  ( .D(n4363), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(shift_op[1]), .QN(\Mpath/the_shift/N112 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_alu_command_reg[OP][1]  ( .D(n4362), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][1] ), .QN(
        \Mpath/the_alu/N467 ) );
  DFFS_X1 \Mcontrol/ir_dx/out_mul_command_reg[0]  ( .D(n4360), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_mul_command [0]), .QN(
        \Mcontrol/st_logic/N34 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_shift_op1_reg[0]  ( .D(n4359), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(shift_op[0]), .QN(\Mpath/the_shift/N105 ) );
  DFFR_X1 \Mcontrol/ir_dx/out_alu_command_reg[OP][0]  ( .D(n4358), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][0] ), .QN(
        \Mpath/the_alu/N468 ) );
  DFFR_X1 \Mcontrol/ir_xm/out_rd1_reg[4]  ( .D(n4356), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/m_sampled_xrd[4] ), .QN(n3045) );
  DFFR_X1 \Mcontrol/ir_xm/out_rd1_reg[3]  ( .D(n4354), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/m_sampled_xrd[3] ), .QN(n3043) );
  DFFR_X1 \Mcontrol/ir_xm/out_rd1_reg[2]  ( .D(n4352), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/m_sampled_xrd[2] ), .QN(n3041) );
  DFFR_X1 \Mcontrol/ir_xm/out_rd1_reg[1]  ( .D(n4350), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/m_sampled_xrd[1] ), .QN(n3039) );
  DFFR_X1 \regfile/rx_5/data_out_reg[0]  ( .D(n4319), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[5][0] ), .QN(n4670) );
  DFFR_X1 \regfile/rx_5/data_out_reg[14]  ( .D(n4318), .CK(CLK), .RN(n7772), 
        .Q(\regfile/reg_out[5][14] ), .QN(n4665) );
  DFFR_X1 \regfile/rx_5/data_out_reg[1]  ( .D(n4317), .CK(CLK), .RN(n7723), 
        .Q(\regfile/reg_out[5][1] ), .QN(n4659) );
  DFFR_X1 \regfile/rx_5/data_out_reg[23]  ( .D(n4316), .CK(CLK), .RN(n7769), 
        .Q(\regfile/reg_out[5][23] ), .QN(n4655) );
  DFFR_X1 \regfile/rx_5/data_out_reg[26]  ( .D(n4315), .CK(CLK), .RN(n7817), 
        .Q(\regfile/reg_out[5][26] ), .QN(n4652) );
  DFFR_X1 \regfile/rx_5/data_out_reg[27]  ( .D(n4314), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[5][27] ), .QN(n4651) );
  DFFR_X1 \regfile/rx_5/data_out_reg[28]  ( .D(n4313), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[5][28] ), .QN(n4650) );
  DFFR_X1 \regfile/rx_5/data_out_reg[29]  ( .D(n4312), .CK(CLK), .RN(n7717), 
        .Q(\regfile/reg_out[5][29] ), .QN(n4649) );
  DFFR_X1 \regfile/rx_5/data_out_reg[2]  ( .D(n4311), .CK(CLK), .RN(n7750), 
        .Q(\regfile/reg_out[5][2] ), .QN(n4648) );
  DFFR_X1 \regfile/rx_5/data_out_reg[30]  ( .D(n4310), .CK(CLK), .RN(n7766), 
        .Q(\regfile/reg_out[5][30] ), .QN(n4647) );
  DFFR_X1 \regfile/rx_5/data_out_reg[3]  ( .D(n4308), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[5][3] ), .QN(n4645) );
  DFFR_X1 \regfile/rx_5/data_out_reg[4]  ( .D(n4307), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[5][4] ), .QN(n4644) );
  DFFR_X1 \regfile/rx_5/data_out_reg[8]  ( .D(n4306), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[5][8] ), .QN(n4640) );
  DFFR_X1 \regfile/rx_19/data_out_reg[0]  ( .D(n4221), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[19][0] ), .QN(n5214) );
  DFFR_X1 \regfile/rx_19/data_out_reg[14]  ( .D(n4220), .CK(CLK), .RN(n7772), 
        .Q(\regfile/reg_out[19][14] ), .QN(n5209) );
  DFFR_X1 \regfile/rx_19/data_out_reg[1]  ( .D(n4219), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[19][1] ), .QN(n5203) );
  DFFR_X1 \regfile/rx_19/data_out_reg[23]  ( .D(n4218), .CK(CLK), .RN(n7768), 
        .Q(\regfile/reg_out[19][23] ), .QN(n5199) );
  DFFR_X1 \regfile/rx_19/data_out_reg[26]  ( .D(n4217), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[19][26] ), .QN(n5196) );
  DFFR_X1 \regfile/rx_19/data_out_reg[27]  ( .D(n4216), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[19][27] ), .QN(n5195) );
  DFFR_X1 \regfile/rx_19/data_out_reg[28]  ( .D(n4215), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[19][28] ), .QN(n5194) );
  DFFR_X1 \regfile/rx_19/data_out_reg[29]  ( .D(n4214), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[19][29] ), .QN(n5193) );
  DFFR_X1 \regfile/rx_19/data_out_reg[2]  ( .D(n4213), .CK(CLK), .RN(n7750), 
        .Q(\regfile/reg_out[19][2] ), .QN(n5192) );
  DFFR_X1 \regfile/rx_19/data_out_reg[30]  ( .D(n4212), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[19][30] ), .QN(n5191) );
  DFFR_X1 \regfile/rx_19/data_out_reg[3]  ( .D(n4210), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[19][3] ), .QN(n5189) );
  DFFR_X1 \regfile/rx_19/data_out_reg[4]  ( .D(n4209), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[19][4] ), .QN(n5188) );
  DFFR_X1 \regfile/rx_19/data_out_reg[8]  ( .D(n4208), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[19][8] ), .QN(n5184) );
  DFFR_X1 \regfile/rx_21/data_out_reg[0]  ( .D(n4207), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[21][0] ), .QN(n5118) );
  DFFR_X1 \regfile/rx_21/data_out_reg[14]  ( .D(n4206), .CK(CLK), .RN(n7771), 
        .Q(\regfile/reg_out[21][14] ), .QN(n5113) );
  DFFR_X1 \regfile/rx_21/data_out_reg[1]  ( .D(n4205), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[21][1] ), .QN(n5107) );
  DFFR_X1 \regfile/rx_21/data_out_reg[23]  ( .D(n4204), .CK(CLK), .RN(n7768), 
        .Q(\regfile/reg_out[21][23] ), .QN(n5103) );
  DFFR_X1 \regfile/rx_21/data_out_reg[26]  ( .D(n4203), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[21][26] ), .QN(n5100) );
  DFFR_X1 \regfile/rx_21/data_out_reg[27]  ( .D(n4202), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[21][27] ), .QN(n5099) );
  DFFR_X1 \regfile/rx_21/data_out_reg[28]  ( .D(n4201), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[21][28] ), .QN(n5098) );
  DFFR_X1 \regfile/rx_21/data_out_reg[29]  ( .D(n4200), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[21][29] ), .QN(n5097) );
  DFFR_X1 \regfile/rx_21/data_out_reg[2]  ( .D(n4199), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[21][2] ), .QN(n5096) );
  DFFR_X1 \regfile/rx_21/data_out_reg[30]  ( .D(n4198), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[21][30] ), .QN(n5095) );
  DFFR_X1 \regfile/rx_21/data_out_reg[3]  ( .D(n4196), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[21][3] ), .QN(n5093) );
  DFFR_X1 \regfile/rx_21/data_out_reg[4]  ( .D(n4195), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[21][4] ), .QN(n5092) );
  DFFR_X1 \regfile/rx_21/data_out_reg[8]  ( .D(n4194), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[21][8] ), .QN(n5088) );
  DFFR_X1 \regfile/rx_25/data_out_reg[0]  ( .D(n4179), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[25][0] ), .QN(n4990) );
  DFFR_X1 \regfile/rx_25/data_out_reg[14]  ( .D(n4178), .CK(CLK), .RN(n7771), 
        .Q(\regfile/reg_out[25][14] ), .QN(n4985) );
  DFFR_X1 \regfile/rx_25/data_out_reg[1]  ( .D(n4177), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[25][1] ), .QN(n4979) );
  DFFR_X1 \regfile/rx_25/data_out_reg[23]  ( .D(n4176), .CK(CLK), .RN(n7768), 
        .Q(\regfile/reg_out[25][23] ), .QN(n4975) );
  DFFR_X1 \regfile/rx_25/data_out_reg[26]  ( .D(n4175), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[25][26] ), .QN(n4972) );
  DFFR_X1 \regfile/rx_25/data_out_reg[27]  ( .D(n4174), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[25][27] ), .QN(n4971) );
  DFFR_X1 \regfile/rx_25/data_out_reg[28]  ( .D(n4173), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[25][28] ), .QN(n4970) );
  DFFR_X1 \regfile/rx_25/data_out_reg[29]  ( .D(n4172), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[25][29] ), .QN(n4969) );
  DFFR_X1 \regfile/rx_25/data_out_reg[2]  ( .D(n4171), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[25][2] ), .QN(n4968) );
  DFFR_X1 \regfile/rx_25/data_out_reg[30]  ( .D(n4170), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[25][30] ), .QN(n4967) );
  DFFR_X1 \regfile/rx_25/data_out_reg[3]  ( .D(n4168), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[25][3] ), .QN(n4965) );
  DFFR_X1 \regfile/rx_25/data_out_reg[4]  ( .D(n4167), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[25][4] ), .QN(n4964) );
  DFFR_X1 \regfile/rx_25/data_out_reg[8]  ( .D(n4166), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[25][8] ), .QN(n4960) );
  DFFR_X1 \regfile/rx_29/data_out_reg[0]  ( .D(n4151), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[29][0] ), .QN(n4862) );
  DFFR_X1 \regfile/rx_29/data_out_reg[14]  ( .D(n4150), .CK(CLK), .RN(n7771), 
        .Q(\regfile/reg_out[29][14] ), .QN(n4857) );
  DFFR_X1 \regfile/rx_29/data_out_reg[1]  ( .D(n4149), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[29][1] ), .QN(n4851) );
  DFFR_X1 \regfile/rx_29/data_out_reg[23]  ( .D(n4148), .CK(CLK), .RN(n7768), 
        .Q(\regfile/reg_out[29][23] ), .QN(n4847) );
  DFFR_X1 \regfile/rx_29/data_out_reg[26]  ( .D(n4147), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[29][26] ), .QN(n4844) );
  DFFR_X1 \regfile/rx_29/data_out_reg[27]  ( .D(n4146), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[29][27] ), .QN(n4843) );
  DFFR_X1 \regfile/rx_29/data_out_reg[28]  ( .D(n4145), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[29][28] ), .QN(n4842) );
  DFFR_X1 \regfile/rx_29/data_out_reg[29]  ( .D(n4144), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[29][29] ), .QN(n4841) );
  DFFR_X1 \regfile/rx_29/data_out_reg[2]  ( .D(n4143), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[29][2] ), .QN(n4840) );
  DFFR_X1 \regfile/rx_29/data_out_reg[30]  ( .D(n4142), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[29][30] ), .QN(n4839) );
  DFFR_X1 \regfile/rx_29/data_out_reg[3]  ( .D(n4140), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[29][3] ), .QN(n4837) );
  DFFR_X1 \regfile/rx_29/data_out_reg[4]  ( .D(n4139), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[29][4] ), .QN(n4836) );
  DFFR_X1 \regfile/rx_29/data_out_reg[8]  ( .D(n4138), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[29][8] ), .QN(n4832) );
  DFFR_X1 \regfile/rx_4/data_out_reg[0]  ( .D(n4109), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[4][0] ), .QN(n4702) );
  DFFR_X1 \regfile/rx_4/data_out_reg[14]  ( .D(n4108), .CK(CLK), .RN(n7771), 
        .Q(\regfile/reg_out[4][14] ), .QN(n4697) );
  DFFR_X1 \regfile/rx_4/data_out_reg[1]  ( .D(n4107), .CK(CLK), .RN(n7721), 
        .Q(\regfile/reg_out[4][1] ), .QN(n4691) );
  DFFR_X1 \regfile/rx_4/data_out_reg[23]  ( .D(n4106), .CK(CLK), .RN(n7767), 
        .Q(\regfile/reg_out[4][23] ), .QN(n4687) );
  DFFR_X1 \regfile/rx_4/data_out_reg[26]  ( .D(n4105), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[4][26] ), .QN(n4684) );
  DFFR_X1 \regfile/rx_4/data_out_reg[27]  ( .D(n4104), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[4][27] ), .QN(n4683) );
  DFFR_X1 \regfile/rx_4/data_out_reg[28]  ( .D(n4103), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[4][28] ), .QN(n4682) );
  DFFR_X1 \regfile/rx_4/data_out_reg[29]  ( .D(n4102), .CK(CLK), .RN(n7742), 
        .Q(\regfile/reg_out[4][29] ), .QN(n4681) );
  DFFR_X1 \regfile/rx_4/data_out_reg[2]  ( .D(n4101), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[4][2] ), .QN(n4680) );
  DFFR_X1 \regfile/rx_4/data_out_reg[30]  ( .D(n4100), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[4][30] ), .QN(n4679) );
  DFFR_X1 \regfile/rx_4/data_out_reg[3]  ( .D(n4098), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[4][3] ), .QN(n4677) );
  DFFR_X1 \regfile/rx_4/data_out_reg[4]  ( .D(n4097), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[4][4] ), .QN(n4676) );
  DFFR_X1 \regfile/rx_4/data_out_reg[8]  ( .D(n4096), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[4][8] ), .QN(n4672) );
  DFFR_X1 \regfile/rx_18/data_out_reg[0]  ( .D(n4011), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[18][0] ), .QN(n5246) );
  DFFR_X1 \regfile/rx_18/data_out_reg[14]  ( .D(n4010), .CK(CLK), .RN(n7770), 
        .Q(\regfile/reg_out[18][14] ), .QN(n5241) );
  DFFR_X1 \regfile/rx_18/data_out_reg[1]  ( .D(n4009), .CK(CLK), .RN(n7721), 
        .Q(\regfile/reg_out[18][1] ), .QN(n5235) );
  DFFR_X1 \regfile/rx_18/data_out_reg[23]  ( .D(n4008), .CK(CLK), .RN(n7767), 
        .Q(\regfile/reg_out[18][23] ), .QN(n5231) );
  DFFR_X1 \regfile/rx_18/data_out_reg[26]  ( .D(n4007), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[18][26] ), .QN(n5228) );
  DFFR_X1 \regfile/rx_18/data_out_reg[27]  ( .D(n4006), .CK(CLK), .RN(n7806), 
        .Q(\regfile/reg_out[18][27] ), .QN(n5227) );
  DFFR_X1 \regfile/rx_18/data_out_reg[28]  ( .D(n4005), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[18][28] ), .QN(n5226) );
  DFFR_X1 \regfile/rx_18/data_out_reg[29]  ( .D(n4004), .CK(CLK), .RN(n7741), 
        .Q(\regfile/reg_out[18][29] ), .QN(n5225) );
  DFFR_X1 \regfile/rx_18/data_out_reg[2]  ( .D(n4003), .CK(CLK), .RN(n7748), 
        .Q(\regfile/reg_out[18][2] ), .QN(n5224) );
  DFFR_X1 \regfile/rx_18/data_out_reg[30]  ( .D(n4002), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[18][30] ), .QN(n5223) );
  DFFR_X1 \regfile/rx_18/data_out_reg[3]  ( .D(n4000), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[18][3] ), .QN(n5221) );
  DFFR_X1 \regfile/rx_18/data_out_reg[4]  ( .D(n3999), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[18][4] ), .QN(n5220) );
  DFFR_X1 \regfile/rx_18/data_out_reg[8]  ( .D(n3998), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[18][8] ), .QN(n5216) );
  DFFR_X1 \regfile/rx_20/data_out_reg[0]  ( .D(n3997), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[20][0] ), .QN(n5150) );
  DFFR_X1 \regfile/rx_20/data_out_reg[14]  ( .D(n3996), .CK(CLK), .RN(n7770), 
        .Q(\regfile/reg_out[20][14] ), .QN(n5145) );
  DFFR_X1 \regfile/rx_20/data_out_reg[1]  ( .D(n3995), .CK(CLK), .RN(n7721), 
        .Q(\regfile/reg_out[20][1] ), .QN(n5139) );
  DFFR_X1 \regfile/rx_20/data_out_reg[23]  ( .D(n3994), .CK(CLK), .RN(n7767), 
        .Q(\regfile/reg_out[20][23] ), .QN(n5135) );
  DFFR_X1 \regfile/rx_20/data_out_reg[26]  ( .D(n3993), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[20][26] ), .QN(n5132) );
  DFFR_X1 \regfile/rx_20/data_out_reg[27]  ( .D(n3992), .CK(CLK), .RN(n7806), 
        .Q(\regfile/reg_out[20][27] ), .QN(n5131) );
  DFFR_X1 \regfile/rx_20/data_out_reg[28]  ( .D(n3991), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[20][28] ), .QN(n5130) );
  DFFR_X1 \regfile/rx_20/data_out_reg[29]  ( .D(n3990), .CK(CLK), .RN(n7741), 
        .Q(\regfile/reg_out[20][29] ), .QN(n5129) );
  DFFR_X1 \regfile/rx_20/data_out_reg[2]  ( .D(n3989), .CK(CLK), .RN(n7748), 
        .Q(\regfile/reg_out[20][2] ), .QN(n5128) );
  DFFR_X1 \regfile/rx_20/data_out_reg[30]  ( .D(n3988), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[20][30] ), .QN(n5127) );
  DFFR_X1 \regfile/rx_20/data_out_reg[3]  ( .D(n3986), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[20][3] ), .QN(n5125) );
  DFFR_X1 \regfile/rx_20/data_out_reg[4]  ( .D(n3985), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[20][4] ), .QN(n5124) );
  DFFR_X1 \regfile/rx_20/data_out_reg[8]  ( .D(n3984), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[20][8] ), .QN(n5120) );
  DFFR_X1 \regfile/rx_24/data_out_reg[0]  ( .D(n3969), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[24][0] ), .QN(n5022) );
  DFFR_X1 \regfile/rx_24/data_out_reg[14]  ( .D(n3968), .CK(CLK), .RN(n7770), 
        .Q(\regfile/reg_out[24][14] ), .QN(n5017) );
  DFFR_X1 \regfile/rx_24/data_out_reg[1]  ( .D(n3967), .CK(CLK), .RN(n7720), 
        .Q(\regfile/reg_out[24][1] ), .QN(n5011) );
  DFFR_X1 \regfile/rx_24/data_out_reg[23]  ( .D(n3966), .CK(CLK), .RN(n7766), 
        .Q(\regfile/reg_out[24][23] ), .QN(n5007) );
  DFFR_X1 \regfile/rx_24/data_out_reg[26]  ( .D(n3965), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[24][26] ), .QN(n5004) );
  DFFR_X1 \regfile/rx_24/data_out_reg[27]  ( .D(n3964), .CK(CLK), .RN(n7806), 
        .Q(\regfile/reg_out[24][27] ), .QN(n5003) );
  DFFR_X1 \regfile/rx_24/data_out_reg[28]  ( .D(n3963), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[24][28] ), .QN(n5002) );
  DFFR_X1 \regfile/rx_24/data_out_reg[29]  ( .D(n3962), .CK(CLK), .RN(n7741), 
        .Q(\regfile/reg_out[24][29] ), .QN(n5001) );
  DFFR_X1 \regfile/rx_24/data_out_reg[2]  ( .D(n3961), .CK(CLK), .RN(n7748), 
        .Q(\regfile/reg_out[24][2] ), .QN(n5000) );
  DFFR_X1 \regfile/rx_24/data_out_reg[30]  ( .D(n3960), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[24][30] ), .QN(n4999) );
  DFFR_X1 \regfile/rx_24/data_out_reg[3]  ( .D(n3958), .CK(CLK), .RN(n7800), 
        .Q(\regfile/reg_out[24][3] ), .QN(n4997) );
  DFFR_X1 \regfile/rx_24/data_out_reg[4]  ( .D(n3957), .CK(CLK), .RN(n7717), 
        .Q(\regfile/reg_out[24][4] ), .QN(n4996) );
  DFFR_X1 \regfile/rx_24/data_out_reg[8]  ( .D(n3956), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[24][8] ), .QN(n4992) );
  DFFR_X1 \regfile/rx_28/data_out_reg[0]  ( .D(n3941), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[28][0] ), .QN(n4894) );
  DFFR_X1 \regfile/rx_28/data_out_reg[14]  ( .D(n3940), .CK(CLK), .RN(n7770), 
        .Q(\regfile/reg_out[28][14] ), .QN(n4889) );
  DFFR_X1 \regfile/rx_28/data_out_reg[1]  ( .D(n3939), .CK(CLK), .RN(n7720), 
        .Q(\regfile/reg_out[28][1] ), .QN(n4883) );
  DFFR_X1 \regfile/rx_28/data_out_reg[23]  ( .D(n3938), .CK(CLK), .RN(n7766), 
        .Q(\regfile/reg_out[28][23] ), .QN(n4879) );
  DFFR_X1 \regfile/rx_28/data_out_reg[26]  ( .D(n3937), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[28][26] ), .QN(n4876) );
  DFFR_X1 \regfile/rx_28/data_out_reg[27]  ( .D(n3936), .CK(CLK), .RN(n7806), 
        .Q(\regfile/reg_out[28][27] ), .QN(n4875) );
  DFFR_X1 \regfile/rx_28/data_out_reg[28]  ( .D(n3935), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[28][28] ), .QN(n4874) );
  DFFR_X1 \regfile/rx_28/data_out_reg[29]  ( .D(n3934), .CK(CLK), .RN(n7741), 
        .Q(\regfile/reg_out[28][29] ), .QN(n4873) );
  DFFR_X1 \regfile/rx_28/data_out_reg[2]  ( .D(n3933), .CK(CLK), .RN(n7748), 
        .Q(\regfile/reg_out[28][2] ), .QN(n4872) );
  DFFR_X1 \regfile/rx_28/data_out_reg[30]  ( .D(n3932), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[28][30] ), .QN(n4871) );
  DFFR_X1 \regfile/rx_28/data_out_reg[3]  ( .D(n3930), .CK(CLK), .RN(n7800), 
        .Q(\regfile/reg_out[28][3] ), .QN(n4869) );
  DFFR_X1 \regfile/rx_28/data_out_reg[4]  ( .D(n3929), .CK(CLK), .RN(n7717), 
        .Q(\regfile/reg_out[28][4] ), .QN(n4868) );
  DFFR_X1 \regfile/rx_28/data_out_reg[8]  ( .D(n3928), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[28][8] ), .QN(n4864) );
  DFFR_X1 \Mcontrol/bvgen/jtype_reg1/data_out_reg[2]  ( .D(n3905), .CK(CLK), 
        .RN(n7754), .QN(\Mcontrol/bvgen/N3 ) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[5]  ( .D(n3895), .CK(CLK), .SN(
        n7823), .Q(\Scc_coproc/ein_exc_word[5] ), .QN(n3028) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[23]  ( .D(n3890), .CK(CLK), .RN(
        n7782), .QN(n6221) );
  DFFR_X1 \Mpath/regM/data_out_reg[9]  ( .D(n3883), .CK(CLK), .RN(n7811), .QN(
        n5526) );
  DFFR_X1 \regfile/rx_5/data_out_reg[9]  ( .D(n3878), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[5][9] ), .QN(n4639) );
  DFFR_X1 \regfile/rx_4/data_out_reg[9]  ( .D(n3877), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[4][9] ), .QN(n4671) );
  DFFR_X1 \regfile/rx_29/data_out_reg[9]  ( .D(n3872), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[29][9] ), .QN(n4831) );
  DFFR_X1 \regfile/rx_28/data_out_reg[9]  ( .D(n3871), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[28][9] ), .QN(n4863) );
  DFFR_X1 \regfile/rx_25/data_out_reg[9]  ( .D(n3868), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[25][9] ), .QN(n4959) );
  DFFR_X1 \regfile/rx_24/data_out_reg[9]  ( .D(n3867), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[24][9] ), .QN(n4991) );
  DFFR_X1 \regfile/rx_21/data_out_reg[9]  ( .D(n3864), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[21][9] ), .QN(n5087) );
  DFFR_X1 \regfile/rx_20/data_out_reg[9]  ( .D(n3863), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[20][9] ), .QN(n5119) );
  DFFR_X1 \regfile/rx_19/data_out_reg[9]  ( .D(n3861), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[19][9] ), .QN(n5183) );
  DFFR_X1 \regfile/rx_18/data_out_reg[9]  ( .D(n3860), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[18][9] ), .QN(n5215) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[9]  ( .D(n3850), .CK(CLK), .RN(
        n7755), .QN(n5722) );
  DFFR_X1 \Scc_coproc/STATUS_REG/data_out_reg[9]  ( .D(n3849), .CK(CLK), .RN(
        n7755), .QN(n5721) );
  DFFR_X1 \Mpath/regB/data_out_reg[9]  ( .D(n3847), .CK(CLK), .RN(n7782), .Q(
        \Mpath/out_regB[9] ), .QN(\Mpath/the_alu/N66 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[7]  ( .D(n3841), .CK(CLK), .RN(n7797), .QN(
        n5533) );
  DFFR_X1 \regfile/rx_5/data_out_reg[7]  ( .D(n3836), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[5][7] ), .QN(n4641) );
  DFFR_X1 \regfile/rx_4/data_out_reg[7]  ( .D(n3835), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[4][7] ), .QN(n4673) );
  DFFR_X1 \regfile/rx_29/data_out_reg[7]  ( .D(n3830), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[29][7] ), .QN(n4833) );
  DFFR_X1 \regfile/rx_28/data_out_reg[7]  ( .D(n3829), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[28][7] ), .QN(n4865) );
  DFFR_X1 \regfile/rx_25/data_out_reg[7]  ( .D(n3826), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[25][7] ), .QN(n4961) );
  DFFR_X1 \regfile/rx_24/data_out_reg[7]  ( .D(n3825), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[24][7] ), .QN(n4993) );
  DFFR_X1 \regfile/rx_21/data_out_reg[7]  ( .D(n3822), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[21][7] ), .QN(n5089) );
  DFFR_X1 \regfile/rx_20/data_out_reg[7]  ( .D(n3821), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[20][7] ), .QN(n5121) );
  DFFR_X1 \regfile/rx_19/data_out_reg[7]  ( .D(n3819), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[19][7] ), .QN(n5185) );
  DFFR_X1 \regfile/rx_18/data_out_reg[7]  ( .D(n3818), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[18][7] ), .QN(n5217) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[7]  ( .D(n3808), .CK(CLK), .RN(
        n7755), .QN(n5726) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[7]  ( .D(n3807), .CK(CLK), .SN(
        n7824), .QN(n5725) );
  DFFR_X1 \Mpath/regM/data_out_reg[6]  ( .D(n3799), .CK(CLK), .RN(n7740), .QN(
        n5536) );
  DFFR_X1 \regfile/rx_5/data_out_reg[6]  ( .D(n3794), .CK(CLK), .RN(n7740), 
        .Q(\regfile/reg_out[5][6] ), .QN(n4642) );
  DFFR_X1 \regfile/rx_4/data_out_reg[6]  ( .D(n3793), .CK(CLK), .RN(n7740), 
        .Q(\regfile/reg_out[4][6] ), .QN(n4674) );
  DFFR_X1 \regfile/rx_29/data_out_reg[6]  ( .D(n3788), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[29][6] ), .QN(n4834) );
  DFFR_X1 \regfile/rx_28/data_out_reg[6]  ( .D(n3787), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[28][6] ), .QN(n4866) );
  DFFR_X1 \regfile/rx_25/data_out_reg[6]  ( .D(n3784), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[25][6] ), .QN(n4962) );
  DFFR_X1 \regfile/rx_24/data_out_reg[6]  ( .D(n3783), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[24][6] ), .QN(n4994) );
  DFFR_X1 \regfile/rx_21/data_out_reg[6]  ( .D(n3780), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[21][6] ), .QN(n5090) );
  DFFR_X1 \regfile/rx_20/data_out_reg[6]  ( .D(n3779), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[20][6] ), .QN(n5122) );
  DFFR_X1 \regfile/rx_19/data_out_reg[6]  ( .D(n3777), .CK(CLK), .RN(n7739), 
        .Q(\regfile/reg_out[19][6] ), .QN(n5186) );
  DFFR_X1 \regfile/rx_18/data_out_reg[6]  ( .D(n3776), .CK(CLK), .RN(n7738), 
        .Q(\regfile/reg_out[18][6] ), .QN(n5218) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[6]  ( .D(n3766), .CK(CLK), .RN(
        n7755), .QN(n5728) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[6]  ( .D(n3765), .CK(CLK), .SN(
        n7823), .QN(n5727) );
  DFFR_X1 \Mpath/regM/data_out_reg[5]  ( .D(n3757), .CK(CLK), .RN(n7800), .QN(
        n5539) );
  DFFR_X1 \regfile/rx_5/data_out_reg[5]  ( .D(n3752), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[5][5] ), .QN(n4643) );
  DFFR_X1 \regfile/rx_4/data_out_reg[5]  ( .D(n3751), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[4][5] ), .QN(n4675) );
  DFFR_X1 \regfile/rx_29/data_out_reg[5]  ( .D(n3746), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[29][5] ), .QN(n4835) );
  DFFR_X1 \regfile/rx_28/data_out_reg[5]  ( .D(n3745), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[28][5] ), .QN(n4867) );
  DFFR_X1 \regfile/rx_25/data_out_reg[5]  ( .D(n3742), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[25][5] ), .QN(n4963) );
  DFFR_X1 \regfile/rx_24/data_out_reg[5]  ( .D(n3741), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[24][5] ), .QN(n4995) );
  DFFR_X1 \regfile/rx_21/data_out_reg[5]  ( .D(n3738), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[21][5] ), .QN(n5091) );
  DFFR_X1 \regfile/rx_20/data_out_reg[5]  ( .D(n3737), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[20][5] ), .QN(n5123) );
  DFFR_X1 \regfile/rx_19/data_out_reg[5]  ( .D(n3735), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[19][5] ), .QN(n5187) );
  DFFR_X1 \regfile/rx_18/data_out_reg[5]  ( .D(n3734), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[18][5] ), .QN(n5219) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[5]  ( .D(n3724), .CK(CLK), .RN(
        n7755), .QN(n5730) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[5]  ( .D(n3723), .CK(CLK), .SN(
        n7825), .QN(n5729) );
  DFFR_X1 \Scc_coproc/CAUSE_REG/data_out_reg[1]  ( .D(n3721), .CK(CLK), .RN(
        n7783), .QN(n6487) );
  DFFR_X1 \Mpath/regB/data_out_reg[5]  ( .D(n3720), .CK(CLK), .RN(n7797), .Q(
        \Mpath/out_regB[5] ), .QN(\Mpath/the_alu/N74 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[2]  ( .D(n3709), .CK(CLK), .RN(n7753), .Q(
        \Mpath/out_regB[2] ), .QN(\Mpath/the_alu/N80 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[3]  ( .D(n3703), .CK(CLK), .RN(n7800), .Q(
        \Mpath/out_regB[3] ), .QN(\Mpath/the_alu/N78 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[4]  ( .D(n3697), .CK(CLK), .RN(n7717), .Q(
        \Mpath/out_regB[4] ), .QN(\Mpath/the_alu/N76 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[8]  ( .D(n3691), .CK(CLK), .RN(n7752), .Q(
        \Mpath/out_regB[8] ), .QN(\Mpath/the_alu/N68 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[13]  ( .D(n3685), .CK(CLK), .RN(n7752), 
        .QN(n5608) );
  DFFR_X1 \regfile/rx_5/data_out_reg[13]  ( .D(n3680), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[5][13] ), .QN(n4666) );
  DFFR_X1 \regfile/rx_4/data_out_reg[13]  ( .D(n3679), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[4][13] ), .QN(n4698) );
  DFFR_X1 \regfile/rx_29/data_out_reg[13]  ( .D(n3674), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[29][13] ), .QN(n4858) );
  DFFR_X1 \regfile/rx_28/data_out_reg[13]  ( .D(n3673), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[28][13] ), .QN(n4890) );
  DFFR_X1 \regfile/rx_25/data_out_reg[13]  ( .D(n3670), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[25][13] ), .QN(n4986) );
  DFFR_X1 \regfile/rx_24/data_out_reg[13]  ( .D(n3669), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[24][13] ), .QN(n5018) );
  DFFR_X1 \regfile/rx_21/data_out_reg[13]  ( .D(n3666), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[21][13] ), .QN(n5114) );
  DFFR_X1 \regfile/rx_20/data_out_reg[13]  ( .D(n3665), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[20][13] ), .QN(n5146) );
  DFFR_X1 \regfile/rx_19/data_out_reg[13]  ( .D(n3663), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[19][13] ), .QN(n5210) );
  DFFR_X1 \regfile/rx_18/data_out_reg[13]  ( .D(n3662), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[18][13] ), .QN(n5242) );
  DFFR_X1 \Mpath/regM/data_out_reg[12]  ( .D(n3646), .CK(CLK), .RN(n7776), 
        .QN(n5611) );
  DFFR_X1 \regfile/rx_5/data_out_reg[12]  ( .D(n3641), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[5][12] ), .QN(n4667) );
  DFFR_X1 \regfile/rx_4/data_out_reg[12]  ( .D(n3640), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[4][12] ), .QN(n4699) );
  DFFR_X1 \regfile/rx_29/data_out_reg[12]  ( .D(n3635), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[29][12] ), .QN(n4859) );
  DFFR_X1 \regfile/rx_28/data_out_reg[12]  ( .D(n3634), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[28][12] ), .QN(n4891) );
  DFFR_X1 \regfile/rx_25/data_out_reg[12]  ( .D(n3631), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[25][12] ), .QN(n4987) );
  DFFR_X1 \regfile/rx_24/data_out_reg[12]  ( .D(n3630), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[24][12] ), .QN(n5019) );
  DFFR_X1 \regfile/rx_21/data_out_reg[12]  ( .D(n3627), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[21][12] ), .QN(n5115) );
  DFFR_X1 \regfile/rx_20/data_out_reg[12]  ( .D(n3626), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[20][12] ), .QN(n5147) );
  DFFR_X1 \regfile/rx_19/data_out_reg[12]  ( .D(n3624), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[19][12] ), .QN(n5211) );
  DFFR_X1 \regfile/rx_18/data_out_reg[12]  ( .D(n3623), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[18][12] ), .QN(n5243) );
  DFFR_X1 \Mpath/regM/data_out_reg[11]  ( .D(n3607), .CK(CLK), .RN(n7737), 
        .QN(n5614) );
  DFFR_X1 \regfile/rx_5/data_out_reg[11]  ( .D(n3602), .CK(CLK), .RN(n7737), 
        .Q(\regfile/reg_out[5][11] ), .QN(n4668) );
  DFFR_X1 \regfile/rx_4/data_out_reg[11]  ( .D(n3601), .CK(CLK), .RN(n7737), 
        .Q(\regfile/reg_out[4][11] ), .QN(n4700) );
  DFFR_X1 \regfile/rx_29/data_out_reg[11]  ( .D(n3596), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[29][11] ), .QN(n4860) );
  DFFR_X1 \regfile/rx_28/data_out_reg[11]  ( .D(n3595), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[28][11] ), .QN(n4892) );
  DFFR_X1 \regfile/rx_25/data_out_reg[11]  ( .D(n3592), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[25][11] ), .QN(n4988) );
  DFFR_X1 \regfile/rx_24/data_out_reg[11]  ( .D(n3591), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[24][11] ), .QN(n5020) );
  DFFR_X1 \regfile/rx_21/data_out_reg[11]  ( .D(n3588), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[21][11] ), .QN(n5116) );
  DFFR_X1 \regfile/rx_20/data_out_reg[11]  ( .D(n3587), .CK(CLK), .RN(n7736), 
        .Q(\regfile/reg_out[20][11] ), .QN(n5148) );
  DFFR_X1 \regfile/rx_19/data_out_reg[11]  ( .D(n3585), .CK(CLK), .RN(n7735), 
        .Q(\regfile/reg_out[19][11] ), .QN(n5212) );
  DFFR_X1 \regfile/rx_18/data_out_reg[11]  ( .D(n3584), .CK(CLK), .RN(n7735), 
        .Q(\regfile/reg_out[18][11] ), .QN(n5244) );
  DFFR_X1 \Mpath/regB/data_out_reg[11]  ( .D(n3574), .CK(CLK), .RN(n7734), .Q(
        \Mpath/out_regB[11] ), .QN(\Mpath/the_alu/N62 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[10]  ( .D(n3568), .CK(CLK), .RN(n7782), 
        .QN(n5617) );
  DFFR_X1 \regfile/rx_5/data_out_reg[10]  ( .D(n3563), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[5][10] ), .QN(n4669) );
  DFFR_X1 \regfile/rx_4/data_out_reg[10]  ( .D(n3562), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[4][10] ), .QN(n4701) );
  DFFR_X1 \regfile/rx_29/data_out_reg[10]  ( .D(n3557), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[29][10] ), .QN(n4861) );
  DFFR_X1 \regfile/rx_28/data_out_reg[10]  ( .D(n3556), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[28][10] ), .QN(n4893) );
  DFFR_X1 \regfile/rx_25/data_out_reg[10]  ( .D(n3553), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[25][10] ), .QN(n4989) );
  DFFR_X1 \regfile/rx_24/data_out_reg[10]  ( .D(n3552), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[24][10] ), .QN(n5021) );
  DFFR_X1 \regfile/rx_21/data_out_reg[10]  ( .D(n3549), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[21][10] ), .QN(n5117) );
  DFFR_X1 \regfile/rx_20/data_out_reg[10]  ( .D(n3548), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[20][10] ), .QN(n5149) );
  DFFR_X1 \regfile/rx_19/data_out_reg[10]  ( .D(n3546), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[19][10] ), .QN(n5213) );
  DFFR_X1 \regfile/rx_18/data_out_reg[10]  ( .D(n3545), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[18][10] ), .QN(n5245) );
  DFFR_X1 \Mpath/regB/data_out_reg[10]  ( .D(n3534), .CK(CLK), .RN(n7779), .Q(
        \Mpath/out_regB[10] ), .QN(\Mpath/the_alu/N64 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[14]  ( .D(n3533), .CK(CLK), .RN(n7790), .Q(
        \Mpath/out_regB[14] ), .QN(\Mpath/the_alu/N56 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[15]  ( .D(n3527), .CK(CLK), .RN(n7779), 
        .QN(n5602) );
  DFFR_X1 \regfile/rx_5/data_out_reg[15]  ( .D(n3522), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[5][15] ), .QN(n4664) );
  DFFR_X1 \regfile/rx_4/data_out_reg[15]  ( .D(n3521), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[4][15] ), .QN(n4696) );
  DFFR_X1 \regfile/rx_29/data_out_reg[15]  ( .D(n3516), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[29][15] ), .QN(n4856) );
  DFFR_X1 \regfile/rx_28/data_out_reg[15]  ( .D(n3515), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[28][15] ), .QN(n4888) );
  DFFR_X1 \regfile/rx_25/data_out_reg[15]  ( .D(n3512), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[25][15] ), .QN(n4984) );
  DFFR_X1 \regfile/rx_24/data_out_reg[15]  ( .D(n3511), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[24][15] ), .QN(n5016) );
  DFFR_X1 \regfile/rx_21/data_out_reg[15]  ( .D(n3508), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[21][15] ), .QN(n5112) );
  DFFR_X1 \regfile/rx_20/data_out_reg[15]  ( .D(n3507), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[20][15] ), .QN(n5144) );
  DFFR_X1 \regfile/rx_19/data_out_reg[15]  ( .D(n3505), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[19][15] ), .QN(n5208) );
  DFFR_X1 \regfile/rx_18/data_out_reg[15]  ( .D(n3504), .CK(CLK), .RN(n7777), 
        .Q(\regfile/reg_out[18][15] ), .QN(n5240) );
  DFFR_X1 \Scc_coproc/EPS_REG/data_out_reg[15]  ( .D(n3494), .CK(CLK), .RN(
        n7754), .QN(n5738) );
  DFFS_X1 \Scc_coproc/STATUS_REG/data_out_reg[15]  ( .D(n3493), .CK(CLK), .SN(
        n7823), .Q(kernel_mode), .QN(n5737) );
  DFFR_X1 \Mpath/regM/data_out_reg[16]  ( .D(n3485), .CK(CLK), .RN(n7793), 
        .QN(n5599) );
  DFFR_X1 \regfile/rx_5/data_out_reg[16]  ( .D(n3480), .CK(CLK), .RN(n7793), 
        .Q(\regfile/reg_out[5][16] ), .QN(n4663) );
  DFFR_X1 \regfile/rx_4/data_out_reg[16]  ( .D(n3479), .CK(CLK), .RN(n7793), 
        .Q(\regfile/reg_out[4][16] ), .QN(n4695) );
  DFFR_X1 \regfile/rx_29/data_out_reg[16]  ( .D(n3474), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[29][16] ), .QN(n4855) );
  DFFR_X1 \regfile/rx_28/data_out_reg[16]  ( .D(n3473), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[28][16] ), .QN(n4887) );
  DFFR_X1 \regfile/rx_25/data_out_reg[16]  ( .D(n3470), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[25][16] ), .QN(n4983) );
  DFFR_X1 \regfile/rx_24/data_out_reg[16]  ( .D(n3469), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[24][16] ), .QN(n5015) );
  DFFR_X1 \regfile/rx_21/data_out_reg[16]  ( .D(n3466), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[21][16] ), .QN(n5111) );
  DFFR_X1 \regfile/rx_20/data_out_reg[16]  ( .D(n3465), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[20][16] ), .QN(n5143) );
  DFFR_X1 \regfile/rx_19/data_out_reg[16]  ( .D(n3463), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[19][16] ), .QN(n5207) );
  DFFR_X1 \regfile/rx_18/data_out_reg[16]  ( .D(n3462), .CK(CLK), .RN(n7791), 
        .Q(\regfile/reg_out[18][16] ), .QN(n5239) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[16]  ( .D(n3447), .CK(CLK), .RN(
        n7785), .QN(n6316) );
  DFFR_X1 \Mpath/regM/data_out_reg[17]  ( .D(n3446), .CK(CLK), .RN(n7752), 
        .QN(n5596) );
  DFFR_X1 \regfile/rx_5/data_out_reg[17]  ( .D(n3441), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[5][17] ), .QN(n4662) );
  DFFR_X1 \regfile/rx_4/data_out_reg[17]  ( .D(n3440), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[4][17] ), .QN(n4694) );
  DFFR_X1 \regfile/rx_29/data_out_reg[17]  ( .D(n3435), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[29][17] ), .QN(n4854) );
  DFFR_X1 \regfile/rx_28/data_out_reg[17]  ( .D(n3434), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[28][17] ), .QN(n4886) );
  DFFR_X1 \regfile/rx_25/data_out_reg[17]  ( .D(n3431), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[25][17] ), .QN(n4982) );
  DFFR_X1 \regfile/rx_24/data_out_reg[17]  ( .D(n3430), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[24][17] ), .QN(n5014) );
  DFFR_X1 \regfile/rx_21/data_out_reg[17]  ( .D(n3427), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[21][17] ), .QN(n5110) );
  DFFR_X1 \regfile/rx_20/data_out_reg[17]  ( .D(n3426), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[20][17] ), .QN(n5142) );
  DFFR_X1 \regfile/rx_19/data_out_reg[17]  ( .D(n3424), .CK(CLK), .RN(n7761), 
        .Q(\regfile/reg_out[19][17] ), .QN(n5206) );
  DFFR_X1 \regfile/rx_18/data_out_reg[17]  ( .D(n3423), .CK(CLK), .RN(n7761), 
        .Q(\regfile/reg_out[18][17] ), .QN(n5238) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[17]  ( .D(n3408), .CK(CLK), .RN(
        n7785), .QN(n6304) );
  DFFR_X1 \Mpath/regM/data_out_reg[18]  ( .D(n3407), .CK(CLK), .RN(n7821), 
        .QN(n5593) );
  DFFR_X1 \regfile/rx_5/data_out_reg[18]  ( .D(n3402), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[5][18] ), .QN(n4661) );
  DFFR_X1 \regfile/rx_4/data_out_reg[18]  ( .D(n3401), .CK(CLK), .RN(n7821), 
        .Q(\regfile/reg_out[4][18] ), .QN(n4693) );
  DFFR_X1 \regfile/rx_29/data_out_reg[18]  ( .D(n3396), .CK(CLK), .RN(n7822), 
        .Q(\regfile/reg_out[29][18] ), .QN(n4853) );
  DFFR_X1 \regfile/rx_28/data_out_reg[18]  ( .D(n3395), .CK(CLK), .RN(n7822), 
        .Q(\regfile/reg_out[28][18] ), .QN(n4885) );
  DFFR_X1 \regfile/rx_25/data_out_reg[18]  ( .D(n3392), .CK(CLK), .RN(n7821), 
        .Q(\regfile/reg_out[25][18] ), .QN(n4981) );
  DFFR_X1 \regfile/rx_24/data_out_reg[18]  ( .D(n3391), .CK(CLK), .RN(n7821), 
        .Q(\regfile/reg_out[24][18] ), .QN(n5013) );
  DFFR_X1 \regfile/rx_21/data_out_reg[18]  ( .D(n3388), .CK(CLK), .RN(n7822), 
        .Q(\regfile/reg_out[21][18] ), .QN(n5109) );
  DFFR_X1 \regfile/rx_20/data_out_reg[18]  ( .D(n3387), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[20][18] ), .QN(n5141) );
  DFFR_X1 \regfile/rx_19/data_out_reg[18]  ( .D(n3385), .CK(CLK), .RN(n7815), 
        .Q(\regfile/reg_out[19][18] ), .QN(n5205) );
  DFFR_X1 \regfile/rx_18/data_out_reg[18]  ( .D(n3384), .CK(CLK), .RN(n7815), 
        .Q(\regfile/reg_out[18][18] ), .QN(n5237) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[18]  ( .D(n3369), .CK(CLK), .RN(
        n7788), .QN(n6290) );
  DFFR_X1 \Mpath/regM/data_out_reg[19]  ( .D(n3368), .CK(CLK), .RN(n7734), 
        .QN(n5590) );
  DFFR_X1 \regfile/rx_5/data_out_reg[19]  ( .D(n3363), .CK(CLK), .RN(n7734), 
        .Q(\regfile/reg_out[5][19] ), .QN(n4660) );
  DFFR_X1 \regfile/rx_4/data_out_reg[19]  ( .D(n3362), .CK(CLK), .RN(n7734), 
        .Q(\regfile/reg_out[4][19] ), .QN(n4692) );
  DFFR_X1 \regfile/rx_29/data_out_reg[19]  ( .D(n3357), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[29][19] ), .QN(n4852) );
  DFFR_X1 \regfile/rx_28/data_out_reg[19]  ( .D(n3356), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[28][19] ), .QN(n4884) );
  DFFR_X1 \regfile/rx_25/data_out_reg[19]  ( .D(n3353), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[25][19] ), .QN(n4980) );
  DFFR_X1 \regfile/rx_24/data_out_reg[19]  ( .D(n3352), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[24][19] ), .QN(n5012) );
  DFFR_X1 \regfile/rx_21/data_out_reg[19]  ( .D(n3349), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[21][19] ), .QN(n5108) );
  DFFR_X1 \regfile/rx_20/data_out_reg[19]  ( .D(n3348), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[20][19] ), .QN(n5140) );
  DFFR_X1 \regfile/rx_19/data_out_reg[19]  ( .D(n3346), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[19][19] ), .QN(n5204) );
  DFFR_X1 \regfile/rx_18/data_out_reg[19]  ( .D(n3345), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[18][19] ), .QN(n5236) );
  DFFR_X1 \Mpath/regB/data_out_reg[19]  ( .D(n3335), .CK(CLK), .RN(n7731), .Q(
        \Mpath/out_regB[19] ), .QN(\Mpath/the_alu/N46 ) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[19]  ( .D(n3330), .CK(CLK), .RN(
        n7788), .QN(n6275) );
  DFFR_X1 \Mpath/regM/data_out_reg[20]  ( .D(n3329), .CK(CLK), .RN(n7770), 
        .QN(n5584) );
  DFFR_X1 \regfile/rx_5/data_out_reg[20]  ( .D(n3324), .CK(CLK), .RN(n7769), 
        .Q(\regfile/reg_out[5][20] ), .QN(n4658) );
  DFFR_X1 \regfile/rx_4/data_out_reg[20]  ( .D(n3323), .CK(CLK), .RN(n7769), 
        .Q(\regfile/reg_out[4][20] ), .QN(n4690) );
  DFFR_X1 \regfile/rx_29/data_out_reg[20]  ( .D(n3318), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[29][20] ), .QN(n4850) );
  DFFR_X1 \regfile/rx_28/data_out_reg[20]  ( .D(n3317), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[28][20] ), .QN(n4882) );
  DFFR_X1 \regfile/rx_25/data_out_reg[20]  ( .D(n3314), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[25][20] ), .QN(n4978) );
  DFFR_X1 \regfile/rx_24/data_out_reg[20]  ( .D(n3313), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[24][20] ), .QN(n5010) );
  DFFR_X1 \regfile/rx_21/data_out_reg[20]  ( .D(n3310), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[21][20] ), .QN(n5106) );
  DFFR_X1 \regfile/rx_20/data_out_reg[20]  ( .D(n3309), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[20][20] ), .QN(n5138) );
  DFFR_X1 \regfile/rx_19/data_out_reg[20]  ( .D(n3307), .CK(CLK), .RN(n7794), 
        .Q(\regfile/reg_out[19][20] ), .QN(n5202) );
  DFFR_X1 \regfile/rx_18/data_out_reg[20]  ( .D(n3306), .CK(CLK), .RN(n7794), 
        .Q(\regfile/reg_out[18][20] ), .QN(n5234) );
  DFFR_X1 \Mpath/regB/data_out_reg[20]  ( .D(n3296), .CK(CLK), .RN(n7790), .Q(
        \Mpath/out_regB[20] ), .QN(\Mpath/the_alu/N44 ) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[20]  ( .D(n3291), .CK(CLK), .RN(
        n7786), .QN(n6262) );
  DFFR_X1 \Mpath/regM/data_out_reg[21]  ( .D(n3290), .CK(CLK), .RN(n7751), 
        .QN(n5581) );
  DFFR_X1 \regfile/rx_5/data_out_reg[21]  ( .D(n3285), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[5][21] ), .QN(n4657) );
  DFFR_X1 \regfile/rx_4/data_out_reg[21]  ( .D(n3284), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[4][21] ), .QN(n4689) );
  DFFR_X1 \regfile/rx_29/data_out_reg[21]  ( .D(n3279), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[29][21] ), .QN(n4849) );
  DFFR_X1 \regfile/rx_28/data_out_reg[21]  ( .D(n3278), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[28][21] ), .QN(n4881) );
  DFFR_X1 \regfile/rx_25/data_out_reg[21]  ( .D(n3275), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[25][21] ), .QN(n4977) );
  DFFR_X1 \regfile/rx_24/data_out_reg[21]  ( .D(n3274), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[24][21] ), .QN(n5009) );
  DFFR_X1 \regfile/rx_21/data_out_reg[21]  ( .D(n3271), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[21][21] ), .QN(n5105) );
  DFFR_X1 \regfile/rx_20/data_out_reg[21]  ( .D(n3270), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[20][21] ), .QN(n5137) );
  DFFR_X1 \regfile/rx_19/data_out_reg[21]  ( .D(n3268), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[19][21] ), .QN(n5201) );
  DFFR_X1 \regfile/rx_18/data_out_reg[21]  ( .D(n3267), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[18][21] ), .QN(n5233) );
  DFFR_X1 \Mpath/regB/data_out_reg[21]  ( .D(n3257), .CK(CLK), .RN(n7751), .Q(
        \Mpath/out_regB[21] ), .QN(\Mpath/the_alu/N42 ) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[21]  ( .D(n3252), .CK(CLK), .RN(
        n7786), .QN(n6246) );
  DFFR_X1 \Mpath/regM/data_out_reg[22]  ( .D(n3251), .CK(CLK), .RN(n7814), 
        .QN(n5578) );
  DFFR_X1 \regfile/rx_5/data_out_reg[22]  ( .D(n3246), .CK(CLK), .RN(n7814), 
        .Q(\regfile/reg_out[5][22] ), .QN(n4656) );
  DFFR_X1 \regfile/rx_4/data_out_reg[22]  ( .D(n3245), .CK(CLK), .RN(n7814), 
        .Q(\regfile/reg_out[4][22] ), .QN(n4688) );
  DFFR_X1 \regfile/rx_29/data_out_reg[22]  ( .D(n3240), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[29][22] ), .QN(n4848) );
  DFFR_X1 \regfile/rx_28/data_out_reg[22]  ( .D(n3239), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[28][22] ), .QN(n4880) );
  DFFR_X1 \regfile/rx_25/data_out_reg[22]  ( .D(n3236), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[25][22] ), .QN(n4976) );
  DFFR_X1 \regfile/rx_24/data_out_reg[22]  ( .D(n3235), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[24][22] ), .QN(n5008) );
  DFFR_X1 \regfile/rx_21/data_out_reg[22]  ( .D(n3232), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[21][22] ), .QN(n5104) );
  DFFR_X1 \regfile/rx_20/data_out_reg[22]  ( .D(n3231), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[20][22] ), .QN(n5136) );
  DFFR_X1 \regfile/rx_19/data_out_reg[22]  ( .D(n3229), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[19][22] ), .QN(n5200) );
  DFFR_X1 \regfile/rx_18/data_out_reg[22]  ( .D(n3228), .CK(CLK), .RN(n7812), 
        .Q(\regfile/reg_out[18][22] ), .QN(n5232) );
  DFFR_X1 \Mpath/regB/data_out_reg[22]  ( .D(n3218), .CK(CLK), .RN(n7789), .Q(
        \Mpath/out_regB[22] ), .QN(\Mpath/the_alu/N40 ) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[22]  ( .D(n3213), .CK(CLK), .RN(
        n7716), .QN(n6234) );
  DFFR_X1 \Mpath/regM/data_out_reg[24]  ( .D(n3212), .CK(CLK), .RN(n7731), 
        .QN(n5572) );
  DFFR_X1 \regfile/rx_5/data_out_reg[24]  ( .D(n3207), .CK(CLK), .RN(n7731), 
        .Q(\regfile/reg_out[5][24] ), .QN(n4654) );
  DFFR_X1 \regfile/rx_4/data_out_reg[24]  ( .D(n3206), .CK(CLK), .RN(n7731), 
        .Q(\regfile/reg_out[4][24] ), .QN(n4686) );
  DFFR_X1 \regfile/rx_29/data_out_reg[24]  ( .D(n3201), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[29][24] ), .QN(n4846) );
  DFFR_X1 \regfile/rx_28/data_out_reg[24]  ( .D(n3200), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[28][24] ), .QN(n4878) );
  DFFR_X1 \regfile/rx_25/data_out_reg[24]  ( .D(n3197), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[25][24] ), .QN(n4974) );
  DFFR_X1 \regfile/rx_24/data_out_reg[24]  ( .D(n3196), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[24][24] ), .QN(n5006) );
  DFFR_X1 \regfile/rx_21/data_out_reg[24]  ( .D(n3193), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[21][24] ), .QN(n5102) );
  DFFR_X1 \regfile/rx_20/data_out_reg[24]  ( .D(n3192), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[20][24] ), .QN(n5134) );
  DFFR_X1 \regfile/rx_19/data_out_reg[24]  ( .D(n3190), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[19][24] ), .QN(n5198) );
  DFFR_X1 \regfile/rx_18/data_out_reg[24]  ( .D(n3189), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[18][24] ), .QN(n5230) );
  DFFR_X1 \Mpath/regB/data_out_reg[24]  ( .D(n3179), .CK(CLK), .RN(n7809), .Q(
        \Mpath/out_regB[24] ), .QN(\Mpath/the_alu/N36 ) );
  DFFR_X1 \Mpath/regM/data_out_reg[25]  ( .D(n3178), .CK(CLK), .RN(n7751), 
        .QN(n5569) );
  DFFR_X1 \regfile/rx_5/data_out_reg[25]  ( .D(n3173), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[5][25] ), .QN(n4653) );
  DFFR_X1 \regfile/rx_4/data_out_reg[25]  ( .D(n3172), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[4][25] ), .QN(n4685) );
  DFFR_X1 \regfile/rx_29/data_out_reg[25]  ( .D(n3167), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[29][25] ), .QN(n4845) );
  DFFR_X1 \regfile/rx_28/data_out_reg[25]  ( .D(n3166), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[28][25] ), .QN(n4877) );
  DFFR_X1 \regfile/rx_25/data_out_reg[25]  ( .D(n3163), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[25][25] ), .QN(n4973) );
  DFFR_X1 \regfile/rx_24/data_out_reg[25]  ( .D(n3162), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[24][25] ), .QN(n5005) );
  DFFR_X1 \regfile/rx_21/data_out_reg[25]  ( .D(n3159), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[21][25] ), .QN(n5101) );
  DFFR_X1 \regfile/rx_20/data_out_reg[25]  ( .D(n3158), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[20][25] ), .QN(n5133) );
  DFFR_X1 \regfile/rx_19/data_out_reg[25]  ( .D(n3156), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[19][25] ), .QN(n5197) );
  DFFR_X1 \regfile/rx_18/data_out_reg[25]  ( .D(n3155), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[18][25] ), .QN(n5229) );
  DFFR_X1 \Mpath/regB/data_out_reg[25]  ( .D(n3145), .CK(CLK), .RN(n7751), .Q(
        \Mpath/out_regB[25] ), .QN(\Mpath/the_alu/N34 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[26]  ( .D(n3144), .CK(CLK), .RN(n7789), .Q(
        \Mpath/out_regB[26] ), .QN(\Mpath/the_alu/N32 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[27]  ( .D(n3143), .CK(CLK), .RN(n7806), .Q(
        \Mpath/out_regB[27] ), .QN(\Mpath/the_alu/N30 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[28]  ( .D(n3142), .CK(CLK), .RN(n7789), .Q(
        \Mpath/out_regB[28] ), .QN(\Mpath/the_alu/N28 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[29]  ( .D(n3141), .CK(CLK), .RN(n7787), .Q(
        \Mpath/out_regB[29] ), .QN(\Mpath/the_alu/N26 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[30]  ( .D(n3140), .CK(CLK), .RN(n7751), .Q(
        \Mpath/out_regB[30] ), .QN(\Mpath/the_alu/N24 ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[0]  ( .D(n3139), .CK(CLK), 
        .RN(n7745), .Q(D_DATA_OUTBUS[0]), .QN(n6441) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[1]  ( .D(n3138), .CK(CLK), 
        .RN(n7720), .Q(D_DATA_OUTBUS[1]), .QN(n6438) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[2]  ( .D(n3137), .CK(CLK), 
        .RN(n7748), .Q(D_DATA_OUTBUS[2]), .QN(n6461) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[3]  ( .D(n3136), .CK(CLK), 
        .RN(n7800), .Q(D_DATA_OUTBUS[3]), .QN(n6458) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[4]  ( .D(n3135), .CK(CLK), 
        .RN(n7717), .Q(D_DATA_OUTBUS[4]), .QN(n6455) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[5]  ( .D(n3134), .CK(CLK), 
        .RN(n7797), .Q(D_DATA_OUTBUS[5]), .QN(n6452) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[6]  ( .D(n3133), .CK(CLK), 
        .RN(n7738), .Q(D_DATA_OUTBUS[6]), .QN(n6449) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[7]  ( .D(n3132), .CK(CLK), 
        .RN(n7817), .Q(D_DATA_OUTBUS[7]), .QN(n6445) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[8]  ( .D(n3131), .CK(CLK), 
        .RN(n7726), .Q(\Mpath/the_memhandle/smdr_out[8] ), .QN(n6442) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[9]  ( .D(n3130), .CK(CLK), 
        .RN(n7782), .Q(\Mpath/the_memhandle/smdr_out[9] ), .QN(n6440) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[10]  ( .D(n3129), .CK(CLK), 
        .RN(n7779), .Q(\Mpath/the_memhandle/smdr_out[10] ), .QN(n6460) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[11]  ( .D(n3128), .CK(CLK), 
        .RN(n7735), .Q(\Mpath/the_memhandle/smdr_out[11] ), .QN(n6457) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[12]  ( .D(n3127), .CK(CLK), 
        .RN(n7773), .Q(\Mpath/the_memhandle/smdr_out[12] ), .QN(n6454) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[13]  ( .D(n3126), .CK(CLK), 
        .RN(n7723), .Q(\Mpath/the_memhandle/smdr_out[13] ), .QN(n6451) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[14]  ( .D(n3125), .CK(CLK), 
        .RN(n7770), .Q(\Mpath/the_memhandle/smdr_out[14] ), .QN(n6448) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[15]  ( .D(n3124), .CK(CLK), 
        .RN(n7776), .Q(\Mpath/the_memhandle/smdr_out[15] ), .QN(n6444) );
  OAI21_X1 U3 ( .B1(n6482), .B2(n7109), .A(n46), .ZN(serve_proc_addr[5]) );
  OAI22_X1 U4 ( .A1(n6484), .A2(n7109), .B1(n5740), .B2(n47), .ZN(
        serve_proc_addr[4]) );
  OAI22_X1 U5 ( .A1(n6487), .A2(n7109), .B1(n5740), .B2(n48), .ZN(
        serve_proc_addr[3]) );
  OAI22_X1 U6 ( .A1(n6489), .A2(n7109), .B1(n5740), .B2(n49), .ZN(
        serve_proc_addr[2]) );
  OAI221_X1 U7 ( .B1(n50), .B2(n51), .C1(n52), .C2(n53), .A(n54), .ZN(n3108)
         );
  AOI22_X1 U8 ( .A1(n55), .A2(n56), .B1(\Mpath/the_memhandle/smdr_out[31] ), 
        .B2(n57), .ZN(n54) );
  OAI221_X1 U9 ( .B1(n58), .B2(n51), .C1(n59), .C2(n53), .A(n60), .ZN(n3109)
         );
  AOI22_X1 U10 ( .A1(n55), .A2(n61), .B1(\Mpath/the_memhandle/smdr_out[30] ), 
        .B2(n57), .ZN(n60) );
  OAI221_X1 U11 ( .B1(n62), .B2(n51), .C1(n63), .C2(n53), .A(n64), .ZN(n3110)
         );
  AOI22_X1 U12 ( .A1(n55), .A2(n65), .B1(\Mpath/the_memhandle/smdr_out[29] ), 
        .B2(n57), .ZN(n64) );
  OAI221_X1 U13 ( .B1(n66), .B2(n51), .C1(n67), .C2(n53), .A(n68), .ZN(n3111)
         );
  AOI22_X1 U14 ( .A1(n55), .A2(n69), .B1(\Mpath/the_memhandle/smdr_out[28] ), 
        .B2(n57), .ZN(n68) );
  OAI221_X1 U15 ( .B1(n70), .B2(n51), .C1(n71), .C2(n53), .A(n72), .ZN(n3112)
         );
  AOI22_X1 U36 ( .A1(n55), .A2(n73), .B1(\Mpath/the_memhandle/smdr_out[27] ), 
        .B2(n57), .ZN(n72) );
  OAI221_X1 U37 ( .B1(n74), .B2(n51), .C1(n75), .C2(n53), .A(n76), .ZN(n3113)
         );
  AOI22_X1 U38 ( .A1(n55), .A2(n77), .B1(\Mpath/the_memhandle/smdr_out[26] ), 
        .B2(n57), .ZN(n76) );
  OAI221_X1 U39 ( .B1(n78), .B2(n51), .C1(n79), .C2(n53), .A(n80), .ZN(n3114)
         );
  AOI22_X1 U40 ( .A1(n55), .A2(n81), .B1(\Mpath/the_memhandle/smdr_out[25] ), 
        .B2(n57), .ZN(n80) );
  OAI221_X1 U41 ( .B1(n82), .B2(n51), .C1(n83), .C2(n53), .A(n84), .ZN(n3115)
         );
  AOI22_X1 U42 ( .A1(n55), .A2(n85), .B1(\Mpath/the_memhandle/smdr_out[24] ), 
        .B2(n57), .ZN(n84) );
  OAI221_X1 U43 ( .B1(n86), .B2(n51), .C1(n87), .C2(n53), .A(n88), .ZN(n3116)
         );
  AOI22_X1 U44 ( .A1(n55), .A2(n89), .B1(\Mpath/the_memhandle/smdr_out[23] ), 
        .B2(n57), .ZN(n88) );
  OAI221_X1 U45 ( .B1(n90), .B2(n51), .C1(n91), .C2(n53), .A(n92), .ZN(n3117)
         );
  AOI22_X1 U46 ( .A1(n55), .A2(n93), .B1(\Mpath/the_memhandle/smdr_out[22] ), 
        .B2(n57), .ZN(n92) );
  OAI221_X1 U47 ( .B1(n94), .B2(n51), .C1(n95), .C2(n53), .A(n96), .ZN(n3118)
         );
  AOI22_X1 U48 ( .A1(n55), .A2(n97), .B1(\Mpath/the_memhandle/smdr_out[21] ), 
        .B2(n57), .ZN(n96) );
  OAI221_X1 U49 ( .B1(n98), .B2(n51), .C1(n99), .C2(n53), .A(n100), .ZN(n3119)
         );
  AOI22_X1 U50 ( .A1(n55), .A2(n101), .B1(\Mpath/the_memhandle/smdr_out[20] ), 
        .B2(n57), .ZN(n100) );
  OAI221_X1 U51 ( .B1(n102), .B2(n51), .C1(n103), .C2(n53), .A(n104), .ZN(
        n3120) );
  AOI22_X1 U52 ( .A1(n55), .A2(n105), .B1(\Mpath/the_memhandle/smdr_out[19] ), 
        .B2(n57), .ZN(n104) );
  OAI221_X1 U53 ( .B1(n106), .B2(n51), .C1(n107), .C2(n53), .A(n108), .ZN(
        n3121) );
  AOI22_X1 U54 ( .A1(n55), .A2(n109), .B1(\Mpath/the_memhandle/smdr_out[18] ), 
        .B2(n57), .ZN(n108) );
  OAI221_X1 U55 ( .B1(n110), .B2(n51), .C1(n111), .C2(n53), .A(n112), .ZN(
        n3122) );
  AOI22_X1 U56 ( .A1(n55), .A2(n113), .B1(\Mpath/the_memhandle/smdr_out[17] ), 
        .B2(n57), .ZN(n112) );
  OAI221_X1 U57 ( .B1(n114), .B2(n51), .C1(n115), .C2(n53), .A(n116), .ZN(
        n3123) );
  AOI22_X1 U58 ( .A1(n55), .A2(n117), .B1(\Mpath/the_memhandle/smdr_out[16] ), 
        .B2(n57), .ZN(n116) );
  OAI221_X1 U59 ( .B1(n118), .B2(n51), .C1(n119), .C2(n53), .A(n120), .ZN(
        n3124) );
  AOI22_X1 U60 ( .A1(n55), .A2(n121), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[15] ), .ZN(n120) );
  OAI221_X1 U61 ( .B1(n122), .B2(n51), .C1(n123), .C2(n53), .A(n124), .ZN(
        n3125) );
  AOI22_X1 U62 ( .A1(n55), .A2(n125), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[14] ), .ZN(n124) );
  OAI221_X1 U63 ( .B1(n126), .B2(n51), .C1(n127), .C2(n53), .A(n128), .ZN(
        n3126) );
  AOI22_X1 U64 ( .A1(n55), .A2(n129), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[13] ), .ZN(n128) );
  OAI221_X1 U65 ( .B1(n130), .B2(n51), .C1(n131), .C2(n53), .A(n132), .ZN(
        n3127) );
  AOI22_X1 U66 ( .A1(n55), .A2(n133), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[12] ), .ZN(n132) );
  OAI221_X1 U67 ( .B1(n134), .B2(n51), .C1(n135), .C2(n53), .A(n136), .ZN(
        n3128) );
  AOI22_X1 U68 ( .A1(n55), .A2(n137), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[11] ), .ZN(n136) );
  OAI221_X1 U69 ( .B1(n138), .B2(n51), .C1(n139), .C2(n53), .A(n140), .ZN(
        n3129) );
  AOI22_X1 U70 ( .A1(n55), .A2(n141), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[10] ), .ZN(n140) );
  OAI221_X1 U71 ( .B1(n142), .B2(n51), .C1(n143), .C2(n53), .A(n144), .ZN(
        n3130) );
  AOI22_X1 U72 ( .A1(n55), .A2(n145), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[9] ), .ZN(n144) );
  OAI221_X1 U73 ( .B1(n146), .B2(n51), .C1(n147), .C2(n53), .A(n148), .ZN(
        n3131) );
  AOI22_X1 U74 ( .A1(n55), .A2(n149), .B1(n57), .B2(
        \Mpath/the_memhandle/smdr_out[8] ), .ZN(n148) );
  OAI221_X1 U75 ( .B1(n150), .B2(n51), .C1(n151), .C2(n53), .A(n152), .ZN(
        n3132) );
  AOI22_X1 U76 ( .A1(n55), .A2(n153), .B1(n57), .B2(D_DATA_OUTBUS[7]), .ZN(
        n152) );
  OAI221_X1 U77 ( .B1(n154), .B2(n51), .C1(n155), .C2(n53), .A(n156), .ZN(
        n3133) );
  AOI22_X1 U78 ( .A1(n55), .A2(n157), .B1(n57), .B2(D_DATA_OUTBUS[6]), .ZN(
        n156) );
  OAI221_X1 U79 ( .B1(n158), .B2(n51), .C1(n159), .C2(n53), .A(n160), .ZN(
        n3134) );
  AOI22_X1 U80 ( .A1(n55), .A2(n161), .B1(n57), .B2(D_DATA_OUTBUS[5]), .ZN(
        n160) );
  OAI221_X1 U81 ( .B1(n162), .B2(n51), .C1(n163), .C2(n53), .A(n164), .ZN(
        n3135) );
  AOI22_X1 U82 ( .A1(n55), .A2(n165), .B1(n57), .B2(D_DATA_OUTBUS[4]), .ZN(
        n164) );
  OAI221_X1 U83 ( .B1(n166), .B2(n51), .C1(n167), .C2(n53), .A(n168), .ZN(
        n3136) );
  AOI22_X1 U84 ( .A1(n55), .A2(n169), .B1(n57), .B2(D_DATA_OUTBUS[3]), .ZN(
        n168) );
  OAI221_X1 U85 ( .B1(n170), .B2(n51), .C1(n171), .C2(n53), .A(n172), .ZN(
        n3137) );
  AOI22_X1 U86 ( .A1(n55), .A2(n173), .B1(n57), .B2(D_DATA_OUTBUS[2]), .ZN(
        n172) );
  OAI221_X1 U87 ( .B1(n174), .B2(n51), .C1(n175), .C2(n53), .A(n176), .ZN(
        n3138) );
  AOI22_X1 U88 ( .A1(n55), .A2(n177), .B1(n57), .B2(D_DATA_OUTBUS[1]), .ZN(
        n176) );
  OAI221_X1 U89 ( .B1(n178), .B2(n51), .C1(n179), .C2(n53), .A(n180), .ZN(
        n3139) );
  AOI22_X1 U90 ( .A1(n55), .A2(n181), .B1(n57), .B2(D_DATA_OUTBUS[0]), .ZN(
        n180) );
  INV_X1 U94 ( .A(n57), .ZN(n183) );
  OAI211_X1 U96 ( .C1(\Mpath/the_alu/N24 ), .C2(net55862), .A(n188), .B(n189), 
        .ZN(n3140) );
  AOI221_X1 U97 ( .B1(n190), .B2(n191), .C1(n192), .C2(n193), .A(n194), .ZN(
        n189) );
  AOI22_X1 U98 ( .A1(n195), .A2(n196), .B1(n197), .B2(n61), .ZN(n188) );
  OAI211_X1 U99 ( .C1(\Mpath/the_alu/N26 ), .C2(net55862), .A(n198), .B(n199), 
        .ZN(n3141) );
  AOI221_X1 U100 ( .B1(n190), .B2(n200), .C1(n192), .C2(n201), .A(n194), .ZN(
        n199) );
  AOI22_X1 U101 ( .A1(n195), .A2(n202), .B1(n197), .B2(n65), .ZN(n198) );
  OAI211_X1 U102 ( .C1(\Mpath/the_alu/N28 ), .C2(net55862), .A(n203), .B(n204), 
        .ZN(n3142) );
  AOI221_X1 U103 ( .B1(n190), .B2(n205), .C1(n192), .C2(n206), .A(n194), .ZN(
        n204) );
  AOI22_X1 U104 ( .A1(n195), .A2(n207), .B1(n197), .B2(n69), .ZN(n203) );
  OAI211_X1 U105 ( .C1(\Mpath/the_alu/N30 ), .C2(net55862), .A(n208), .B(n209), 
        .ZN(n3143) );
  AOI221_X1 U106 ( .B1(n190), .B2(n210), .C1(n192), .C2(n211), .A(n194), .ZN(
        n209) );
  AOI21_X1 U107 ( .B1(n212), .B2(n213), .A(n214), .ZN(n194) );
  NAND2_X1 U108 ( .A1(n5854), .A2(n215), .ZN(n212) );
  AOI22_X1 U109 ( .A1(n195), .A2(n216), .B1(n197), .B2(n73), .ZN(n208) );
  NAND3_X1 U110 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n3144) );
  AOI222_X1 U111 ( .A1(net55898), .A2(n221), .B1(n195), .B2(n222), .C1(n197), 
        .C2(n77), .ZN(n219) );
  AOI21_X1 U112 ( .B1(n5891), .B2(n223), .A(n224), .ZN(n218) );
  AOI22_X1 U113 ( .A1(n192), .A2(n225), .B1(n5890), .B2(n190), .ZN(n217) );
  NAND3_X1 U114 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n3145) );
  AOI222_X1 U115 ( .A1(net55898), .A2(n229), .B1(n195), .B2(n230), .C1(n197), 
        .C2(n81), .ZN(n228) );
  AOI21_X1 U116 ( .B1(n5902), .B2(n223), .A(n224), .ZN(n227) );
  AOI22_X1 U117 ( .A1(n192), .A2(n231), .B1(n5901), .B2(n190), .ZN(n226) );
  OAI221_X1 U118 ( .B1(n79), .B2(n6554), .C1(\Mpath/the_alu/N33 ), .C2(
        net55856), .A(n233), .ZN(n3146) );
  AOI22_X1 U119 ( .A1(n6556), .A2(n231), .B1(n6560), .B2(n236), .ZN(n233) );
  OAI22_X1 U120 ( .A1(n237), .A2(n238), .B1(n79), .B2(n239), .ZN(n3147) );
  OAI22_X1 U121 ( .A1(n240), .A2(n241), .B1(n79), .B2(n7318), .ZN(n3148) );
  OAI22_X1 U122 ( .A1(n243), .A2(n244), .B1(n79), .B2(n7370), .ZN(n3149) );
  OAI22_X1 U124 ( .A1(n246), .A2(n247), .B1(n79), .B2(n248), .ZN(n3150) );
  OAI22_X1 U125 ( .A1(n249), .A2(n250), .B1(n79), .B2(n251), .ZN(n3151) );
  OAI22_X1 U126 ( .A1(n252), .A2(n253), .B1(n79), .B2(n7271), .ZN(n3152) );
  OAI22_X1 U127 ( .A1(n255), .A2(n256), .B1(n79), .B2(n257), .ZN(n3153) );
  OAI22_X1 U129 ( .A1(n258), .A2(n259), .B1(n79), .B2(n7117), .ZN(n3154) );
  OAI22_X1 U130 ( .A1(n7115), .A2(n5229), .B1(n79), .B2(n262), .ZN(n3155) );
  OAI22_X1 U131 ( .A1(n263), .A2(n5197), .B1(n79), .B2(n7158), .ZN(n3156) );
  OAI22_X1 U132 ( .A1(n6895), .A2(n266), .B1(n79), .B2(n6898), .ZN(n3157) );
  OAI22_X1 U133 ( .A1(n268), .A2(n5133), .B1(n79), .B2(n269), .ZN(n3158) );
  OAI22_X1 U134 ( .A1(n270), .A2(n5101), .B1(n79), .B2(n271), .ZN(n3159) );
  OAI22_X1 U135 ( .A1(n272), .A2(n273), .B1(n79), .B2(n274), .ZN(n3160) );
  OAI22_X1 U136 ( .A1(n275), .A2(n276), .B1(n79), .B2(n7363), .ZN(n3161) );
  OAI22_X1 U137 ( .A1(n278), .A2(n5005), .B1(n79), .B2(n7276), .ZN(n3162) );
  OAI22_X1 U138 ( .A1(n7122), .A2(n4973), .B1(n79), .B2(n281), .ZN(n3163) );
  OAI22_X1 U139 ( .A1(n282), .A2(n283), .B1(n79), .B2(n284), .ZN(n3164) );
  OAI22_X1 U140 ( .A1(n7119), .A2(n286), .B1(n79), .B2(n287), .ZN(n3165) );
  OAI22_X1 U141 ( .A1(n288), .A2(n4877), .B1(n79), .B2(n289), .ZN(n3166) );
  OAI22_X1 U142 ( .A1(n290), .A2(n4845), .B1(n79), .B2(n291), .ZN(n3167) );
  OAI22_X1 U143 ( .A1(n292), .A2(n293), .B1(n79), .B2(n294), .ZN(n3168) );
  OAI22_X1 U145 ( .A1(n295), .A2(n296), .B1(n79), .B2(n297), .ZN(n3169) );
  OAI22_X1 U147 ( .A1(n298), .A2(n299), .B1(n79), .B2(n300), .ZN(n3170) );
  OAI22_X1 U148 ( .A1(n6558), .A2(n302), .B1(n79), .B2(n7076), .ZN(n3171) );
  OAI22_X1 U150 ( .A1(n304), .A2(n4685), .B1(n79), .B2(n7113), .ZN(n3172) );
  OAI22_X1 U151 ( .A1(n7112), .A2(n4653), .B1(n79), .B2(n307), .ZN(n3173) );
  OAI22_X1 U152 ( .A1(n308), .A2(n309), .B1(n79), .B2(n310), .ZN(n3174) );
  OAI22_X1 U153 ( .A1(n7074), .A2(n312), .B1(n79), .B2(n313), .ZN(n3175) );
  OAI22_X1 U154 ( .A1(n314), .A2(n315), .B1(n79), .B2(n7210), .ZN(n3176) );
  OAI22_X1 U155 ( .A1(n317), .A2(n318), .B1(n79), .B2(n7209), .ZN(n3177) );
  OAI221_X1 U157 ( .B1(n5895), .B2(n320), .C1(n5745), .C2(n5569), .A(n321), 
        .ZN(n230) );
  OAI22_X1 U158 ( .A1(n5569), .A2(net55842), .B1(n78), .B2(net55906), .ZN(
        n3178) );
  INV_X1 U159 ( .A(n231), .ZN(n78) );
  OAI22_X1 U160 ( .A1(n5698), .A2(n322), .B1(n5699), .B2(n323), .ZN(n231) );
  NAND3_X1 U161 ( .A1(n324), .A2(n325), .A3(n326), .ZN(n3179) );
  AOI222_X1 U162 ( .A1(net55898), .A2(n327), .B1(n195), .B2(n328), .C1(n197), 
        .C2(n85), .ZN(n326) );
  AOI21_X1 U163 ( .B1(n5912), .B2(n223), .A(n224), .ZN(n325) );
  AND2_X1 U164 ( .A1(n329), .A2(n330), .ZN(n224) );
  AND2_X1 U165 ( .A1(n331), .A2(n329), .ZN(n223) );
  AOI22_X1 U166 ( .A1(n192), .A2(n332), .B1(n5911), .B2(n190), .ZN(n324) );
  AND2_X1 U167 ( .A1(n333), .A2(n329), .ZN(n190) );
  OAI221_X1 U168 ( .B1(n83), .B2(n6554), .C1(\Mpath/the_alu/N35 ), .C2(
        net55856), .A(n334), .ZN(n3180) );
  AOI22_X1 U169 ( .A1(n6556), .A2(n332), .B1(n6560), .B2(n335), .ZN(n334) );
  OAI22_X1 U170 ( .A1(n237), .A2(n336), .B1(n83), .B2(n239), .ZN(n3181) );
  OAI22_X1 U171 ( .A1(n240), .A2(n337), .B1(n83), .B2(n7318), .ZN(n3182) );
  OAI22_X1 U172 ( .A1(n243), .A2(n338), .B1(n83), .B2(n7370), .ZN(n3183) );
  OAI22_X1 U174 ( .A1(n246), .A2(n339), .B1(n83), .B2(n248), .ZN(n3184) );
  OAI22_X1 U175 ( .A1(n249), .A2(n340), .B1(n83), .B2(n251), .ZN(n3185) );
  OAI22_X1 U176 ( .A1(n252), .A2(n341), .B1(n83), .B2(n7271), .ZN(n3186) );
  OAI22_X1 U177 ( .A1(n255), .A2(n342), .B1(n83), .B2(n257), .ZN(n3187) );
  OAI22_X1 U179 ( .A1(n258), .A2(n343), .B1(n83), .B2(n7117), .ZN(n3188) );
  OAI22_X1 U180 ( .A1(n7115), .A2(n5230), .B1(n83), .B2(n262), .ZN(n3189) );
  OAI22_X1 U181 ( .A1(n263), .A2(n5198), .B1(n83), .B2(n7158), .ZN(n3190) );
  OAI22_X1 U182 ( .A1(n6897), .A2(n344), .B1(n83), .B2(n6898), .ZN(n3191) );
  OAI22_X1 U183 ( .A1(n268), .A2(n5134), .B1(n83), .B2(n269), .ZN(n3192) );
  OAI22_X1 U184 ( .A1(n270), .A2(n5102), .B1(n83), .B2(n271), .ZN(n3193) );
  OAI22_X1 U185 ( .A1(n272), .A2(n345), .B1(n83), .B2(n274), .ZN(n3194) );
  OAI22_X1 U186 ( .A1(n275), .A2(n346), .B1(n83), .B2(n7363), .ZN(n3195) );
  OAI22_X1 U187 ( .A1(n278), .A2(n5006), .B1(n83), .B2(n7276), .ZN(n3196) );
  OAI22_X1 U188 ( .A1(n7122), .A2(n4974), .B1(n83), .B2(n281), .ZN(n3197) );
  OAI22_X1 U189 ( .A1(n282), .A2(n347), .B1(n83), .B2(n284), .ZN(n3198) );
  OAI22_X1 U190 ( .A1(n7119), .A2(n348), .B1(n83), .B2(n287), .ZN(n3199) );
  OAI22_X1 U191 ( .A1(n288), .A2(n4878), .B1(n83), .B2(n289), .ZN(n3200) );
  OAI22_X1 U192 ( .A1(n290), .A2(n4846), .B1(n83), .B2(n291), .ZN(n3201) );
  OAI22_X1 U193 ( .A1(n292), .A2(n349), .B1(n83), .B2(n294), .ZN(n3202) );
  OAI22_X1 U195 ( .A1(n295), .A2(n350), .B1(n83), .B2(n297), .ZN(n3203) );
  OAI22_X1 U197 ( .A1(n298), .A2(n351), .B1(n83), .B2(n300), .ZN(n3204) );
  OAI22_X1 U198 ( .A1(n6559), .A2(n352), .B1(n83), .B2(n7076), .ZN(n3205) );
  OAI22_X1 U200 ( .A1(n304), .A2(n4686), .B1(n83), .B2(n7113), .ZN(n3206) );
  OAI22_X1 U201 ( .A1(n7112), .A2(n4654), .B1(n83), .B2(n307), .ZN(n3207) );
  OAI22_X1 U202 ( .A1(n308), .A2(n353), .B1(n83), .B2(n310), .ZN(n3208) );
  OAI22_X1 U203 ( .A1(n7074), .A2(n354), .B1(n83), .B2(n313), .ZN(n3209) );
  OAI22_X1 U204 ( .A1(n314), .A2(n355), .B1(n83), .B2(n7210), .ZN(n3210) );
  OAI22_X1 U205 ( .A1(n317), .A2(n356), .B1(n83), .B2(n7209), .ZN(n3211) );
  OAI221_X1 U207 ( .B1(n5905), .B2(n320), .C1(n5745), .C2(n5572), .A(n321), 
        .ZN(n328) );
  OAI22_X1 U208 ( .A1(n5572), .A2(net55842), .B1(n82), .B2(net55906), .ZN(
        n3212) );
  INV_X1 U209 ( .A(n332), .ZN(n82) );
  OAI22_X1 U210 ( .A1(n5706), .A2(n322), .B1(n5707), .B2(n323), .ZN(n332) );
  OAI221_X1 U211 ( .B1(n357), .B2(n358), .C1(n6234), .C2(n359), .A(n360), .ZN(
        n3213) );
  AOI22_X1 U212 ( .A1(\Mcontrol/bvgen/d_curr_pc[22] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [22]), .B2(n362), .ZN(n360) );
  OAI222_X1 U213 ( .A1(n363), .A2(n364), .B1(n365), .B2(n366), .C1(net55850), 
        .C2(n358), .ZN(n3214) );
  OAI22_X1 U215 ( .A1(net55888), .A2(n365), .B1(net55830), .B2(n363), .ZN(
        n3215) );
  INV_X1 U218 ( .A(n367), .ZN(n3216) );
  AOI22_X1 U219 ( .A1(n7189), .A2(\Mcontrol/f_currpc[22] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[22] ), .ZN(n367) );
  OAI221_X1 U222 ( .B1(n374), .B2(n214), .C1(\Mpath/the_alu/N40 ), .C2(
        net55858), .A(n375), .ZN(n3218) );
  AOI222_X1 U223 ( .A1(n197), .A2(n93), .B1(n192), .B2(n376), .C1(n195), .C2(
        n377), .ZN(n375) );
  OAI221_X1 U224 ( .B1(n91), .B2(n232), .C1(\Mpath/the_alu/N39 ), .C2(net55858), .A(n378), .ZN(n3219) );
  AOI22_X1 U225 ( .A1(n6556), .A2(n376), .B1(n6560), .B2(n379), .ZN(n378) );
  OAI22_X1 U226 ( .A1(n237), .A2(n380), .B1(n91), .B2(n239), .ZN(n3220) );
  OAI22_X1 U227 ( .A1(n240), .A2(n381), .B1(n91), .B2(n7318), .ZN(n3221) );
  OAI22_X1 U228 ( .A1(n243), .A2(n382), .B1(n91), .B2(n7370), .ZN(n3222) );
  OAI22_X1 U230 ( .A1(n246), .A2(n383), .B1(n91), .B2(n248), .ZN(n3223) );
  OAI22_X1 U231 ( .A1(n249), .A2(n384), .B1(n91), .B2(n251), .ZN(n3224) );
  OAI22_X1 U232 ( .A1(n252), .A2(n385), .B1(n91), .B2(n7271), .ZN(n3225) );
  OAI22_X1 U233 ( .A1(n255), .A2(n386), .B1(n91), .B2(n257), .ZN(n3226) );
  OAI22_X1 U235 ( .A1(n258), .A2(n387), .B1(n91), .B2(n7117), .ZN(n3227) );
  OAI22_X1 U236 ( .A1(n7115), .A2(n5232), .B1(n91), .B2(n262), .ZN(n3228) );
  OAI22_X1 U237 ( .A1(n263), .A2(n5200), .B1(n91), .B2(n7158), .ZN(n3229) );
  OAI22_X1 U238 ( .A1(n6896), .A2(n388), .B1(n91), .B2(n6898), .ZN(n3230) );
  OAI22_X1 U239 ( .A1(n268), .A2(n5136), .B1(n91), .B2(n269), .ZN(n3231) );
  OAI22_X1 U240 ( .A1(n270), .A2(n5104), .B1(n91), .B2(n271), .ZN(n3232) );
  OAI22_X1 U241 ( .A1(n272), .A2(n389), .B1(n91), .B2(n274), .ZN(n3233) );
  OAI22_X1 U242 ( .A1(n275), .A2(n390), .B1(n91), .B2(n7363), .ZN(n3234) );
  OAI22_X1 U243 ( .A1(n278), .A2(n5008), .B1(n91), .B2(n7276), .ZN(n3235) );
  OAI22_X1 U244 ( .A1(n7122), .A2(n4976), .B1(n91), .B2(n281), .ZN(n3236) );
  OAI22_X1 U245 ( .A1(n282), .A2(n391), .B1(n91), .B2(n284), .ZN(n3237) );
  OAI22_X1 U246 ( .A1(n7119), .A2(n392), .B1(n91), .B2(n287), .ZN(n3238) );
  OAI22_X1 U247 ( .A1(n288), .A2(n4880), .B1(n91), .B2(n289), .ZN(n3239) );
  OAI22_X1 U248 ( .A1(n290), .A2(n4848), .B1(n91), .B2(n291), .ZN(n3240) );
  OAI22_X1 U249 ( .A1(n292), .A2(n393), .B1(n91), .B2(n294), .ZN(n3241) );
  OAI22_X1 U251 ( .A1(n295), .A2(n394), .B1(n91), .B2(n297), .ZN(n3242) );
  OAI22_X1 U253 ( .A1(n298), .A2(n395), .B1(n91), .B2(n300), .ZN(n3243) );
  OAI22_X1 U254 ( .A1(n6558), .A2(n396), .B1(n91), .B2(n7076), .ZN(n3244) );
  OAI22_X1 U256 ( .A1(n304), .A2(n4688), .B1(n91), .B2(n7113), .ZN(n3245) );
  OAI22_X1 U257 ( .A1(n7112), .A2(n4656), .B1(n91), .B2(n307), .ZN(n3246) );
  OAI22_X1 U258 ( .A1(n308), .A2(n397), .B1(n91), .B2(n310), .ZN(n3247) );
  OAI22_X1 U259 ( .A1(n7074), .A2(n398), .B1(n91), .B2(n313), .ZN(n3248) );
  OAI22_X1 U260 ( .A1(n314), .A2(n399), .B1(n91), .B2(n7210), .ZN(n3249) );
  OAI22_X1 U261 ( .A1(n317), .A2(n400), .B1(n91), .B2(n7209), .ZN(n3250) );
  OAI221_X1 U263 ( .B1(n5803), .B2(n320), .C1(n5745), .C2(n5578), .A(n321), 
        .ZN(n377) );
  OAI22_X1 U264 ( .A1(n5578), .A2(net55842), .B1(n90), .B2(net55902), .ZN(
        n3251) );
  INV_X1 U265 ( .A(n376), .ZN(n90) );
  OAI222_X1 U266 ( .A1(n401), .A2(n323), .B1(n6235), .B2(n402), .C1(n403), 
        .C2(n322), .ZN(n376) );
  INV_X1 U267 ( .A(n6238), .ZN(n403) );
  INV_X1 U268 ( .A(n6237), .ZN(n401) );
  OAI221_X1 U269 ( .B1(n357), .B2(n404), .C1(n6246), .C2(n359), .A(n405), .ZN(
        n3252) );
  AOI22_X1 U270 ( .A1(\Mcontrol/bvgen/d_curr_pc[21] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [21]), .B2(n362), .ZN(n405) );
  OAI222_X1 U271 ( .A1(n364), .A2(n406), .B1(n366), .B2(n407), .C1(net55848), 
        .C2(n404), .ZN(n3253) );
  OAI22_X1 U273 ( .A1(net55888), .A2(n407), .B1(net55832), .B2(n406), .ZN(
        n3254) );
  INV_X1 U276 ( .A(n408), .ZN(n3255) );
  AOI22_X1 U277 ( .A1(n7189), .A2(\Mcontrol/f_currpc[21] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[21] ), .ZN(n408) );
  OAI221_X1 U280 ( .B1(n410), .B2(n214), .C1(\Mpath/the_alu/N42 ), .C2(
        net55858), .A(n411), .ZN(n3257) );
  AOI222_X1 U281 ( .A1(n197), .A2(n97), .B1(n192), .B2(n412), .C1(n195), .C2(
        n413), .ZN(n411) );
  OAI221_X1 U282 ( .B1(n95), .B2(n6554), .C1(\Mpath/the_alu/N41 ), .C2(
        net55858), .A(n414), .ZN(n3258) );
  AOI22_X1 U283 ( .A1(n6556), .A2(n412), .B1(n6560), .B2(n415), .ZN(n414) );
  OAI22_X1 U284 ( .A1(n237), .A2(n416), .B1(n95), .B2(n239), .ZN(n3259) );
  OAI22_X1 U285 ( .A1(n240), .A2(n417), .B1(n95), .B2(n7318), .ZN(n3260) );
  OAI22_X1 U286 ( .A1(n243), .A2(n418), .B1(n95), .B2(n7370), .ZN(n3261) );
  OAI22_X1 U288 ( .A1(n246), .A2(n419), .B1(n95), .B2(n248), .ZN(n3262) );
  OAI22_X1 U289 ( .A1(n249), .A2(n420), .B1(n95), .B2(n251), .ZN(n3263) );
  OAI22_X1 U290 ( .A1(n252), .A2(n421), .B1(n95), .B2(n7271), .ZN(n3264) );
  OAI22_X1 U291 ( .A1(n255), .A2(n422), .B1(n95), .B2(n257), .ZN(n3265) );
  OAI22_X1 U293 ( .A1(n258), .A2(n423), .B1(n95), .B2(n7117), .ZN(n3266) );
  OAI22_X1 U294 ( .A1(n7115), .A2(n5233), .B1(n95), .B2(n262), .ZN(n3267) );
  OAI22_X1 U295 ( .A1(n263), .A2(n5201), .B1(n95), .B2(n7158), .ZN(n3268) );
  OAI22_X1 U296 ( .A1(n6896), .A2(n424), .B1(n95), .B2(n6898), .ZN(n3269) );
  OAI22_X1 U297 ( .A1(n268), .A2(n5137), .B1(n95), .B2(n269), .ZN(n3270) );
  OAI22_X1 U298 ( .A1(n270), .A2(n5105), .B1(n95), .B2(n271), .ZN(n3271) );
  OAI22_X1 U299 ( .A1(n272), .A2(n425), .B1(n95), .B2(n274), .ZN(n3272) );
  OAI22_X1 U300 ( .A1(n275), .A2(n426), .B1(n95), .B2(n7363), .ZN(n3273) );
  OAI22_X1 U301 ( .A1(n278), .A2(n5009), .B1(n95), .B2(n7276), .ZN(n3274) );
  OAI22_X1 U302 ( .A1(n7122), .A2(n4977), .B1(n95), .B2(n281), .ZN(n3275) );
  OAI22_X1 U303 ( .A1(n282), .A2(n427), .B1(n95), .B2(n284), .ZN(n3276) );
  OAI22_X1 U304 ( .A1(n7119), .A2(n428), .B1(n95), .B2(n287), .ZN(n3277) );
  OAI22_X1 U305 ( .A1(n288), .A2(n4881), .B1(n95), .B2(n289), .ZN(n3278) );
  OAI22_X1 U306 ( .A1(n290), .A2(n4849), .B1(n95), .B2(n291), .ZN(n3279) );
  OAI22_X1 U307 ( .A1(n292), .A2(n429), .B1(n95), .B2(n294), .ZN(n3280) );
  OAI22_X1 U309 ( .A1(n295), .A2(n430), .B1(n95), .B2(n297), .ZN(n3281) );
  OAI22_X1 U311 ( .A1(n298), .A2(n431), .B1(n95), .B2(n300), .ZN(n3282) );
  OAI22_X1 U312 ( .A1(n6558), .A2(n432), .B1(n95), .B2(n7076), .ZN(n3283) );
  OAI22_X1 U314 ( .A1(n304), .A2(n4689), .B1(n95), .B2(n7113), .ZN(n3284) );
  OAI22_X1 U315 ( .A1(n7112), .A2(n4657), .B1(n95), .B2(n307), .ZN(n3285) );
  OAI22_X1 U316 ( .A1(n308), .A2(n433), .B1(n95), .B2(n310), .ZN(n3286) );
  OAI22_X1 U317 ( .A1(n7074), .A2(n434), .B1(n95), .B2(n313), .ZN(n3287) );
  OAI22_X1 U318 ( .A1(n314), .A2(n435), .B1(n95), .B2(n7210), .ZN(n3288) );
  OAI22_X1 U319 ( .A1(n317), .A2(n436), .B1(n95), .B2(n7209), .ZN(n3289) );
  OAI221_X1 U321 ( .B1(n5814), .B2(n320), .C1(n5745), .C2(n5581), .A(n321), 
        .ZN(n413) );
  OAI22_X1 U322 ( .A1(n5581), .A2(net55844), .B1(n94), .B2(net55904), .ZN(
        n3290) );
  INV_X1 U323 ( .A(n412), .ZN(n94) );
  OAI222_X1 U324 ( .A1(n437), .A2(n323), .B1(n6247), .B2(n402), .C1(n438), 
        .C2(n322), .ZN(n412) );
  INV_X1 U325 ( .A(n6250), .ZN(n438) );
  INV_X1 U326 ( .A(n6249), .ZN(n437) );
  OAI221_X1 U327 ( .B1(n357), .B2(n439), .C1(n6262), .C2(n359), .A(n440), .ZN(
        n3291) );
  AOI22_X1 U328 ( .A1(\Mcontrol/bvgen/d_curr_pc[20] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [20]), .B2(n362), .ZN(n440) );
  OAI222_X1 U329 ( .A1(n364), .A2(n441), .B1(n366), .B2(n442), .C1(net55848), 
        .C2(n439), .ZN(n3292) );
  OAI22_X1 U331 ( .A1(net55886), .A2(n442), .B1(net55830), .B2(n441), .ZN(
        n3293) );
  INV_X1 U334 ( .A(n443), .ZN(n3294) );
  AOI22_X1 U335 ( .A1(n7189), .A2(\Mcontrol/f_currpc[20] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[20] ), .ZN(n443) );
  INV_X1 U336 ( .A(n444), .ZN(n3295) );
  OAI221_X1 U338 ( .B1(n445), .B2(n214), .C1(\Mpath/the_alu/N44 ), .C2(
        net55858), .A(n446), .ZN(n3296) );
  AOI222_X1 U339 ( .A1(n197), .A2(n101), .B1(n192), .B2(n447), .C1(n195), .C2(
        n448), .ZN(n446) );
  OAI221_X1 U340 ( .B1(n99), .B2(n232), .C1(\Mpath/the_alu/N43 ), .C2(net55860), .A(n449), .ZN(n3297) );
  AOI22_X1 U341 ( .A1(n6556), .A2(n447), .B1(n6560), .B2(n450), .ZN(n449) );
  OAI22_X1 U342 ( .A1(n237), .A2(n451), .B1(n99), .B2(n239), .ZN(n3298) );
  OAI22_X1 U343 ( .A1(n240), .A2(n452), .B1(n99), .B2(n7318), .ZN(n3299) );
  OAI22_X1 U344 ( .A1(n243), .A2(n453), .B1(n99), .B2(n7370), .ZN(n3300) );
  OAI22_X1 U346 ( .A1(n246), .A2(n454), .B1(n99), .B2(n248), .ZN(n3301) );
  OAI22_X1 U347 ( .A1(n249), .A2(n455), .B1(n99), .B2(n251), .ZN(n3302) );
  OAI22_X1 U348 ( .A1(n252), .A2(n456), .B1(n99), .B2(n7271), .ZN(n3303) );
  OAI22_X1 U349 ( .A1(n255), .A2(n457), .B1(n99), .B2(n257), .ZN(n3304) );
  OAI22_X1 U351 ( .A1(n258), .A2(n458), .B1(n99), .B2(n7117), .ZN(n3305) );
  OAI22_X1 U352 ( .A1(n7115), .A2(n5234), .B1(n99), .B2(n262), .ZN(n3306) );
  OAI22_X1 U353 ( .A1(n263), .A2(n5202), .B1(n99), .B2(n7158), .ZN(n3307) );
  OAI22_X1 U354 ( .A1(n6895), .A2(n459), .B1(n99), .B2(n6898), .ZN(n3308) );
  OAI22_X1 U355 ( .A1(n268), .A2(n5138), .B1(n99), .B2(n269), .ZN(n3309) );
  OAI22_X1 U356 ( .A1(n270), .A2(n5106), .B1(n99), .B2(n271), .ZN(n3310) );
  OAI22_X1 U357 ( .A1(n272), .A2(n460), .B1(n99), .B2(n274), .ZN(n3311) );
  OAI22_X1 U358 ( .A1(n275), .A2(n461), .B1(n99), .B2(n7363), .ZN(n3312) );
  OAI22_X1 U359 ( .A1(n278), .A2(n5010), .B1(n99), .B2(n7276), .ZN(n3313) );
  OAI22_X1 U360 ( .A1(n7122), .A2(n4978), .B1(n99), .B2(n281), .ZN(n3314) );
  OAI22_X1 U361 ( .A1(n282), .A2(n462), .B1(n99), .B2(n284), .ZN(n3315) );
  OAI22_X1 U362 ( .A1(n7119), .A2(n463), .B1(n99), .B2(n287), .ZN(n3316) );
  OAI22_X1 U363 ( .A1(n288), .A2(n4882), .B1(n99), .B2(n289), .ZN(n3317) );
  OAI22_X1 U364 ( .A1(n290), .A2(n4850), .B1(n99), .B2(n291), .ZN(n3318) );
  OAI22_X1 U365 ( .A1(n292), .A2(n464), .B1(n99), .B2(n294), .ZN(n3319) );
  OAI22_X1 U367 ( .A1(n295), .A2(n465), .B1(n99), .B2(n297), .ZN(n3320) );
  OAI22_X1 U369 ( .A1(n298), .A2(n466), .B1(n99), .B2(n300), .ZN(n3321) );
  OAI22_X1 U370 ( .A1(n6558), .A2(n467), .B1(n99), .B2(n7076), .ZN(n3322) );
  OAI22_X1 U372 ( .A1(n304), .A2(n4690), .B1(n99), .B2(n7113), .ZN(n3323) );
  OAI22_X1 U373 ( .A1(n7112), .A2(n4658), .B1(n99), .B2(n307), .ZN(n3324) );
  OAI22_X1 U374 ( .A1(n308), .A2(n468), .B1(n99), .B2(n310), .ZN(n3325) );
  OAI22_X1 U375 ( .A1(n7074), .A2(n469), .B1(n99), .B2(n313), .ZN(n3326) );
  OAI22_X1 U376 ( .A1(n314), .A2(n470), .B1(n99), .B2(n7210), .ZN(n3327) );
  OAI22_X1 U377 ( .A1(n317), .A2(n471), .B1(n99), .B2(n7209), .ZN(n3328) );
  OAI221_X1 U379 ( .B1(n5824), .B2(n320), .C1(n5745), .C2(n5584), .A(n321), 
        .ZN(n448) );
  OAI22_X1 U380 ( .A1(n5584), .A2(net55844), .B1(n98), .B2(net55904), .ZN(
        n3329) );
  INV_X1 U381 ( .A(n447), .ZN(n98) );
  OAI222_X1 U382 ( .A1(n472), .A2(n323), .B1(n6263), .B2(n402), .C1(n473), 
        .C2(n322), .ZN(n447) );
  INV_X1 U383 ( .A(n6266), .ZN(n473) );
  INV_X1 U384 ( .A(n6265), .ZN(n472) );
  OAI221_X1 U385 ( .B1(n357), .B2(n474), .C1(n6275), .C2(n359), .A(n475), .ZN(
        n3330) );
  AOI22_X1 U386 ( .A1(\Mcontrol/bvgen/d_curr_pc[19] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [19]), .B2(n362), .ZN(n475) );
  OAI222_X1 U387 ( .A1(n364), .A2(n476), .B1(n366), .B2(n477), .C1(net55848), 
        .C2(n474), .ZN(n3331) );
  OAI22_X1 U389 ( .A1(net55886), .A2(n477), .B1(net55830), .B2(n476), .ZN(
        n3332) );
  INV_X1 U392 ( .A(n478), .ZN(n3333) );
  AOI22_X1 U393 ( .A1(n7189), .A2(\Mcontrol/f_currpc[19] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[19] ), .ZN(n478) );
  INV_X1 U394 ( .A(n479), .ZN(n3334) );
  AOI221_X1 U395 ( .B1(n371), .B2(\Mcontrol/f_currpc[19] ), .C1(
        I_ADDR_OUTBUS[19]), .C2(n372), .A(n373), .ZN(n479) );
  OAI221_X1 U396 ( .B1(n480), .B2(n214), .C1(\Mpath/the_alu/N46 ), .C2(
        net55860), .A(n481), .ZN(n3335) );
  AOI222_X1 U397 ( .A1(n197), .A2(n105), .B1(n192), .B2(n482), .C1(n195), .C2(
        n483), .ZN(n481) );
  INV_X1 U398 ( .A(break_code[19]), .ZN(n480) );
  OAI221_X1 U399 ( .B1(n103), .B2(n232), .C1(\Mpath/the_alu/N45 ), .C2(
        net55860), .A(n484), .ZN(n3336) );
  AOI22_X1 U400 ( .A1(n6556), .A2(n482), .B1(n6560), .B2(n485), .ZN(n484) );
  OAI22_X1 U401 ( .A1(n237), .A2(n486), .B1(n103), .B2(n239), .ZN(n3337) );
  OAI22_X1 U402 ( .A1(n240), .A2(n487), .B1(n103), .B2(n7318), .ZN(n3338) );
  OAI22_X1 U403 ( .A1(n243), .A2(n488), .B1(n103), .B2(n7370), .ZN(n3339) );
  OAI22_X1 U405 ( .A1(n246), .A2(n489), .B1(n103), .B2(n248), .ZN(n3340) );
  OAI22_X1 U406 ( .A1(n249), .A2(n490), .B1(n103), .B2(n251), .ZN(n3341) );
  OAI22_X1 U407 ( .A1(n252), .A2(n491), .B1(n103), .B2(n7271), .ZN(n3342) );
  OAI22_X1 U408 ( .A1(n255), .A2(n492), .B1(n103), .B2(n257), .ZN(n3343) );
  OAI22_X1 U410 ( .A1(n258), .A2(n493), .B1(n103), .B2(n7117), .ZN(n3344) );
  OAI22_X1 U411 ( .A1(n7115), .A2(n5236), .B1(n103), .B2(n262), .ZN(n3345) );
  OAI22_X1 U412 ( .A1(n263), .A2(n5204), .B1(n103), .B2(n7158), .ZN(n3346) );
  OAI22_X1 U413 ( .A1(n6895), .A2(n494), .B1(n103), .B2(n6898), .ZN(n3347) );
  OAI22_X1 U414 ( .A1(n268), .A2(n5140), .B1(n103), .B2(n269), .ZN(n3348) );
  OAI22_X1 U415 ( .A1(n270), .A2(n5108), .B1(n103), .B2(n271), .ZN(n3349) );
  OAI22_X1 U416 ( .A1(n272), .A2(n495), .B1(n103), .B2(n274), .ZN(n3350) );
  OAI22_X1 U417 ( .A1(n275), .A2(n496), .B1(n103), .B2(n7363), .ZN(n3351) );
  OAI22_X1 U418 ( .A1(n278), .A2(n5012), .B1(n103), .B2(n7276), .ZN(n3352) );
  OAI22_X1 U419 ( .A1(n7122), .A2(n4980), .B1(n103), .B2(n281), .ZN(n3353) );
  OAI22_X1 U420 ( .A1(n282), .A2(n497), .B1(n103), .B2(n284), .ZN(n3354) );
  OAI22_X1 U421 ( .A1(n7119), .A2(n498), .B1(n103), .B2(n287), .ZN(n3355) );
  OAI22_X1 U422 ( .A1(n288), .A2(n4884), .B1(n103), .B2(n289), .ZN(n3356) );
  OAI22_X1 U423 ( .A1(n290), .A2(n4852), .B1(n103), .B2(n291), .ZN(n3357) );
  OAI22_X1 U424 ( .A1(n292), .A2(n499), .B1(n103), .B2(n294), .ZN(n3358) );
  OAI22_X1 U426 ( .A1(n295), .A2(n500), .B1(n103), .B2(n297), .ZN(n3359) );
  OAI22_X1 U428 ( .A1(n298), .A2(n501), .B1(n103), .B2(n300), .ZN(n3360) );
  OAI22_X1 U429 ( .A1(n6559), .A2(n502), .B1(n103), .B2(n7076), .ZN(n3361) );
  OAI22_X1 U431 ( .A1(n304), .A2(n4692), .B1(n103), .B2(n7113), .ZN(n3362) );
  OAI22_X1 U432 ( .A1(n7112), .A2(n4660), .B1(n103), .B2(n307), .ZN(n3363) );
  OAI22_X1 U433 ( .A1(n308), .A2(n503), .B1(n103), .B2(n310), .ZN(n3364) );
  OAI22_X1 U434 ( .A1(n7074), .A2(n504), .B1(n103), .B2(n313), .ZN(n3365) );
  OAI22_X1 U435 ( .A1(n314), .A2(n505), .B1(n103), .B2(n7210), .ZN(n3366) );
  OAI22_X1 U436 ( .A1(n317), .A2(n506), .B1(n103), .B2(n7209), .ZN(n3367) );
  OAI221_X1 U438 ( .B1(n5834), .B2(n320), .C1(n5745), .C2(n5590), .A(n321), 
        .ZN(n483) );
  OAI22_X1 U439 ( .A1(n5590), .A2(net55844), .B1(n102), .B2(net55902), .ZN(
        n3368) );
  INV_X1 U440 ( .A(n482), .ZN(n102) );
  OAI222_X1 U441 ( .A1(n507), .A2(n323), .B1(n6276), .B2(n402), .C1(n508), 
        .C2(n322), .ZN(n482) );
  INV_X1 U442 ( .A(n6279), .ZN(n508) );
  INV_X1 U443 ( .A(n6278), .ZN(n507) );
  OAI221_X1 U444 ( .B1(n357), .B2(n509), .C1(n6290), .C2(n359), .A(n510), .ZN(
        n3369) );
  AOI22_X1 U445 ( .A1(\Mcontrol/bvgen/d_curr_pc[18] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [18]), .B2(n362), .ZN(n510) );
  OAI222_X1 U446 ( .A1(n364), .A2(n511), .B1(n366), .B2(n512), .C1(net55846), 
        .C2(n509), .ZN(n3370) );
  OAI22_X1 U448 ( .A1(net55880), .A2(n512), .B1(net55832), .B2(n511), .ZN(
        n3371) );
  INV_X1 U451 ( .A(n513), .ZN(n3372) );
  AOI22_X1 U452 ( .A1(n7189), .A2(\Mcontrol/f_currpc[18] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[18] ), .ZN(n513) );
  INV_X1 U453 ( .A(n514), .ZN(n3373) );
  AOI221_X1 U454 ( .B1(n371), .B2(\Mcontrol/f_currpc[18] ), .C1(n372), .C2(
        n7873), .A(n373), .ZN(n514) );
  OAI221_X1 U455 ( .B1(n515), .B2(n214), .C1(\Mpath/the_alu/N48 ), .C2(
        net55860), .A(n516), .ZN(n3374) );
  AOI222_X1 U456 ( .A1(n197), .A2(n109), .B1(n192), .B2(n517), .C1(n195), .C2(
        n518), .ZN(n516) );
  INV_X1 U457 ( .A(break_code[18]), .ZN(n515) );
  OAI221_X1 U458 ( .B1(n107), .B2(n232), .C1(\Mpath/the_alu/N47 ), .C2(
        net55860), .A(n519), .ZN(n3375) );
  AOI22_X1 U459 ( .A1(n6556), .A2(n517), .B1(n6560), .B2(n520), .ZN(n519) );
  OAI22_X1 U460 ( .A1(n237), .A2(n521), .B1(n107), .B2(n239), .ZN(n3376) );
  OAI22_X1 U461 ( .A1(n240), .A2(n522), .B1(n107), .B2(n7318), .ZN(n3377) );
  OAI22_X1 U462 ( .A1(n243), .A2(n523), .B1(n107), .B2(n7370), .ZN(n3378) );
  OAI22_X1 U464 ( .A1(n246), .A2(n524), .B1(n107), .B2(n248), .ZN(n3379) );
  OAI22_X1 U465 ( .A1(n249), .A2(n525), .B1(n107), .B2(n251), .ZN(n3380) );
  OAI22_X1 U466 ( .A1(n252), .A2(n526), .B1(n107), .B2(n7271), .ZN(n3381) );
  OAI22_X1 U467 ( .A1(n255), .A2(n527), .B1(n107), .B2(n257), .ZN(n3382) );
  OAI22_X1 U469 ( .A1(n258), .A2(n528), .B1(n107), .B2(n7117), .ZN(n3383) );
  OAI22_X1 U470 ( .A1(n7115), .A2(n5237), .B1(n107), .B2(n262), .ZN(n3384) );
  OAI22_X1 U471 ( .A1(n263), .A2(n5205), .B1(n107), .B2(n7158), .ZN(n3385) );
  OAI22_X1 U472 ( .A1(n6897), .A2(n529), .B1(n107), .B2(n6898), .ZN(n3386) );
  OAI22_X1 U473 ( .A1(n268), .A2(n5141), .B1(n107), .B2(n269), .ZN(n3387) );
  OAI22_X1 U474 ( .A1(n270), .A2(n5109), .B1(n107), .B2(n271), .ZN(n3388) );
  OAI22_X1 U475 ( .A1(n272), .A2(n530), .B1(n107), .B2(n274), .ZN(n3389) );
  OAI22_X1 U476 ( .A1(n275), .A2(n531), .B1(n107), .B2(n7363), .ZN(n3390) );
  OAI22_X1 U477 ( .A1(n278), .A2(n5013), .B1(n107), .B2(n7276), .ZN(n3391) );
  OAI22_X1 U478 ( .A1(n7122), .A2(n4981), .B1(n107), .B2(n281), .ZN(n3392) );
  OAI22_X1 U479 ( .A1(n282), .A2(n532), .B1(n107), .B2(n284), .ZN(n3393) );
  OAI22_X1 U480 ( .A1(n7119), .A2(n533), .B1(n107), .B2(n287), .ZN(n3394) );
  OAI22_X1 U481 ( .A1(n288), .A2(n4885), .B1(n107), .B2(n289), .ZN(n3395) );
  OAI22_X1 U482 ( .A1(n290), .A2(n4853), .B1(n107), .B2(n291), .ZN(n3396) );
  OAI22_X1 U483 ( .A1(n292), .A2(n534), .B1(n107), .B2(n294), .ZN(n3397) );
  OAI22_X1 U485 ( .A1(n295), .A2(n535), .B1(n107), .B2(n297), .ZN(n3398) );
  OAI22_X1 U487 ( .A1(n298), .A2(n536), .B1(n107), .B2(n300), .ZN(n3399) );
  OAI22_X1 U488 ( .A1(n6559), .A2(n537), .B1(n107), .B2(n7076), .ZN(n3400) );
  OAI22_X1 U490 ( .A1(n304), .A2(n4693), .B1(n107), .B2(n7113), .ZN(n3401) );
  OAI22_X1 U491 ( .A1(n7112), .A2(n4661), .B1(n107), .B2(n307), .ZN(n3402) );
  OAI22_X1 U492 ( .A1(n308), .A2(n538), .B1(n107), .B2(n310), .ZN(n3403) );
  OAI22_X1 U493 ( .A1(n7074), .A2(n539), .B1(n107), .B2(n313), .ZN(n3404) );
  OAI22_X1 U494 ( .A1(n314), .A2(n540), .B1(n107), .B2(n7210), .ZN(n3405) );
  OAI22_X1 U495 ( .A1(n317), .A2(n541), .B1(n107), .B2(n7209), .ZN(n3406) );
  OAI221_X1 U497 ( .B1(n5859), .B2(n320), .C1(n5745), .C2(n5593), .A(n321), 
        .ZN(n518) );
  OAI22_X1 U498 ( .A1(n5593), .A2(net55842), .B1(n106), .B2(net55900), .ZN(
        n3407) );
  INV_X1 U499 ( .A(n517), .ZN(n106) );
  OAI222_X1 U500 ( .A1(n542), .A2(n323), .B1(n6291), .B2(n402), .C1(n543), 
        .C2(n322), .ZN(n517) );
  INV_X1 U501 ( .A(n6294), .ZN(n543) );
  INV_X1 U502 ( .A(n6293), .ZN(n542) );
  OAI221_X1 U503 ( .B1(n357), .B2(n544), .C1(n6304), .C2(n359), .A(n545), .ZN(
        n3408) );
  AOI22_X1 U504 ( .A1(\Mcontrol/bvgen/d_curr_pc[17] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [17]), .B2(n362), .ZN(n545) );
  OAI222_X1 U505 ( .A1(n364), .A2(n546), .B1(n366), .B2(n547), .C1(net55848), 
        .C2(n544), .ZN(n3409) );
  OAI22_X1 U507 ( .A1(net55878), .A2(n547), .B1(net55830), .B2(n546), .ZN(
        n3410) );
  INV_X1 U510 ( .A(n548), .ZN(n3411) );
  AOI22_X1 U511 ( .A1(n7189), .A2(\Mcontrol/f_currpc[17] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[17] ), .ZN(n548) );
  INV_X1 U512 ( .A(n549), .ZN(n3412) );
  AOI221_X1 U513 ( .B1(n371), .B2(\Mcontrol/f_currpc[17] ), .C1(n372), .C2(
        n7874), .A(n373), .ZN(n549) );
  OAI221_X1 U514 ( .B1(n550), .B2(n214), .C1(\Mpath/the_alu/N50 ), .C2(
        net55860), .A(n551), .ZN(n3413) );
  AOI222_X1 U515 ( .A1(n197), .A2(n113), .B1(n192), .B2(n552), .C1(n195), .C2(
        n553), .ZN(n551) );
  INV_X1 U516 ( .A(break_code[17]), .ZN(n550) );
  OAI221_X1 U517 ( .B1(n111), .B2(n232), .C1(\Mpath/the_alu/N49 ), .C2(
        net55860), .A(n554), .ZN(n3414) );
  AOI22_X1 U518 ( .A1(n6556), .A2(n552), .B1(n6560), .B2(n555), .ZN(n554) );
  OAI22_X1 U519 ( .A1(n237), .A2(n556), .B1(n111), .B2(n239), .ZN(n3415) );
  OAI22_X1 U520 ( .A1(n240), .A2(n557), .B1(n111), .B2(n7318), .ZN(n3416) );
  OAI22_X1 U521 ( .A1(n243), .A2(n558), .B1(n111), .B2(n7370), .ZN(n3417) );
  OAI22_X1 U523 ( .A1(n246), .A2(n559), .B1(n111), .B2(n248), .ZN(n3418) );
  OAI22_X1 U524 ( .A1(n249), .A2(n560), .B1(n111), .B2(n251), .ZN(n3419) );
  OAI22_X1 U525 ( .A1(n252), .A2(n561), .B1(n111), .B2(n7271), .ZN(n3420) );
  OAI22_X1 U526 ( .A1(n255), .A2(n562), .B1(n111), .B2(n257), .ZN(n3421) );
  OAI22_X1 U528 ( .A1(n258), .A2(n563), .B1(n111), .B2(n7117), .ZN(n3422) );
  OAI22_X1 U529 ( .A1(n7115), .A2(n5238), .B1(n111), .B2(n262), .ZN(n3423) );
  OAI22_X1 U530 ( .A1(n263), .A2(n5206), .B1(n111), .B2(n7158), .ZN(n3424) );
  OAI22_X1 U531 ( .A1(n6896), .A2(n564), .B1(n111), .B2(n6898), .ZN(n3425) );
  OAI22_X1 U532 ( .A1(n268), .A2(n5142), .B1(n111), .B2(n269), .ZN(n3426) );
  OAI22_X1 U533 ( .A1(n270), .A2(n5110), .B1(n111), .B2(n271), .ZN(n3427) );
  OAI22_X1 U534 ( .A1(n272), .A2(n565), .B1(n111), .B2(n274), .ZN(n3428) );
  OAI22_X1 U535 ( .A1(n275), .A2(n566), .B1(n111), .B2(n7363), .ZN(n3429) );
  OAI22_X1 U536 ( .A1(n278), .A2(n5014), .B1(n111), .B2(n7276), .ZN(n3430) );
  OAI22_X1 U537 ( .A1(n7122), .A2(n4982), .B1(n111), .B2(n281), .ZN(n3431) );
  OAI22_X1 U538 ( .A1(n282), .A2(n567), .B1(n111), .B2(n284), .ZN(n3432) );
  OAI22_X1 U539 ( .A1(n7119), .A2(n568), .B1(n111), .B2(n287), .ZN(n3433) );
  OAI22_X1 U540 ( .A1(n288), .A2(n4886), .B1(n111), .B2(n289), .ZN(n3434) );
  OAI22_X1 U541 ( .A1(n290), .A2(n4854), .B1(n111), .B2(n291), .ZN(n3435) );
  OAI22_X1 U542 ( .A1(n292), .A2(n569), .B1(n111), .B2(n294), .ZN(n3436) );
  OAI22_X1 U544 ( .A1(n295), .A2(n570), .B1(n111), .B2(n297), .ZN(n3437) );
  OAI22_X1 U546 ( .A1(n298), .A2(n571), .B1(n111), .B2(n300), .ZN(n3438) );
  OAI22_X1 U547 ( .A1(n6558), .A2(n572), .B1(n111), .B2(n7076), .ZN(n3439) );
  OAI22_X1 U549 ( .A1(n304), .A2(n4694), .B1(n111), .B2(n7113), .ZN(n3440) );
  OAI22_X1 U550 ( .A1(n7112), .A2(n4662), .B1(n111), .B2(n307), .ZN(n3441) );
  OAI22_X1 U551 ( .A1(n308), .A2(n573), .B1(n111), .B2(n310), .ZN(n3442) );
  OAI22_X1 U552 ( .A1(n7074), .A2(n574), .B1(n111), .B2(n313), .ZN(n3443) );
  OAI22_X1 U553 ( .A1(n314), .A2(n575), .B1(n111), .B2(n7210), .ZN(n3444) );
  OAI22_X1 U554 ( .A1(n317), .A2(n576), .B1(n111), .B2(n7209), .ZN(n3445) );
  OAI221_X1 U556 ( .B1(n5940), .B2(n320), .C1(n5745), .C2(n5596), .A(n321), 
        .ZN(n553) );
  OAI22_X1 U557 ( .A1(n5596), .A2(net55846), .B1(n110), .B2(net55904), .ZN(
        n3446) );
  INV_X1 U558 ( .A(n552), .ZN(n110) );
  OAI222_X1 U559 ( .A1(n577), .A2(n323), .B1(n6305), .B2(n402), .C1(n578), 
        .C2(n322), .ZN(n552) );
  INV_X1 U560 ( .A(n6308), .ZN(n578) );
  INV_X1 U561 ( .A(n6307), .ZN(n577) );
  OAI221_X1 U562 ( .B1(n357), .B2(n579), .C1(n6316), .C2(n359), .A(n580), .ZN(
        n3447) );
  AOI22_X1 U563 ( .A1(\Mcontrol/bvgen/d_curr_pc[16] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [16]), .B2(n362), .ZN(n580) );
  OAI222_X1 U564 ( .A1(n364), .A2(n581), .B1(n366), .B2(n582), .C1(net55848), 
        .C2(n579), .ZN(n3448) );
  OAI22_X1 U566 ( .A1(net55878), .A2(n582), .B1(net55832), .B2(n581), .ZN(
        n3449) );
  INV_X1 U569 ( .A(n583), .ZN(n3450) );
  AOI22_X1 U570 ( .A1(n7189), .A2(\Mcontrol/f_currpc[16] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[16] ), .ZN(n583) );
  INV_X1 U571 ( .A(n584), .ZN(n3451) );
  AOI221_X1 U572 ( .B1(n371), .B2(\Mcontrol/f_currpc[16] ), .C1(n372), .C2(
        n7875), .A(n373), .ZN(n584) );
  OAI221_X1 U573 ( .B1(n585), .B2(n214), .C1(\Mpath/the_alu/N52 ), .C2(
        net55858), .A(n586), .ZN(n3452) );
  AOI222_X1 U574 ( .A1(n197), .A2(n117), .B1(n192), .B2(n587), .C1(n195), .C2(
        n588), .ZN(n586) );
  INV_X1 U575 ( .A(break_code[16]), .ZN(n585) );
  OAI221_X1 U576 ( .B1(n115), .B2(n232), .C1(\Mpath/the_alu/N51 ), .C2(
        net55860), .A(n589), .ZN(n3453) );
  AOI22_X1 U577 ( .A1(n6556), .A2(n587), .B1(n6560), .B2(n590), .ZN(n589) );
  OAI22_X1 U578 ( .A1(n237), .A2(n591), .B1(n115), .B2(n239), .ZN(n3454) );
  OAI22_X1 U579 ( .A1(n240), .A2(n592), .B1(n115), .B2(n7318), .ZN(n3455) );
  OAI22_X1 U580 ( .A1(n243), .A2(n593), .B1(n115), .B2(n7370), .ZN(n3456) );
  OAI22_X1 U582 ( .A1(n246), .A2(n594), .B1(n115), .B2(n248), .ZN(n3457) );
  OAI22_X1 U583 ( .A1(n249), .A2(n595), .B1(n115), .B2(n251), .ZN(n3458) );
  OAI22_X1 U584 ( .A1(n252), .A2(n596), .B1(n115), .B2(n7271), .ZN(n3459) );
  OAI22_X1 U585 ( .A1(n255), .A2(n597), .B1(n115), .B2(n257), .ZN(n3460) );
  OAI22_X1 U587 ( .A1(n258), .A2(n598), .B1(n115), .B2(n7117), .ZN(n3461) );
  OAI22_X1 U588 ( .A1(n7115), .A2(n5239), .B1(n115), .B2(n262), .ZN(n3462) );
  OAI22_X1 U589 ( .A1(n263), .A2(n5207), .B1(n115), .B2(n7158), .ZN(n3463) );
  OAI22_X1 U590 ( .A1(n6897), .A2(n599), .B1(n115), .B2(n6898), .ZN(n3464) );
  OAI22_X1 U591 ( .A1(n268), .A2(n5143), .B1(n115), .B2(n269), .ZN(n3465) );
  OAI22_X1 U592 ( .A1(n270), .A2(n5111), .B1(n115), .B2(n271), .ZN(n3466) );
  OAI22_X1 U593 ( .A1(n272), .A2(n600), .B1(n115), .B2(n274), .ZN(n3467) );
  OAI22_X1 U594 ( .A1(n275), .A2(n601), .B1(n115), .B2(n7363), .ZN(n3468) );
  OAI22_X1 U595 ( .A1(n278), .A2(n5015), .B1(n115), .B2(n7276), .ZN(n3469) );
  OAI22_X1 U596 ( .A1(n7122), .A2(n4983), .B1(n115), .B2(n281), .ZN(n3470) );
  OAI22_X1 U597 ( .A1(n282), .A2(n602), .B1(n115), .B2(n284), .ZN(n3471) );
  OAI22_X1 U598 ( .A1(n7119), .A2(n603), .B1(n115), .B2(n287), .ZN(n3472) );
  OAI22_X1 U599 ( .A1(n288), .A2(n4887), .B1(n115), .B2(n289), .ZN(n3473) );
  OAI22_X1 U600 ( .A1(n290), .A2(n4855), .B1(n115), .B2(n291), .ZN(n3474) );
  OAI22_X1 U601 ( .A1(n292), .A2(n604), .B1(n115), .B2(n294), .ZN(n3475) );
  OAI22_X1 U603 ( .A1(n295), .A2(n605), .B1(n115), .B2(n297), .ZN(n3476) );
  OAI22_X1 U605 ( .A1(n298), .A2(n606), .B1(n115), .B2(n300), .ZN(n3477) );
  OAI22_X1 U606 ( .A1(n6558), .A2(n607), .B1(n115), .B2(n7076), .ZN(n3478) );
  OAI22_X1 U608 ( .A1(n304), .A2(n4695), .B1(n115), .B2(n7113), .ZN(n3479) );
  OAI22_X1 U609 ( .A1(n7112), .A2(n4663), .B1(n115), .B2(n307), .ZN(n3480) );
  OAI22_X1 U610 ( .A1(n308), .A2(n608), .B1(n115), .B2(n310), .ZN(n3481) );
  OAI22_X1 U611 ( .A1(n7074), .A2(n609), .B1(n115), .B2(n313), .ZN(n3482) );
  OAI22_X1 U612 ( .A1(n314), .A2(n610), .B1(n115), .B2(n7210), .ZN(n3483) );
  OAI22_X1 U613 ( .A1(n317), .A2(n611), .B1(n115), .B2(n7209), .ZN(n3484) );
  OAI221_X1 U615 ( .B1(n5961), .B2(n320), .C1(n5745), .C2(n5599), .A(n321), 
        .ZN(n588) );
  OAI22_X1 U616 ( .A1(n5599), .A2(net55846), .B1(n114), .B2(net55900), .ZN(
        n3485) );
  INV_X1 U617 ( .A(n587), .ZN(n114) );
  OAI222_X1 U618 ( .A1(n612), .A2(n323), .B1(n6317), .B2(n402), .C1(n613), 
        .C2(n322), .ZN(n587) );
  INV_X1 U619 ( .A(n6320), .ZN(n613) );
  INV_X1 U620 ( .A(n6319), .ZN(n612) );
  OAI221_X1 U621 ( .B1(n357), .B2(n614), .C1(n359), .C2(n615), .A(n616), .ZN(
        n3486) );
  AOI22_X1 U622 ( .A1(\Mcontrol/bvgen/d_curr_pc[15] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [15]), .B2(n362), .ZN(n616) );
  OAI222_X1 U624 ( .A1(n364), .A2(n617), .B1(n366), .B2(n618), .C1(net55848), 
        .C2(n614), .ZN(n3487) );
  OAI22_X1 U626 ( .A1(net55878), .A2(n618), .B1(net55832), .B2(n617), .ZN(
        n3488) );
  INV_X1 U629 ( .A(n619), .ZN(n3489) );
  AOI22_X1 U630 ( .A1(n7189), .A2(\Mcontrol/f_currpc[15] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[15] ), .ZN(n619) );
  INV_X1 U631 ( .A(n620), .ZN(n3490) );
  AOI221_X1 U632 ( .B1(n371), .B2(\Mcontrol/f_currpc[15] ), .C1(n372), .C2(
        n7876), .A(n373), .ZN(n620) );
  OAI221_X1 U633 ( .B1(n621), .B2(n214), .C1(\Mpath/the_alu/N54 ), .C2(
        net55856), .A(n622), .ZN(n3491) );
  AOI222_X1 U634 ( .A1(n197), .A2(n121), .B1(n192), .B2(n623), .C1(n195), .C2(
        n624), .ZN(n622) );
  INV_X1 U635 ( .A(break_code[15]), .ZN(n621) );
  OAI22_X1 U636 ( .A1(n5737), .A2(net55916), .B1(net55832), .B2(n625), .ZN(
        n3492) );
  OAI22_X1 U637 ( .A1(n5738), .A2(n626), .B1(n5737), .B2(n627), .ZN(n3493) );
  OAI222_X1 U638 ( .A1(n625), .A2(n628), .B1(n5737), .B2(n629), .C1(n5738), 
        .C2(n359), .ZN(n3494) );
  OAI221_X1 U640 ( .B1(n119), .B2(n232), .C1(\Mpath/the_alu/N53 ), .C2(
        net55856), .A(n630), .ZN(n3495) );
  AOI22_X1 U641 ( .A1(n6556), .A2(n623), .B1(n6560), .B2(n631), .ZN(n630) );
  OAI22_X1 U642 ( .A1(n237), .A2(n632), .B1(n119), .B2(n239), .ZN(n3496) );
  OAI22_X1 U643 ( .A1(n240), .A2(n633), .B1(n119), .B2(n7318), .ZN(n3497) );
  OAI22_X1 U644 ( .A1(n243), .A2(n634), .B1(n119), .B2(n7370), .ZN(n3498) );
  OAI22_X1 U646 ( .A1(n246), .A2(n635), .B1(n119), .B2(n248), .ZN(n3499) );
  OAI22_X1 U647 ( .A1(n249), .A2(n636), .B1(n119), .B2(n251), .ZN(n3500) );
  OAI22_X1 U648 ( .A1(n252), .A2(n637), .B1(n119), .B2(n7271), .ZN(n3501) );
  OAI22_X1 U649 ( .A1(n255), .A2(n638), .B1(n119), .B2(n257), .ZN(n3502) );
  OAI22_X1 U651 ( .A1(n258), .A2(n639), .B1(n119), .B2(n7117), .ZN(n3503) );
  OAI22_X1 U652 ( .A1(n7115), .A2(n5240), .B1(n119), .B2(n262), .ZN(n3504) );
  OAI22_X1 U653 ( .A1(n263), .A2(n5208), .B1(n119), .B2(n7158), .ZN(n3505) );
  OAI22_X1 U654 ( .A1(n6895), .A2(n640), .B1(n119), .B2(n6898), .ZN(n3506) );
  OAI22_X1 U655 ( .A1(n268), .A2(n5144), .B1(n119), .B2(n269), .ZN(n3507) );
  OAI22_X1 U656 ( .A1(n270), .A2(n5112), .B1(n119), .B2(n271), .ZN(n3508) );
  OAI22_X1 U657 ( .A1(n272), .A2(n641), .B1(n119), .B2(n274), .ZN(n3509) );
  OAI22_X1 U658 ( .A1(n275), .A2(n642), .B1(n119), .B2(n7363), .ZN(n3510) );
  OAI22_X1 U659 ( .A1(n278), .A2(n5016), .B1(n119), .B2(n7276), .ZN(n3511) );
  OAI22_X1 U660 ( .A1(n7122), .A2(n4984), .B1(n119), .B2(n281), .ZN(n3512) );
  OAI22_X1 U661 ( .A1(n282), .A2(n643), .B1(n119), .B2(n284), .ZN(n3513) );
  OAI22_X1 U662 ( .A1(n7119), .A2(n644), .B1(n119), .B2(n287), .ZN(n3514) );
  OAI22_X1 U663 ( .A1(n288), .A2(n4888), .B1(n119), .B2(n289), .ZN(n3515) );
  OAI22_X1 U664 ( .A1(n290), .A2(n4856), .B1(n119), .B2(n291), .ZN(n3516) );
  OAI22_X1 U665 ( .A1(n292), .A2(n645), .B1(n119), .B2(n294), .ZN(n3517) );
  OAI22_X1 U667 ( .A1(n295), .A2(n646), .B1(n119), .B2(n297), .ZN(n3518) );
  OAI22_X1 U669 ( .A1(n298), .A2(n647), .B1(n119), .B2(n300), .ZN(n3519) );
  OAI22_X1 U670 ( .A1(n6559), .A2(n648), .B1(n119), .B2(n7076), .ZN(n3520) );
  OAI22_X1 U672 ( .A1(n304), .A2(n4696), .B1(n119), .B2(n7113), .ZN(n3521) );
  OAI22_X1 U673 ( .A1(n7112), .A2(n4664), .B1(n119), .B2(n307), .ZN(n3522) );
  OAI22_X1 U674 ( .A1(n308), .A2(n649), .B1(n119), .B2(n310), .ZN(n3523) );
  OAI22_X1 U675 ( .A1(n7074), .A2(n650), .B1(n119), .B2(n313), .ZN(n3524) );
  OAI22_X1 U676 ( .A1(n314), .A2(n651), .B1(n119), .B2(n7210), .ZN(n3525) );
  OAI22_X1 U677 ( .A1(n317), .A2(n652), .B1(n119), .B2(n7209), .ZN(n3526) );
  OAI211_X1 U679 ( .C1(n5789), .C2(n653), .A(n654), .B(n655), .ZN(n624) );
  AOI22_X1 U680 ( .A1(n656), .A2(n6541), .B1(n657), .B2(n658), .ZN(n655) );
  INV_X1 U681 ( .A(n5602), .ZN(n657) );
  OAI22_X1 U682 ( .A1(n5602), .A2(net55844), .B1(n118), .B2(net55908), .ZN(
        n3527) );
  INV_X1 U683 ( .A(n623), .ZN(n118) );
  OAI222_X1 U684 ( .A1(n659), .A2(n323), .B1(n6329), .B2(n402), .C1(n660), 
        .C2(n322), .ZN(n623) );
  INV_X1 U685 ( .A(n6333), .ZN(n660) );
  INV_X1 U686 ( .A(n6332), .ZN(n659) );
  OAI221_X1 U687 ( .B1(n357), .B2(n661), .C1(n359), .C2(n662), .A(n663), .ZN(
        n3528) );
  AOI22_X1 U688 ( .A1(\Mcontrol/bvgen/d_curr_pc[14] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [14]), .B2(n362), .ZN(n663) );
  OAI222_X1 U690 ( .A1(n364), .A2(n664), .B1(n366), .B2(n665), .C1(net55846), 
        .C2(n661), .ZN(n3529) );
  OAI22_X1 U692 ( .A1(net55878), .A2(n665), .B1(net55832), .B2(n664), .ZN(
        n3530) );
  INV_X1 U695 ( .A(n666), .ZN(n3531) );
  AOI22_X1 U696 ( .A1(n7189), .A2(\Mcontrol/f_currpc[14] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[14] ), .ZN(n666) );
  INV_X1 U697 ( .A(n667), .ZN(n3532) );
  AOI221_X1 U698 ( .B1(n371), .B2(\Mcontrol/f_currpc[14] ), .C1(n372), .C2(
        n7877), .A(n373), .ZN(n667) );
  OAI221_X1 U699 ( .B1(n668), .B2(n214), .C1(\Mpath/the_alu/N56 ), .C2(
        net55858), .A(n669), .ZN(n3533) );
  AOI222_X1 U700 ( .A1(n197), .A2(n125), .B1(n192), .B2(n670), .C1(n195), .C2(
        n671), .ZN(n669) );
  INV_X1 U701 ( .A(break_code[14]), .ZN(n668) );
  OAI221_X1 U702 ( .B1(n672), .B2(n214), .C1(\Mpath/the_alu/N64 ), .C2(
        net55856), .A(n673), .ZN(n3534) );
  AOI222_X1 U703 ( .A1(n197), .A2(n141), .B1(n192), .B2(n674), .C1(n195), .C2(
        n675), .ZN(n673) );
  INV_X1 U704 ( .A(break_code[10]), .ZN(n672) );
  OAI221_X1 U705 ( .B1(n357), .B2(n676), .C1(n359), .C2(n677), .A(n678), .ZN(
        n3535) );
  AOI22_X1 U706 ( .A1(\Mcontrol/bvgen/d_curr_pc[10] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [10]), .B2(n362), .ZN(n678) );
  OAI221_X1 U708 ( .B1(n139), .B2(n232), .C1(\Mpath/the_alu/N63 ), .C2(
        net55856), .A(n679), .ZN(n3536) );
  AOI22_X1 U709 ( .A1(n6556), .A2(n674), .B1(n6560), .B2(n680), .ZN(n679) );
  OAI22_X1 U710 ( .A1(n237), .A2(n681), .B1(n139), .B2(n239), .ZN(n3537) );
  OAI22_X1 U711 ( .A1(n240), .A2(n682), .B1(n139), .B2(n7318), .ZN(n3538) );
  OAI22_X1 U712 ( .A1(n243), .A2(n683), .B1(n139), .B2(n7370), .ZN(n3539) );
  OAI22_X1 U714 ( .A1(n246), .A2(n684), .B1(n139), .B2(n248), .ZN(n3540) );
  OAI22_X1 U715 ( .A1(n249), .A2(n685), .B1(n139), .B2(n251), .ZN(n3541) );
  OAI22_X1 U716 ( .A1(n252), .A2(n686), .B1(n139), .B2(n7271), .ZN(n3542) );
  OAI22_X1 U717 ( .A1(n255), .A2(n687), .B1(n139), .B2(n257), .ZN(n3543) );
  OAI22_X1 U719 ( .A1(n258), .A2(n688), .B1(n139), .B2(n7117), .ZN(n3544) );
  OAI22_X1 U720 ( .A1(n7115), .A2(n5245), .B1(n139), .B2(n262), .ZN(n3545) );
  OAI22_X1 U721 ( .A1(n263), .A2(n5213), .B1(n139), .B2(n7158), .ZN(n3546) );
  OAI22_X1 U722 ( .A1(n6897), .A2(n689), .B1(n139), .B2(n6898), .ZN(n3547) );
  OAI22_X1 U723 ( .A1(n268), .A2(n5149), .B1(n139), .B2(n269), .ZN(n3548) );
  OAI22_X1 U724 ( .A1(n270), .A2(n5117), .B1(n139), .B2(n271), .ZN(n3549) );
  OAI22_X1 U725 ( .A1(n272), .A2(n690), .B1(n139), .B2(n274), .ZN(n3550) );
  OAI22_X1 U726 ( .A1(n275), .A2(n691), .B1(n139), .B2(n7363), .ZN(n3551) );
  OAI22_X1 U727 ( .A1(n278), .A2(n5021), .B1(n139), .B2(n7276), .ZN(n3552) );
  OAI22_X1 U728 ( .A1(n7122), .A2(n4989), .B1(n139), .B2(n281), .ZN(n3553) );
  OAI22_X1 U729 ( .A1(n282), .A2(n692), .B1(n139), .B2(n284), .ZN(n3554) );
  OAI22_X1 U730 ( .A1(n7119), .A2(n693), .B1(n139), .B2(n287), .ZN(n3555) );
  OAI22_X1 U731 ( .A1(n288), .A2(n4893), .B1(n139), .B2(n289), .ZN(n3556) );
  OAI22_X1 U732 ( .A1(n290), .A2(n4861), .B1(n139), .B2(n291), .ZN(n3557) );
  OAI22_X1 U733 ( .A1(n292), .A2(n694), .B1(n139), .B2(n294), .ZN(n3558) );
  OAI22_X1 U735 ( .A1(n295), .A2(n695), .B1(n139), .B2(n297), .ZN(n3559) );
  OAI22_X1 U737 ( .A1(n298), .A2(n696), .B1(n139), .B2(n300), .ZN(n3560) );
  OAI22_X1 U738 ( .A1(n6559), .A2(n697), .B1(n139), .B2(n7076), .ZN(n3561) );
  OAI22_X1 U740 ( .A1(n304), .A2(n4701), .B1(n139), .B2(n7113), .ZN(n3562) );
  OAI22_X1 U741 ( .A1(n7112), .A2(n4669), .B1(n139), .B2(n307), .ZN(n3563) );
  OAI22_X1 U742 ( .A1(n308), .A2(n698), .B1(n139), .B2(n310), .ZN(n3564) );
  OAI22_X1 U743 ( .A1(n7074), .A2(n699), .B1(n139), .B2(n313), .ZN(n3565) );
  OAI22_X1 U744 ( .A1(n314), .A2(n700), .B1(n139), .B2(n7210), .ZN(n3566) );
  OAI22_X1 U745 ( .A1(n317), .A2(n701), .B1(n139), .B2(n7209), .ZN(n3567) );
  OAI211_X1 U747 ( .C1(n5856), .C2(n653), .A(n654), .B(n702), .ZN(n675) );
  AOI22_X1 U748 ( .A1(n656), .A2(n6531), .B1(n703), .B2(n658), .ZN(n702) );
  INV_X1 U749 ( .A(n5617), .ZN(n703) );
  OAI22_X1 U750 ( .A1(n5617), .A2(net55844), .B1(n138), .B2(net55908), .ZN(
        n3568) );
  INV_X1 U751 ( .A(n674), .ZN(n138) );
  OAI222_X1 U752 ( .A1(n704), .A2(n323), .B1(n6391), .B2(n402), .C1(n705), 
        .C2(n322), .ZN(n674) );
  INV_X1 U753 ( .A(n6395), .ZN(n705) );
  INV_X1 U754 ( .A(n6394), .ZN(n704) );
  OAI221_X1 U755 ( .B1(n357), .B2(n706), .C1(n359), .C2(n707), .A(n708), .ZN(
        n3569) );
  AOI22_X1 U756 ( .A1(\Mcontrol/bvgen/d_curr_pc[11] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [11]), .B2(n362), .ZN(n708) );
  OAI222_X1 U758 ( .A1(n364), .A2(n709), .B1(n366), .B2(n710), .C1(net55848), 
        .C2(n706), .ZN(n3570) );
  OAI22_X1 U760 ( .A1(net55878), .A2(n710), .B1(net55830), .B2(n709), .ZN(
        n3571) );
  INV_X1 U763 ( .A(n711), .ZN(n3572) );
  AOI22_X1 U764 ( .A1(n7189), .A2(\Mcontrol/f_currpc[11] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[11] ), .ZN(n711) );
  INV_X1 U765 ( .A(n712), .ZN(n3573) );
  AOI221_X1 U766 ( .B1(n371), .B2(\Mcontrol/f_currpc[11] ), .C1(n372), .C2(
        n7880), .A(n373), .ZN(n712) );
  OAI221_X1 U767 ( .B1(n713), .B2(n214), .C1(\Mpath/the_alu/N62 ), .C2(
        net55858), .A(n714), .ZN(n3574) );
  AOI222_X1 U768 ( .A1(n197), .A2(n137), .B1(n192), .B2(n715), .C1(n195), .C2(
        n716), .ZN(n714) );
  INV_X1 U769 ( .A(break_code[11]), .ZN(n713) );
  OAI221_X1 U770 ( .B1(n135), .B2(n232), .C1(\Mpath/the_alu/N61 ), .C2(
        net55858), .A(n717), .ZN(n3575) );
  AOI22_X1 U771 ( .A1(n6556), .A2(n715), .B1(n6560), .B2(n718), .ZN(n717) );
  OAI22_X1 U772 ( .A1(n237), .A2(n719), .B1(n135), .B2(n239), .ZN(n3576) );
  OAI22_X1 U773 ( .A1(n240), .A2(n720), .B1(n135), .B2(n7318), .ZN(n3577) );
  OAI22_X1 U774 ( .A1(n243), .A2(n721), .B1(n135), .B2(n7370), .ZN(n3578) );
  OAI22_X1 U776 ( .A1(n246), .A2(n722), .B1(n135), .B2(n248), .ZN(n3579) );
  OAI22_X1 U777 ( .A1(n249), .A2(n723), .B1(n135), .B2(n251), .ZN(n3580) );
  OAI22_X1 U778 ( .A1(n252), .A2(n724), .B1(n135), .B2(n7271), .ZN(n3581) );
  OAI22_X1 U779 ( .A1(n255), .A2(n725), .B1(n135), .B2(n257), .ZN(n3582) );
  OAI22_X1 U781 ( .A1(n258), .A2(n726), .B1(n135), .B2(n7117), .ZN(n3583) );
  OAI22_X1 U782 ( .A1(n7115), .A2(n5244), .B1(n135), .B2(n262), .ZN(n3584) );
  OAI22_X1 U783 ( .A1(n263), .A2(n5212), .B1(n135), .B2(n7158), .ZN(n3585) );
  OAI22_X1 U784 ( .A1(n6896), .A2(n727), .B1(n135), .B2(n6898), .ZN(n3586) );
  OAI22_X1 U785 ( .A1(n268), .A2(n5148), .B1(n135), .B2(n269), .ZN(n3587) );
  OAI22_X1 U786 ( .A1(n270), .A2(n5116), .B1(n135), .B2(n271), .ZN(n3588) );
  OAI22_X1 U787 ( .A1(n272), .A2(n728), .B1(n135), .B2(n274), .ZN(n3589) );
  OAI22_X1 U788 ( .A1(n275), .A2(n729), .B1(n135), .B2(n7363), .ZN(n3590) );
  OAI22_X1 U789 ( .A1(n278), .A2(n5020), .B1(n135), .B2(n7276), .ZN(n3591) );
  OAI22_X1 U790 ( .A1(n7122), .A2(n4988), .B1(n135), .B2(n281), .ZN(n3592) );
  OAI22_X1 U791 ( .A1(n282), .A2(n730), .B1(n135), .B2(n284), .ZN(n3593) );
  OAI22_X1 U792 ( .A1(n7119), .A2(n731), .B1(n135), .B2(n287), .ZN(n3594) );
  OAI22_X1 U793 ( .A1(n288), .A2(n4892), .B1(n135), .B2(n289), .ZN(n3595) );
  OAI22_X1 U794 ( .A1(n290), .A2(n4860), .B1(n135), .B2(n291), .ZN(n3596) );
  OAI22_X1 U795 ( .A1(n292), .A2(n732), .B1(n135), .B2(n294), .ZN(n3597) );
  OAI22_X1 U797 ( .A1(n295), .A2(n733), .B1(n135), .B2(n297), .ZN(n3598) );
  OAI22_X1 U799 ( .A1(n298), .A2(n734), .B1(n135), .B2(n300), .ZN(n3599) );
  OAI22_X1 U800 ( .A1(n6558), .A2(n735), .B1(n135), .B2(n7076), .ZN(n3600) );
  OAI22_X1 U802 ( .A1(n304), .A2(n4700), .B1(n135), .B2(n7113), .ZN(n3601) );
  OAI22_X1 U803 ( .A1(n7112), .A2(n4668), .B1(n135), .B2(n307), .ZN(n3602) );
  OAI22_X1 U804 ( .A1(n308), .A2(n736), .B1(n135), .B2(n310), .ZN(n3603) );
  OAI22_X1 U805 ( .A1(n7074), .A2(n737), .B1(n135), .B2(n313), .ZN(n3604) );
  OAI22_X1 U806 ( .A1(n314), .A2(n738), .B1(n135), .B2(n7210), .ZN(n3605) );
  OAI22_X1 U807 ( .A1(n317), .A2(n739), .B1(n135), .B2(n7209), .ZN(n3606) );
  OAI211_X1 U809 ( .C1(n5831), .C2(n653), .A(n654), .B(n740), .ZN(n716) );
  AOI22_X1 U810 ( .A1(n656), .A2(n6533), .B1(n741), .B2(n658), .ZN(n740) );
  INV_X1 U811 ( .A(n5614), .ZN(n741) );
  OAI22_X1 U812 ( .A1(n5614), .A2(net55846), .B1(n134), .B2(net55908), .ZN(
        n3607) );
  INV_X1 U813 ( .A(n715), .ZN(n134) );
  OAI222_X1 U814 ( .A1(n742), .A2(n323), .B1(n6377), .B2(n402), .C1(n743), 
        .C2(n322), .ZN(n715) );
  INV_X1 U815 ( .A(n6381), .ZN(n743) );
  INV_X1 U816 ( .A(n6380), .ZN(n742) );
  OAI221_X1 U817 ( .B1(n357), .B2(n744), .C1(n359), .C2(n745), .A(n746), .ZN(
        n3608) );
  AOI22_X1 U818 ( .A1(\Mcontrol/bvgen/d_curr_pc[12] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [12]), .B2(n362), .ZN(n746) );
  OAI222_X1 U820 ( .A1(n364), .A2(n747), .B1(n366), .B2(n748), .C1(net55850), 
        .C2(n744), .ZN(n3609) );
  OAI22_X1 U822 ( .A1(net55878), .A2(n748), .B1(net55832), .B2(n747), .ZN(
        n3610) );
  INV_X1 U825 ( .A(n749), .ZN(n3611) );
  AOI22_X1 U826 ( .A1(n7189), .A2(\Mcontrol/f_currpc[12] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[12] ), .ZN(n749) );
  INV_X1 U827 ( .A(n750), .ZN(n3612) );
  AOI221_X1 U828 ( .B1(n371), .B2(\Mcontrol/f_currpc[12] ), .C1(n372), .C2(
        n7879), .A(n373), .ZN(n750) );
  OAI221_X1 U829 ( .B1(n751), .B2(n214), .C1(\Mpath/the_alu/N60 ), .C2(
        net55858), .A(n752), .ZN(n3613) );
  AOI222_X1 U830 ( .A1(n197), .A2(n133), .B1(n192), .B2(n753), .C1(n195), .C2(
        n754), .ZN(n752) );
  INV_X1 U831 ( .A(break_code[12]), .ZN(n751) );
  OAI221_X1 U832 ( .B1(n131), .B2(n232), .C1(\Mpath/the_alu/N59 ), .C2(
        net55858), .A(n755), .ZN(n3614) );
  AOI22_X1 U833 ( .A1(n6556), .A2(n753), .B1(n6560), .B2(n756), .ZN(n755) );
  OAI22_X1 U834 ( .A1(n237), .A2(n757), .B1(n131), .B2(n239), .ZN(n3615) );
  OAI22_X1 U835 ( .A1(n240), .A2(n758), .B1(n131), .B2(n7318), .ZN(n3616) );
  OAI22_X1 U836 ( .A1(n243), .A2(n759), .B1(n131), .B2(n7370), .ZN(n3617) );
  OAI22_X1 U838 ( .A1(n246), .A2(n760), .B1(n131), .B2(n248), .ZN(n3618) );
  OAI22_X1 U839 ( .A1(n249), .A2(n761), .B1(n131), .B2(n251), .ZN(n3619) );
  OAI22_X1 U840 ( .A1(n252), .A2(n762), .B1(n131), .B2(n7271), .ZN(n3620) );
  OAI22_X1 U841 ( .A1(n255), .A2(n763), .B1(n131), .B2(n257), .ZN(n3621) );
  OAI22_X1 U843 ( .A1(n258), .A2(n764), .B1(n131), .B2(n7117), .ZN(n3622) );
  OAI22_X1 U844 ( .A1(n7115), .A2(n5243), .B1(n131), .B2(n262), .ZN(n3623) );
  OAI22_X1 U845 ( .A1(n263), .A2(n5211), .B1(n131), .B2(n7158), .ZN(n3624) );
  OAI22_X1 U846 ( .A1(n6896), .A2(n765), .B1(n131), .B2(n6898), .ZN(n3625) );
  OAI22_X1 U847 ( .A1(n268), .A2(n5147), .B1(n131), .B2(n269), .ZN(n3626) );
  OAI22_X1 U848 ( .A1(n270), .A2(n5115), .B1(n131), .B2(n271), .ZN(n3627) );
  OAI22_X1 U849 ( .A1(n272), .A2(n766), .B1(n131), .B2(n274), .ZN(n3628) );
  OAI22_X1 U850 ( .A1(n275), .A2(n767), .B1(n131), .B2(n7363), .ZN(n3629) );
  OAI22_X1 U851 ( .A1(n278), .A2(n5019), .B1(n131), .B2(n7276), .ZN(n3630) );
  OAI22_X1 U852 ( .A1(n7122), .A2(n4987), .B1(n131), .B2(n281), .ZN(n3631) );
  OAI22_X1 U853 ( .A1(n282), .A2(n768), .B1(n131), .B2(n284), .ZN(n3632) );
  OAI22_X1 U854 ( .A1(n7119), .A2(n769), .B1(n131), .B2(n287), .ZN(n3633) );
  OAI22_X1 U855 ( .A1(n288), .A2(n4891), .B1(n131), .B2(n289), .ZN(n3634) );
  OAI22_X1 U856 ( .A1(n290), .A2(n4859), .B1(n131), .B2(n291), .ZN(n3635) );
  OAI22_X1 U857 ( .A1(n292), .A2(n770), .B1(n131), .B2(n294), .ZN(n3636) );
  OAI22_X1 U859 ( .A1(n295), .A2(n771), .B1(n131), .B2(n297), .ZN(n3637) );
  OAI22_X1 U861 ( .A1(n298), .A2(n772), .B1(n131), .B2(n300), .ZN(n3638) );
  OAI22_X1 U862 ( .A1(n6559), .A2(n773), .B1(n131), .B2(n7076), .ZN(n3639) );
  OAI22_X1 U864 ( .A1(n304), .A2(n4699), .B1(n131), .B2(n7113), .ZN(n3640) );
  OAI22_X1 U865 ( .A1(n7112), .A2(n4667), .B1(n131), .B2(n307), .ZN(n3641) );
  OAI22_X1 U866 ( .A1(n308), .A2(n774), .B1(n131), .B2(n310), .ZN(n3642) );
  OAI22_X1 U867 ( .A1(n7074), .A2(n775), .B1(n131), .B2(n313), .ZN(n3643) );
  OAI22_X1 U868 ( .A1(n314), .A2(n776), .B1(n131), .B2(n7210), .ZN(n3644) );
  OAI22_X1 U869 ( .A1(n317), .A2(n777), .B1(n131), .B2(n7209), .ZN(n3645) );
  OAI211_X1 U871 ( .C1(n5821), .C2(n653), .A(n654), .B(n778), .ZN(n754) );
  AOI22_X1 U872 ( .A1(n656), .A2(n6535), .B1(n779), .B2(n658), .ZN(n778) );
  INV_X1 U873 ( .A(n5611), .ZN(n779) );
  OAI22_X1 U874 ( .A1(n5611), .A2(net55846), .B1(n130), .B2(net55908), .ZN(
        n3646) );
  INV_X1 U875 ( .A(n753), .ZN(n130) );
  OAI222_X1 U876 ( .A1(n780), .A2(n323), .B1(n6365), .B2(n402), .C1(n781), 
        .C2(n322), .ZN(n753) );
  INV_X1 U877 ( .A(n6369), .ZN(n781) );
  INV_X1 U878 ( .A(n6368), .ZN(n780) );
  OAI221_X1 U879 ( .B1(n357), .B2(n782), .C1(n359), .C2(n783), .A(n784), .ZN(
        n3647) );
  AOI22_X1 U880 ( .A1(\Mcontrol/bvgen/d_curr_pc[13] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [13]), .B2(n362), .ZN(n784) );
  OAI222_X1 U882 ( .A1(n364), .A2(n785), .B1(n366), .B2(n786), .C1(net55850), 
        .C2(n782), .ZN(n3648) );
  OAI22_X1 U884 ( .A1(net55878), .A2(n786), .B1(net55834), .B2(n785), .ZN(
        n3649) );
  INV_X1 U887 ( .A(n787), .ZN(n3650) );
  AOI22_X1 U888 ( .A1(n7189), .A2(\Mcontrol/f_currpc[13] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[13] ), .ZN(n787) );
  INV_X1 U889 ( .A(n788), .ZN(n3651) );
  AOI221_X1 U890 ( .B1(n371), .B2(\Mcontrol/f_currpc[13] ), .C1(n372), .C2(
        n7878), .A(n373), .ZN(n788) );
  OAI221_X1 U891 ( .B1(n789), .B2(n214), .C1(\Mpath/the_alu/N58 ), .C2(
        net55854), .A(n790), .ZN(n3652) );
  AOI222_X1 U892 ( .A1(n197), .A2(n129), .B1(n192), .B2(n791), .C1(n195), .C2(
        n792), .ZN(n790) );
  INV_X1 U893 ( .A(break_code[13]), .ZN(n789) );
  OAI221_X1 U894 ( .B1(n127), .B2(n232), .C1(\Mpath/the_alu/N57 ), .C2(
        net55854), .A(n793), .ZN(n3653) );
  AOI22_X1 U895 ( .A1(n6556), .A2(n791), .B1(n6560), .B2(n794), .ZN(n793) );
  OAI22_X1 U896 ( .A1(n237), .A2(n795), .B1(n127), .B2(n239), .ZN(n3654) );
  OAI22_X1 U897 ( .A1(n240), .A2(n796), .B1(n127), .B2(n7318), .ZN(n3655) );
  OAI22_X1 U898 ( .A1(n243), .A2(n797), .B1(n127), .B2(n7370), .ZN(n3656) );
  OAI22_X1 U900 ( .A1(n246), .A2(n798), .B1(n127), .B2(n248), .ZN(n3657) );
  OAI22_X1 U901 ( .A1(n249), .A2(n799), .B1(n127), .B2(n251), .ZN(n3658) );
  OAI22_X1 U902 ( .A1(n252), .A2(n800), .B1(n127), .B2(n7271), .ZN(n3659) );
  OAI22_X1 U903 ( .A1(n255), .A2(n801), .B1(n127), .B2(n257), .ZN(n3660) );
  OAI22_X1 U905 ( .A1(n258), .A2(n802), .B1(n127), .B2(n7117), .ZN(n3661) );
  OAI22_X1 U906 ( .A1(n7115), .A2(n5242), .B1(n127), .B2(n262), .ZN(n3662) );
  OAI22_X1 U907 ( .A1(n263), .A2(n5210), .B1(n127), .B2(n7158), .ZN(n3663) );
  OAI22_X1 U908 ( .A1(n6895), .A2(n803), .B1(n127), .B2(n6898), .ZN(n3664) );
  OAI22_X1 U909 ( .A1(n268), .A2(n5146), .B1(n127), .B2(n269), .ZN(n3665) );
  OAI22_X1 U910 ( .A1(n270), .A2(n5114), .B1(n127), .B2(n271), .ZN(n3666) );
  OAI22_X1 U911 ( .A1(n272), .A2(n804), .B1(n127), .B2(n274), .ZN(n3667) );
  OAI22_X1 U912 ( .A1(n275), .A2(n805), .B1(n127), .B2(n7363), .ZN(n3668) );
  OAI22_X1 U913 ( .A1(n278), .A2(n5018), .B1(n127), .B2(n7276), .ZN(n3669) );
  OAI22_X1 U914 ( .A1(n7122), .A2(n4986), .B1(n127), .B2(n281), .ZN(n3670) );
  OAI22_X1 U915 ( .A1(n282), .A2(n806), .B1(n127), .B2(n284), .ZN(n3671) );
  OAI22_X1 U916 ( .A1(n7119), .A2(n807), .B1(n127), .B2(n287), .ZN(n3672) );
  OAI22_X1 U917 ( .A1(n288), .A2(n4890), .B1(n127), .B2(n289), .ZN(n3673) );
  OAI22_X1 U918 ( .A1(n290), .A2(n4858), .B1(n127), .B2(n291), .ZN(n3674) );
  OAI22_X1 U919 ( .A1(n292), .A2(n808), .B1(n127), .B2(n294), .ZN(n3675) );
  OAI22_X1 U921 ( .A1(n295), .A2(n809), .B1(n127), .B2(n297), .ZN(n3676) );
  OAI22_X1 U923 ( .A1(n298), .A2(n810), .B1(n127), .B2(n300), .ZN(n3677) );
  OAI22_X1 U924 ( .A1(n6559), .A2(n811), .B1(n127), .B2(n7076), .ZN(n3678) );
  OAI22_X1 U926 ( .A1(n304), .A2(n4698), .B1(n127), .B2(n7113), .ZN(n3679) );
  OAI22_X1 U927 ( .A1(n7112), .A2(n4666), .B1(n127), .B2(n307), .ZN(n3680) );
  OAI22_X1 U928 ( .A1(n308), .A2(n812), .B1(n127), .B2(n310), .ZN(n3681) );
  OAI22_X1 U929 ( .A1(n7074), .A2(n813), .B1(n127), .B2(n313), .ZN(n3682) );
  OAI22_X1 U930 ( .A1(n314), .A2(n814), .B1(n127), .B2(n7210), .ZN(n3683) );
  OAI22_X1 U931 ( .A1(n317), .A2(n815), .B1(n127), .B2(n7209), .ZN(n3684) );
  OAI211_X1 U933 ( .C1(n5811), .C2(n653), .A(n654), .B(n816), .ZN(n792) );
  AOI22_X1 U934 ( .A1(n656), .A2(n6537), .B1(n817), .B2(n658), .ZN(n816) );
  INV_X1 U935 ( .A(n5608), .ZN(n817) );
  OAI22_X1 U936 ( .A1(n5608), .A2(net55846), .B1(n126), .B2(net55906), .ZN(
        n3685) );
  INV_X1 U937 ( .A(n791), .ZN(n126) );
  OAI222_X1 U938 ( .A1(n818), .A2(n323), .B1(n6353), .B2(n402), .C1(n819), 
        .C2(n322), .ZN(n791) );
  INV_X1 U939 ( .A(n6357), .ZN(n819) );
  INV_X1 U940 ( .A(n6356), .ZN(n818) );
  OAI221_X1 U941 ( .B1(n357), .B2(n820), .C1(n359), .C2(n821), .A(n822), .ZN(
        n3686) );
  AOI22_X1 U942 ( .A1(\Mcontrol/bvgen/d_curr_pc[8] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [8]), .B2(n362), .ZN(n822) );
  OAI222_X1 U944 ( .A1(n364), .A2(n823), .B1(n366), .B2(n824), .C1(net55850), 
        .C2(n820), .ZN(n3687) );
  OAI22_X1 U946 ( .A1(net55876), .A2(n824), .B1(net55834), .B2(n823), .ZN(
        n3688) );
  INV_X1 U949 ( .A(n825), .ZN(n3689) );
  AOI22_X1 U950 ( .A1(n7189), .A2(\Mcontrol/f_currpc[8] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[8] ), .ZN(n825) );
  INV_X1 U951 ( .A(n826), .ZN(n3690) );
  OAI221_X1 U953 ( .B1(n827), .B2(n214), .C1(\Mpath/the_alu/N68 ), .C2(
        net55854), .A(n828), .ZN(n3691) );
  AOI222_X1 U954 ( .A1(n197), .A2(n149), .B1(n192), .B2(n829), .C1(n195), .C2(
        n830), .ZN(n828) );
  INV_X1 U955 ( .A(break_code[8]), .ZN(n827) );
  OAI221_X1 U956 ( .B1(n357), .B2(n831), .C1(n359), .C2(n832), .A(n833), .ZN(
        n3692) );
  AOI22_X1 U957 ( .A1(\Mcontrol/bvgen/d_curr_pc[4] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [4]), .B2(n362), .ZN(n833) );
  OAI222_X1 U959 ( .A1(n364), .A2(n834), .B1(n366), .B2(n835), .C1(net55850), 
        .C2(n831), .ZN(n3693) );
  OAI22_X1 U961 ( .A1(net55876), .A2(n835), .B1(net55828), .B2(n834), .ZN(
        n3694) );
  INV_X1 U964 ( .A(n836), .ZN(n3695) );
  AOI22_X1 U965 ( .A1(n7189), .A2(\Mcontrol/f_currpc[4] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[4] ), .ZN(n836) );
  INV_X1 U966 ( .A(n837), .ZN(n3696) );
  OAI221_X1 U968 ( .B1(n838), .B2(n214), .C1(\Mpath/the_alu/N76 ), .C2(
        net55854), .A(n839), .ZN(n3697) );
  AOI222_X1 U969 ( .A1(n197), .A2(n165), .B1(n192), .B2(n840), .C1(n195), .C2(
        n841), .ZN(n839) );
  INV_X1 U970 ( .A(break_code[4]), .ZN(n838) );
  OAI221_X1 U971 ( .B1(n357), .B2(n842), .C1(n359), .C2(n843), .A(n844), .ZN(
        n3698) );
  AOI22_X1 U972 ( .A1(\Mcontrol/bvgen/d_curr_pc[3] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [3]), .B2(n362), .ZN(n844) );
  OAI222_X1 U974 ( .A1(n364), .A2(n845), .B1(n366), .B2(n846), .C1(net55850), 
        .C2(n842), .ZN(n3699) );
  OAI22_X1 U976 ( .A1(net55876), .A2(n846), .B1(net55826), .B2(n845), .ZN(
        n3700) );
  INV_X1 U979 ( .A(n847), .ZN(n3701) );
  AOI22_X1 U980 ( .A1(n7189), .A2(\Mcontrol/f_currpc[3] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[3] ), .ZN(n847) );
  INV_X1 U981 ( .A(n848), .ZN(n3702) );
  OAI221_X1 U983 ( .B1(n849), .B2(n214), .C1(\Mpath/the_alu/N78 ), .C2(
        net55854), .A(n850), .ZN(n3703) );
  AOI222_X1 U984 ( .A1(n197), .A2(n169), .B1(n192), .B2(n851), .C1(n195), .C2(
        n852), .ZN(n850) );
  INV_X1 U985 ( .A(n7311), .ZN(n849) );
  OAI221_X1 U986 ( .B1(n357), .B2(n853), .C1(n359), .C2(n854), .A(n855), .ZN(
        n3704) );
  AOI22_X1 U987 ( .A1(\Mcontrol/bvgen/d_curr_pc[2] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [2]), .B2(n362), .ZN(n855) );
  OAI222_X1 U989 ( .A1(n364), .A2(n856), .B1(n366), .B2(n857), .C1(net55848), 
        .C2(n853), .ZN(n3705) );
  OAI22_X1 U991 ( .A1(net55876), .A2(n857), .B1(net55830), .B2(n856), .ZN(
        n3706) );
  INV_X1 U994 ( .A(n858), .ZN(n3707) );
  AOI22_X1 U995 ( .A1(n7189), .A2(\Mcontrol/f_currpc[2] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[2] ), .ZN(n858) );
  INV_X1 U996 ( .A(n859), .ZN(n3708) );
  OAI221_X1 U998 ( .B1(n860), .B2(n214), .C1(\Mpath/the_alu/N80 ), .C2(
        net55854), .A(n861), .ZN(n3709) );
  AOI222_X1 U999 ( .A1(n197), .A2(n173), .B1(n192), .B2(n862), .C1(n195), .C2(
        n863), .ZN(n861) );
  INV_X1 U1000 ( .A(n7353), .ZN(n860) );
  OAI221_X1 U1001 ( .B1(n357), .B2(n864), .C1(n359), .C2(n865), .A(n866), .ZN(
        n3710) );
  AOI22_X1 U1002 ( .A1(\Mcontrol/bvgen/d_curr_pc[1] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [1]), .B2(n362), .ZN(n866) );
  OAI222_X1 U1004 ( .A1(n364), .A2(n867), .B1(n366), .B2(n868), .C1(net55850), 
        .C2(n864), .ZN(n3711) );
  OAI22_X1 U1006 ( .A1(net55876), .A2(n868), .B1(net55828), .B2(n867), .ZN(
        n3712) );
  OAI22_X1 U1008 ( .A1(n7030), .A2(n869), .B1(n7189), .B2(n868), .ZN(n3713) );
  OAI21_X1 U1010 ( .B1(n372), .B2(n869), .A(n870), .ZN(n3714) );
  NAND3_X1 U1011 ( .A1(n7083), .A2(n6547), .A3(n372), .ZN(n870) );
  OAI221_X1 U1013 ( .B1(n357), .B2(n872), .C1(n359), .C2(n873), .A(n874), .ZN(
        n3715) );
  AOI22_X1 U1014 ( .A1(\Mcontrol/bvgen/d_curr_pc[5] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [5]), .B2(n362), .ZN(n874) );
  OAI222_X1 U1016 ( .A1(n364), .A2(n875), .B1(n366), .B2(n876), .C1(net55848), 
        .C2(n872), .ZN(n3716) );
  OAI22_X1 U1018 ( .A1(net55876), .A2(n876), .B1(net55830), .B2(n875), .ZN(
        n3717) );
  INV_X1 U1021 ( .A(n877), .ZN(n3718) );
  AOI22_X1 U1022 ( .A1(n7189), .A2(\Mcontrol/f_currpc[5] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[5] ), .ZN(n877) );
  INV_X1 U1023 ( .A(n878), .ZN(n3719) );
  OAI221_X1 U1025 ( .B1(n879), .B2(n214), .C1(\Mpath/the_alu/N74 ), .C2(
        net55854), .A(n880), .ZN(n3720) );
  AOI222_X1 U1026 ( .A1(n197), .A2(n161), .B1(n192), .B2(n881), .C1(n195), 
        .C2(n882), .ZN(n880) );
  INV_X1 U1027 ( .A(break_code[5]), .ZN(n879) );
  OAI22_X1 U1028 ( .A1(n6487), .A2(n7110), .B1(serve_exception), .B2(n48), 
        .ZN(n3721) );
  AOI22_X1 U1029 ( .A1(\Scc_coproc/x_exc_word[1] ), .A2(n883), .B1(n884), .B2(
        n885), .ZN(n48) );
  INV_X1 U1030 ( .A(n886), .ZN(n884) );
  AOI211_X1 U1031 ( .C1(n5741), .C2(n5742), .A(\Scc_coproc/interrupt[7] ), .B(
        \Scc_coproc/interrupt[6] ), .ZN(n886) );
  OAI22_X1 U1032 ( .A1(n5729), .A2(net55916), .B1(net55830), .B2(n887), .ZN(
        n3722) );
  OAI22_X1 U1033 ( .A1(n5730), .A2(n626), .B1(n5729), .B2(n627), .ZN(n3723) );
  OAI222_X1 U1034 ( .A1(n628), .A2(n887), .B1(n5729), .B2(n629), .C1(n5730), 
        .C2(n359), .ZN(n3724) );
  OAI221_X1 U1036 ( .B1(n159), .B2(n232), .C1(\Mpath/the_alu/N73 ), .C2(
        net55854), .A(n888), .ZN(n3725) );
  AOI22_X1 U1037 ( .A1(n6556), .A2(n881), .B1(n6560), .B2(n889), .ZN(n888) );
  OAI22_X1 U1038 ( .A1(n237), .A2(n890), .B1(n159), .B2(n239), .ZN(n3726) );
  OAI22_X1 U1039 ( .A1(n240), .A2(n891), .B1(n159), .B2(n7318), .ZN(n3727) );
  OAI22_X1 U1040 ( .A1(n243), .A2(n892), .B1(n159), .B2(n7370), .ZN(n3728) );
  OAI22_X1 U1042 ( .A1(n246), .A2(n893), .B1(n159), .B2(n248), .ZN(n3729) );
  OAI22_X1 U1043 ( .A1(n249), .A2(n894), .B1(n159), .B2(n251), .ZN(n3730) );
  OAI22_X1 U1044 ( .A1(n252), .A2(n895), .B1(n159), .B2(n7271), .ZN(n3731) );
  OAI22_X1 U1045 ( .A1(n255), .A2(n896), .B1(n159), .B2(n257), .ZN(n3732) );
  OAI22_X1 U1047 ( .A1(n258), .A2(n897), .B1(n159), .B2(n7117), .ZN(n3733) );
  OAI22_X1 U1048 ( .A1(n7115), .A2(n5219), .B1(n159), .B2(n262), .ZN(n3734) );
  OAI22_X1 U1049 ( .A1(n263), .A2(n5187), .B1(n159), .B2(n7158), .ZN(n3735) );
  OAI22_X1 U1050 ( .A1(n6895), .A2(n898), .B1(n159), .B2(n6898), .ZN(n3736) );
  OAI22_X1 U1051 ( .A1(n268), .A2(n5123), .B1(n159), .B2(n269), .ZN(n3737) );
  OAI22_X1 U1052 ( .A1(n270), .A2(n5091), .B1(n159), .B2(n271), .ZN(n3738) );
  OAI22_X1 U1053 ( .A1(n272), .A2(n899), .B1(n159), .B2(n274), .ZN(n3739) );
  OAI22_X1 U1054 ( .A1(n275), .A2(n900), .B1(n159), .B2(n7363), .ZN(n3740) );
  OAI22_X1 U1055 ( .A1(n278), .A2(n4995), .B1(n159), .B2(n7276), .ZN(n3741) );
  OAI22_X1 U1056 ( .A1(n7122), .A2(n4963), .B1(n159), .B2(n281), .ZN(n3742) );
  OAI22_X1 U1057 ( .A1(n282), .A2(n901), .B1(n159), .B2(n284), .ZN(n3743) );
  OAI22_X1 U1058 ( .A1(n7119), .A2(n902), .B1(n159), .B2(n287), .ZN(n3744) );
  OAI22_X1 U1059 ( .A1(n288), .A2(n4867), .B1(n159), .B2(n289), .ZN(n3745) );
  OAI22_X1 U1060 ( .A1(n290), .A2(n4835), .B1(n159), .B2(n291), .ZN(n3746) );
  OAI22_X1 U1061 ( .A1(n292), .A2(n903), .B1(n159), .B2(n294), .ZN(n3747) );
  OAI22_X1 U1063 ( .A1(n295), .A2(n904), .B1(n159), .B2(n297), .ZN(n3748) );
  OAI22_X1 U1065 ( .A1(n298), .A2(n905), .B1(n159), .B2(n300), .ZN(n3749) );
  OAI22_X1 U1066 ( .A1(n6559), .A2(n906), .B1(n159), .B2(n7076), .ZN(n3750) );
  OAI22_X1 U1068 ( .A1(n304), .A2(n4675), .B1(n159), .B2(n7113), .ZN(n3751) );
  OAI22_X1 U1069 ( .A1(n7112), .A2(n4643), .B1(n159), .B2(n307), .ZN(n3752) );
  OAI22_X1 U1070 ( .A1(n308), .A2(n907), .B1(n159), .B2(n310), .ZN(n3753) );
  OAI22_X1 U1071 ( .A1(n7074), .A2(n908), .B1(n159), .B2(n313), .ZN(n3754) );
  OAI22_X1 U1072 ( .A1(n314), .A2(n909), .B1(n159), .B2(n7210), .ZN(n3755) );
  OAI22_X1 U1073 ( .A1(n317), .A2(n910), .B1(n159), .B2(n7209), .ZN(n3756) );
  OAI211_X1 U1075 ( .C1(n5745), .C2(n5539), .A(n911), .B(n912), .ZN(n882) );
  AOI222_X1 U1076 ( .A1(n913), .A2(n6537), .B1(n6516), .B2(n914), .C1(n915), 
        .C2(n6524), .ZN(n912) );
  AOI22_X1 U1077 ( .A1(n5813), .A2(n916), .B1(n5810), .B2(n917), .ZN(n911) );
  OAI22_X1 U1078 ( .A1(n5539), .A2(net55846), .B1(n158), .B2(net55906), .ZN(
        n3757) );
  INV_X1 U1079 ( .A(n881), .ZN(n158) );
  OAI222_X1 U1080 ( .A1(n918), .A2(n323), .B1(n6163), .B2(n402), .C1(n919), 
        .C2(n322), .ZN(n881) );
  INV_X1 U1081 ( .A(n6167), .ZN(n919) );
  INV_X1 U1082 ( .A(n6166), .ZN(n918) );
  OAI221_X1 U1083 ( .B1(n357), .B2(n920), .C1(n359), .C2(n921), .A(n922), .ZN(
        n3758) );
  AOI22_X1 U1084 ( .A1(\Mcontrol/bvgen/d_curr_pc[6] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [6]), .B2(n362), .ZN(n922) );
  OAI222_X1 U1086 ( .A1(n364), .A2(n923), .B1(n366), .B2(n924), .C1(net55848), 
        .C2(n920), .ZN(n3759) );
  OAI22_X1 U1088 ( .A1(net55876), .A2(n924), .B1(net55828), .B2(n923), .ZN(
        n3760) );
  INV_X1 U1091 ( .A(n925), .ZN(n3761) );
  AOI22_X1 U1092 ( .A1(n7189), .A2(\Mcontrol/f_currpc[6] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[6] ), .ZN(n925) );
  INV_X1 U1093 ( .A(n926), .ZN(n3762) );
  AOI221_X1 U1094 ( .B1(n371), .B2(\Mcontrol/f_currpc[6] ), .C1(n372), .C2(
        n7884), .A(n373), .ZN(n926) );
  OAI221_X1 U1095 ( .B1(n927), .B2(n214), .C1(\Mpath/the_alu/N72 ), .C2(
        net55856), .A(n928), .ZN(n3763) );
  AOI222_X1 U1096 ( .A1(n197), .A2(n157), .B1(n192), .B2(n929), .C1(n195), 
        .C2(n930), .ZN(n928) );
  INV_X1 U1097 ( .A(break_code[6]), .ZN(n927) );
  OAI22_X1 U1098 ( .A1(n5727), .A2(net55912), .B1(net55830), .B2(n931), .ZN(
        n3764) );
  OAI22_X1 U1099 ( .A1(n5728), .A2(n626), .B1(n5727), .B2(n627), .ZN(n3765) );
  OAI222_X1 U1100 ( .A1(n628), .A2(n931), .B1(n5727), .B2(n629), .C1(n5728), 
        .C2(n359), .ZN(n3766) );
  OAI221_X1 U1102 ( .B1(n155), .B2(n232), .C1(\Mpath/the_alu/N71 ), .C2(
        net55856), .A(n932), .ZN(n3767) );
  AOI22_X1 U1103 ( .A1(n6556), .A2(n929), .B1(n6560), .B2(n933), .ZN(n932) );
  OAI22_X1 U1104 ( .A1(n237), .A2(n934), .B1(n155), .B2(n239), .ZN(n3768) );
  OAI22_X1 U1105 ( .A1(n240), .A2(n935), .B1(n155), .B2(n7318), .ZN(n3769) );
  OAI22_X1 U1106 ( .A1(n243), .A2(n936), .B1(n155), .B2(n7370), .ZN(n3770) );
  OAI22_X1 U1108 ( .A1(n246), .A2(n937), .B1(n155), .B2(n248), .ZN(n3771) );
  OAI22_X1 U1109 ( .A1(n249), .A2(n938), .B1(n155), .B2(n251), .ZN(n3772) );
  OAI22_X1 U1110 ( .A1(n252), .A2(n939), .B1(n155), .B2(n7271), .ZN(n3773) );
  OAI22_X1 U1111 ( .A1(n255), .A2(n940), .B1(n155), .B2(n257), .ZN(n3774) );
  OAI22_X1 U1113 ( .A1(n258), .A2(n941), .B1(n155), .B2(n7117), .ZN(n3775) );
  OAI22_X1 U1114 ( .A1(n7115), .A2(n5218), .B1(n155), .B2(n262), .ZN(n3776) );
  OAI22_X1 U1115 ( .A1(n263), .A2(n5186), .B1(n155), .B2(n7158), .ZN(n3777) );
  OAI22_X1 U1116 ( .A1(n6897), .A2(n942), .B1(n155), .B2(n6898), .ZN(n3778) );
  OAI22_X1 U1117 ( .A1(n268), .A2(n5122), .B1(n155), .B2(n269), .ZN(n3779) );
  OAI22_X1 U1118 ( .A1(n270), .A2(n5090), .B1(n155), .B2(n271), .ZN(n3780) );
  OAI22_X1 U1119 ( .A1(n272), .A2(n943), .B1(n155), .B2(n274), .ZN(n3781) );
  OAI22_X1 U1120 ( .A1(n275), .A2(n944), .B1(n155), .B2(n7363), .ZN(n3782) );
  OAI22_X1 U1121 ( .A1(n278), .A2(n4994), .B1(n155), .B2(n7276), .ZN(n3783) );
  OAI22_X1 U1122 ( .A1(n7122), .A2(n4962), .B1(n155), .B2(n281), .ZN(n3784) );
  OAI22_X1 U1123 ( .A1(n282), .A2(n945), .B1(n155), .B2(n284), .ZN(n3785) );
  OAI22_X1 U1124 ( .A1(n7119), .A2(n946), .B1(n155), .B2(n287), .ZN(n3786) );
  OAI22_X1 U1125 ( .A1(n288), .A2(n4866), .B1(n155), .B2(n289), .ZN(n3787) );
  OAI22_X1 U1126 ( .A1(n290), .A2(n4834), .B1(n155), .B2(n291), .ZN(n3788) );
  OAI22_X1 U1127 ( .A1(n292), .A2(n947), .B1(n155), .B2(n294), .ZN(n3789) );
  OAI22_X1 U1129 ( .A1(n295), .A2(n948), .B1(n155), .B2(n297), .ZN(n3790) );
  OAI22_X1 U1131 ( .A1(n298), .A2(n949), .B1(n155), .B2(n300), .ZN(n3791) );
  OAI22_X1 U1132 ( .A1(n6558), .A2(n950), .B1(n155), .B2(n7076), .ZN(n3792) );
  OAI22_X1 U1134 ( .A1(n304), .A2(n4674), .B1(n155), .B2(n7113), .ZN(n3793) );
  OAI22_X1 U1135 ( .A1(n7112), .A2(n4642), .B1(n155), .B2(n307), .ZN(n3794) );
  OAI22_X1 U1136 ( .A1(n308), .A2(n951), .B1(n155), .B2(n310), .ZN(n3795) );
  OAI22_X1 U1137 ( .A1(n7074), .A2(n952), .B1(n155), .B2(n313), .ZN(n3796) );
  OAI22_X1 U1138 ( .A1(n314), .A2(n953), .B1(n155), .B2(n7210), .ZN(n3797) );
  OAI22_X1 U1139 ( .A1(n317), .A2(n954), .B1(n155), .B2(n7209), .ZN(n3798) );
  OAI211_X1 U1141 ( .C1(n5745), .C2(n5536), .A(n955), .B(n956), .ZN(n930) );
  AOI222_X1 U1142 ( .A1(n913), .A2(n6539), .B1(n6514), .B2(n914), .C1(n915), 
        .C2(n6525), .ZN(n956) );
  AOI22_X1 U1143 ( .A1(n5801), .A2(n916), .B1(n5798), .B2(n917), .ZN(n955) );
  OAI22_X1 U1144 ( .A1(n5536), .A2(net55844), .B1(n154), .B2(net55902), .ZN(
        n3799) );
  INV_X1 U1145 ( .A(n929), .ZN(n154) );
  OAI222_X1 U1146 ( .A1(n957), .A2(n323), .B1(n6151), .B2(n402), .C1(n958), 
        .C2(n322), .ZN(n929) );
  INV_X1 U1147 ( .A(n6155), .ZN(n958) );
  INV_X1 U1148 ( .A(n6154), .ZN(n957) );
  OAI221_X1 U1149 ( .B1(n357), .B2(n959), .C1(n359), .C2(n960), .A(n961), .ZN(
        n3800) );
  AOI22_X1 U1150 ( .A1(\Mcontrol/bvgen/d_curr_pc[7] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [7]), .B2(n362), .ZN(n961) );
  OAI222_X1 U1152 ( .A1(n364), .A2(n962), .B1(n366), .B2(n963), .C1(net55848), 
        .C2(n959), .ZN(n3801) );
  OAI22_X1 U1154 ( .A1(net55874), .A2(n963), .B1(net55830), .B2(n962), .ZN(
        n3802) );
  INV_X1 U1157 ( .A(n964), .ZN(n3803) );
  AOI22_X1 U1158 ( .A1(n7189), .A2(\Mcontrol/f_currpc[7] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[7] ), .ZN(n964) );
  INV_X1 U1159 ( .A(n965), .ZN(n3804) );
  AOI221_X1 U1160 ( .B1(n371), .B2(\Mcontrol/f_currpc[7] ), .C1(n372), .C2(
        n7883), .A(n373), .ZN(n965) );
  OAI221_X1 U1161 ( .B1(n966), .B2(n214), .C1(\Mpath/the_alu/N70 ), .C2(
        net55856), .A(n967), .ZN(n3805) );
  AOI222_X1 U1162 ( .A1(n197), .A2(n153), .B1(n192), .B2(n968), .C1(n195), 
        .C2(n969), .ZN(n967) );
  INV_X1 U1163 ( .A(break_code[7]), .ZN(n966) );
  OAI22_X1 U1164 ( .A1(n5725), .A2(net55916), .B1(net55828), .B2(n970), .ZN(
        n3806) );
  OAI22_X1 U1165 ( .A1(n5726), .A2(n626), .B1(n5725), .B2(n627), .ZN(n3807) );
  OAI222_X1 U1166 ( .A1(n628), .A2(n970), .B1(n5725), .B2(n629), .C1(n5726), 
        .C2(n359), .ZN(n3808) );
  OAI221_X1 U1168 ( .B1(n151), .B2(n232), .C1(\Mpath/the_alu/N69 ), .C2(
        net55852), .A(n971), .ZN(n3809) );
  AOI22_X1 U1169 ( .A1(n6556), .A2(n968), .B1(n6560), .B2(n972), .ZN(n971) );
  OAI22_X1 U1170 ( .A1(n237), .A2(n973), .B1(n151), .B2(n239), .ZN(n3810) );
  OAI22_X1 U1171 ( .A1(n240), .A2(n974), .B1(n151), .B2(n7318), .ZN(n3811) );
  OAI22_X1 U1172 ( .A1(n243), .A2(n975), .B1(n151), .B2(n7370), .ZN(n3812) );
  OAI22_X1 U1174 ( .A1(n246), .A2(n976), .B1(n151), .B2(n248), .ZN(n3813) );
  OAI22_X1 U1175 ( .A1(n249), .A2(n977), .B1(n151), .B2(n251), .ZN(n3814) );
  OAI22_X1 U1176 ( .A1(n252), .A2(n978), .B1(n151), .B2(n7271), .ZN(n3815) );
  OAI22_X1 U1177 ( .A1(n255), .A2(n979), .B1(n151), .B2(n257), .ZN(n3816) );
  OAI22_X1 U1179 ( .A1(n258), .A2(n980), .B1(n151), .B2(n7117), .ZN(n3817) );
  OAI22_X1 U1180 ( .A1(n7115), .A2(n5217), .B1(n151), .B2(n262), .ZN(n3818) );
  OAI22_X1 U1181 ( .A1(n263), .A2(n5185), .B1(n151), .B2(n7158), .ZN(n3819) );
  OAI22_X1 U1182 ( .A1(n6896), .A2(n981), .B1(n151), .B2(n6898), .ZN(n3820) );
  OAI22_X1 U1183 ( .A1(n268), .A2(n5121), .B1(n151), .B2(n269), .ZN(n3821) );
  OAI22_X1 U1184 ( .A1(n270), .A2(n5089), .B1(n151), .B2(n271), .ZN(n3822) );
  OAI22_X1 U1185 ( .A1(n272), .A2(n982), .B1(n151), .B2(n274), .ZN(n3823) );
  OAI22_X1 U1186 ( .A1(n275), .A2(n983), .B1(n151), .B2(n7363), .ZN(n3824) );
  OAI22_X1 U1187 ( .A1(n278), .A2(n4993), .B1(n151), .B2(n7276), .ZN(n3825) );
  OAI22_X1 U1188 ( .A1(n7122), .A2(n4961), .B1(n151), .B2(n281), .ZN(n3826) );
  OAI22_X1 U1189 ( .A1(n282), .A2(n984), .B1(n151), .B2(n284), .ZN(n3827) );
  OAI22_X1 U1190 ( .A1(n7119), .A2(n985), .B1(n151), .B2(n287), .ZN(n3828) );
  OAI22_X1 U1191 ( .A1(n288), .A2(n4865), .B1(n151), .B2(n289), .ZN(n3829) );
  OAI22_X1 U1192 ( .A1(n290), .A2(n4833), .B1(n151), .B2(n291), .ZN(n3830) );
  OAI22_X1 U1193 ( .A1(n292), .A2(n986), .B1(n151), .B2(n294), .ZN(n3831) );
  OAI22_X1 U1195 ( .A1(n295), .A2(n987), .B1(n151), .B2(n297), .ZN(n3832) );
  OAI22_X1 U1197 ( .A1(n298), .A2(n988), .B1(n151), .B2(n300), .ZN(n3833) );
  OAI22_X1 U1198 ( .A1(n6559), .A2(n989), .B1(n151), .B2(n7076), .ZN(n3834) );
  OAI22_X1 U1200 ( .A1(n304), .A2(n4673), .B1(n151), .B2(n7113), .ZN(n3835) );
  OAI22_X1 U1201 ( .A1(n7112), .A2(n4641), .B1(n151), .B2(n307), .ZN(n3836) );
  OAI22_X1 U1202 ( .A1(n308), .A2(n990), .B1(n151), .B2(n310), .ZN(n3837) );
  OAI22_X1 U1203 ( .A1(n7074), .A2(n991), .B1(n151), .B2(n313), .ZN(n3838) );
  OAI22_X1 U1204 ( .A1(n314), .A2(n992), .B1(n151), .B2(n7210), .ZN(n3839) );
  OAI22_X1 U1205 ( .A1(n317), .A2(n993), .B1(n151), .B2(n7209), .ZN(n3840) );
  OAI222_X1 U1207 ( .A1(n5785), .A2(n658), .B1(n994), .B2(n995), .C1(n5745), 
        .C2(n5533), .ZN(n969) );
  AOI221_X1 U1208 ( .B1(n5786), .B2(n6540), .C1(n5787), .C2(n6544), .A(n5788), 
        .ZN(n994) );
  OAI22_X1 U1209 ( .A1(n5533), .A2(net55846), .B1(n150), .B2(net55904), .ZN(
        n3841) );
  INV_X1 U1210 ( .A(n968), .ZN(n150) );
  OAI222_X1 U1211 ( .A1(n996), .A2(n323), .B1(n6139), .B2(n402), .C1(n997), 
        .C2(n322), .ZN(n968) );
  INV_X1 U1212 ( .A(n6143), .ZN(n997) );
  INV_X1 U1213 ( .A(n6142), .ZN(n996) );
  OAI221_X1 U1214 ( .B1(n357), .B2(n998), .C1(n359), .C2(n999), .A(n1000), 
        .ZN(n3842) );
  AOI22_X1 U1215 ( .A1(\Mcontrol/bvgen/d_curr_pc[9] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [9]), .B2(n362), .ZN(n1000) );
  OAI222_X1 U1217 ( .A1(n364), .A2(n1001), .B1(n366), .B2(n1002), .C1(net55848), .C2(n998), .ZN(n3843) );
  OAI22_X1 U1219 ( .A1(net55874), .A2(n1002), .B1(net55832), .B2(n1001), .ZN(
        n3844) );
  INV_X1 U1222 ( .A(n1003), .ZN(n3845) );
  AOI22_X1 U1223 ( .A1(n7189), .A2(\Mcontrol/f_currpc[9] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[9] ), .ZN(n1003) );
  INV_X1 U1224 ( .A(n1004), .ZN(n3846) );
  AOI221_X1 U1225 ( .B1(n371), .B2(\Mcontrol/f_currpc[9] ), .C1(n372), .C2(
        n7882), .A(n373), .ZN(n1004) );
  OAI221_X1 U1226 ( .B1(n1005), .B2(n214), .C1(\Mpath/the_alu/N66 ), .C2(
        net55852), .A(n1006), .ZN(n3847) );
  AOI222_X1 U1227 ( .A1(n197), .A2(n145), .B1(n192), .B2(n1007), .C1(n195), 
        .C2(n1008), .ZN(n1006) );
  INV_X1 U1228 ( .A(break_code[9]), .ZN(n1005) );
  OAI22_X1 U1229 ( .A1(n5721), .A2(net55912), .B1(net55828), .B2(n1009), .ZN(
        n3848) );
  OAI22_X1 U1230 ( .A1(n5722), .A2(n626), .B1(n5721), .B2(n627), .ZN(n3849) );
  OAI222_X1 U1231 ( .A1(n628), .A2(n1009), .B1(n5721), .B2(n629), .C1(n5722), 
        .C2(n359), .ZN(n3850) );
  OAI221_X1 U1233 ( .B1(n143), .B2(n232), .C1(\Mpath/the_alu/N65 ), .C2(
        net55852), .A(n1010), .ZN(n3851) );
  AOI22_X1 U1234 ( .A1(n6556), .A2(n1007), .B1(n6560), .B2(n1011), .ZN(n1010)
         );
  OAI22_X1 U1235 ( .A1(n237), .A2(n1012), .B1(n143), .B2(n239), .ZN(n3852) );
  OAI22_X1 U1236 ( .A1(n240), .A2(n1013), .B1(n143), .B2(n7318), .ZN(n3853) );
  OAI22_X1 U1237 ( .A1(n243), .A2(n1014), .B1(n143), .B2(n7370), .ZN(n3854) );
  OAI22_X1 U1239 ( .A1(n246), .A2(n1015), .B1(n143), .B2(n248), .ZN(n3855) );
  OAI22_X1 U1240 ( .A1(n249), .A2(n1016), .B1(n143), .B2(n251), .ZN(n3856) );
  OAI22_X1 U1241 ( .A1(n252), .A2(n1017), .B1(n143), .B2(n7271), .ZN(n3857) );
  OAI22_X1 U1242 ( .A1(n255), .A2(n1018), .B1(n143), .B2(n257), .ZN(n3858) );
  OAI22_X1 U1244 ( .A1(n258), .A2(n1019), .B1(n143), .B2(n7117), .ZN(n3859) );
  OAI22_X1 U1245 ( .A1(n7115), .A2(n5215), .B1(n143), .B2(n262), .ZN(n3860) );
  OAI22_X1 U1246 ( .A1(n263), .A2(n5183), .B1(n143), .B2(n7158), .ZN(n3861) );
  OAI22_X1 U1247 ( .A1(n6897), .A2(n1020), .B1(n143), .B2(n6898), .ZN(n3862)
         );
  OAI22_X1 U1248 ( .A1(n268), .A2(n5119), .B1(n143), .B2(n269), .ZN(n3863) );
  OAI22_X1 U1249 ( .A1(n270), .A2(n5087), .B1(n143), .B2(n271), .ZN(n3864) );
  OAI22_X1 U1250 ( .A1(n272), .A2(n1021), .B1(n143), .B2(n274), .ZN(n3865) );
  OAI22_X1 U1251 ( .A1(n275), .A2(n1022), .B1(n143), .B2(n7363), .ZN(n3866) );
  OAI22_X1 U1252 ( .A1(n278), .A2(n4991), .B1(n143), .B2(n7276), .ZN(n3867) );
  OAI22_X1 U1253 ( .A1(n7122), .A2(n4959), .B1(n143), .B2(n281), .ZN(n3868) );
  OAI22_X1 U1254 ( .A1(n282), .A2(n1023), .B1(n143), .B2(n284), .ZN(n3869) );
  OAI22_X1 U1255 ( .A1(n7119), .A2(n1024), .B1(n143), .B2(n287), .ZN(n3870) );
  OAI22_X1 U1256 ( .A1(n288), .A2(n4863), .B1(n143), .B2(n289), .ZN(n3871) );
  OAI22_X1 U1257 ( .A1(n290), .A2(n4831), .B1(n143), .B2(n291), .ZN(n3872) );
  OAI22_X1 U1258 ( .A1(n292), .A2(n1025), .B1(n143), .B2(n294), .ZN(n3873) );
  OAI22_X1 U1260 ( .A1(n295), .A2(n1026), .B1(n143), .B2(n297), .ZN(n3874) );
  OAI22_X1 U1262 ( .A1(n298), .A2(n1027), .B1(n143), .B2(n300), .ZN(n3875) );
  OAI22_X1 U1263 ( .A1(n6558), .A2(n1028), .B1(n143), .B2(n7076), .ZN(n3876)
         );
  OAI22_X1 U1265 ( .A1(n304), .A2(n4671), .B1(n143), .B2(n7113), .ZN(n3877) );
  OAI22_X1 U1266 ( .A1(n7112), .A2(n4639), .B1(n143), .B2(n307), .ZN(n3878) );
  OAI22_X1 U1267 ( .A1(n308), .A2(n1029), .B1(n143), .B2(n310), .ZN(n3879) );
  OAI22_X1 U1268 ( .A1(n7074), .A2(n1030), .B1(n143), .B2(n313), .ZN(n3880) );
  OAI22_X1 U1269 ( .A1(n314), .A2(n1031), .B1(n143), .B2(n7210), .ZN(n3881) );
  OAI22_X1 U1270 ( .A1(n317), .A2(n1032), .B1(n143), .B2(n7209), .ZN(n3882) );
  OAI211_X1 U1272 ( .C1(n5936), .C2(n653), .A(n654), .B(n1033), .ZN(n1008) );
  AOI22_X1 U1273 ( .A1(n656), .A2(n6529), .B1(n1034), .B2(n658), .ZN(n1033) );
  INV_X1 U1274 ( .A(n5526), .ZN(n1034) );
  OAI22_X1 U1275 ( .A1(n5526), .A2(net55842), .B1(n142), .B2(net55902), .ZN(
        n3883) );
  INV_X1 U1276 ( .A(n1007), .ZN(n142) );
  OAI222_X1 U1277 ( .A1(n1035), .A2(n323), .B1(n6114), .B2(n402), .C1(n1036), 
        .C2(n322), .ZN(n1007) );
  INV_X1 U1278 ( .A(n6118), .ZN(n1036) );
  INV_X1 U1279 ( .A(n6117), .ZN(n1035) );
  INV_X1 U1280 ( .A(n1037), .ZN(n3884) );
  AOI22_X1 U1281 ( .A1(serve_exception), .A2(\Scc_coproc/cause[5] ), .B1(n7109), .B2(n1038), .ZN(n1037) );
  OAI222_X1 U1282 ( .A1(n364), .A2(n1039), .B1(n366), .B2(n1040), .C1(net55850), .C2(n1041), .ZN(n3885) );
  OAI22_X1 U1283 ( .A1(net55874), .A2(n1040), .B1(net55830), .B2(n1039), .ZN(
        n3886) );
  OAI22_X1 U1285 ( .A1(n7030), .A2(n1042), .B1(n7189), .B2(n1040), .ZN(n3887)
         );
  OAI22_X1 U1287 ( .A1(n372), .A2(n1042), .B1(n1043), .B2(n1044), .ZN(n3888)
         );
  NAND2_X1 U1288 ( .A1(n372), .A2(n6547), .ZN(n1044) );
  OAI221_X1 U1290 ( .B1(n357), .B2(n1041), .C1(n359), .C2(n1045), .A(n1046), 
        .ZN(n3889) );
  AOI22_X1 U1291 ( .A1(\Mcontrol/bvgen/d_curr_pc[0] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [0]), .B2(n362), .ZN(n1046) );
  OAI221_X1 U1294 ( .B1(n357), .B2(n1047), .C1(n6221), .C2(n359), .A(n1048), 
        .ZN(n3890) );
  AOI22_X1 U1295 ( .A1(\Mcontrol/bvgen/d_curr_pc[23] ), .A2(n361), .B1(
        \Mcontrol/bvgen/x_curr_pc [23]), .B2(n362), .ZN(n1048) );
  OAI21_X1 U1298 ( .B1(net55824), .B2(n1052), .A(n1053), .ZN(n3891) );
  OAI22_X1 U1299 ( .A1(net55822), .A2(n1054), .B1(n1055), .B2(net55898), .ZN(
        n3892) );
  NOR2_X1 U1300 ( .A1(n1056), .A2(\Scc_coproc/din_exc_word[4] ), .ZN(n1055) );
  OAI21_X1 U1301 ( .B1(net55824), .B2(n1057), .A(n1053), .ZN(n3893) );
  OAI21_X1 U1302 ( .B1(net55824), .B2(n1058), .A(n1053), .ZN(n3894) );
  OAI21_X1 U1303 ( .B1(n1059), .B2(n1060), .A(net55824), .ZN(n1053) );
  OAI22_X1 U1304 ( .A1(net55822), .A2(n3028), .B1(n1061), .B2(net55902), .ZN(
        n3895) );
  AOI22_X1 U1305 ( .A1(n1056), .A2(n1060), .B1(\Scc_coproc/din_exc_word[5] ), 
        .B2(n1059), .ZN(n1061) );
  INV_X1 U1306 ( .A(n1059), .ZN(n1056) );
  NAND2_X1 U1307 ( .A1(\Scc_coproc/din_exc_word[0] ), .A2(\Scc_coproc/N562 ), 
        .ZN(n1059) );
  OAI21_X1 U1308 ( .B1(n7189), .B2(n1062), .A(n1063), .ZN(n3896) );
  OAI21_X1 U1310 ( .B1(n7189), .B2(n1064), .A(n1063), .ZN(n3897) );
  OAI222_X1 U1312 ( .A1(n364), .A2(n1065), .B1(n366), .B2(n1066), .C1(net55846), .C2(n676), .ZN(n3898) );
  OAI22_X1 U1314 ( .A1(net55874), .A2(n1066), .B1(net55828), .B2(n1065), .ZN(
        n3899) );
  INV_X1 U1317 ( .A(n1067), .ZN(n3900) );
  AOI22_X1 U1318 ( .A1(n7189), .A2(\Mcontrol/f_currpc[10] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[10] ), .ZN(n1067) );
  OAI222_X1 U1319 ( .A1(n364), .A2(n1068), .B1(n366), .B2(n1069), .C1(net55846), .C2(n1047), .ZN(n3901) );
  NAND2_X1 U1321 ( .A1(n1050), .A2(net55824), .ZN(n366) );
  INV_X1 U1322 ( .A(n1051), .ZN(n1050) );
  NAND2_X1 U1323 ( .A1(net55840), .A2(n1051), .ZN(n364) );
  NAND2_X1 U1324 ( .A1(n1070), .A2(\Mcontrol/bvgen/x_jump_type[0] ), .ZN(n1051) );
  INV_X1 U1325 ( .A(\Mcontrol/bvgen/N9 ), .ZN(n1070) );
  OAI22_X1 U1326 ( .A1(net55874), .A2(n1069), .B1(net55826), .B2(n1068), .ZN(
        n3902) );
  INV_X1 U1329 ( .A(n1071), .ZN(n3903) );
  AOI22_X1 U1330 ( .A1(n7189), .A2(\Mcontrol/f_currpc[23] ), .B1(n7030), .B2(
        \Mcontrol/bvgen/d_curr_pc[23] ), .ZN(n1071) );
  INV_X1 U1331 ( .A(n1072), .ZN(n3904) );
  AOI22_X1 U1332 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(net55822), .B1(net55910), .B2(\Mcontrol/bvgen/x_jump_type[0] ), .ZN(n1072) );
  OAI22_X1 U1333 ( .A1(n1073), .A2(net55912), .B1(net55828), .B2(
        \Mcontrol/bvgen/N3 ), .ZN(n3905) );
  INV_X1 U1334 ( .A(\Mcontrol/d_jump_type[2] ), .ZN(n1073) );
  OAI221_X1 U1335 ( .B1(n123), .B2(n232), .C1(\Mpath/the_alu/N55 ), .C2(
        net55852), .A(n1074), .ZN(n3906) );
  AOI22_X1 U1336 ( .A1(n6556), .A2(n670), .B1(n6560), .B2(n1075), .ZN(n1074)
         );
  OAI221_X1 U1337 ( .B1(n175), .B2(n232), .C1(\Mpath/the_alu/N81 ), .C2(
        net55852), .A(n1076), .ZN(n3907) );
  AOI22_X1 U1338 ( .A1(n6556), .A2(n1077), .B1(n6560), .B2(n1078), .ZN(n1076)
         );
  OAI221_X1 U1339 ( .B1(n87), .B2(n232), .C1(\Mpath/the_alu/N37 ), .C2(
        net55854), .A(n1079), .ZN(n3908) );
  AOI22_X1 U1340 ( .A1(n6556), .A2(n1080), .B1(n6560), .B2(n1081), .ZN(n1079)
         );
  OAI221_X1 U1341 ( .B1(n171), .B2(n232), .C1(\Mpath/the_alu/N79 ), .C2(
        net55854), .A(n1082), .ZN(n3909) );
  AOI22_X1 U1342 ( .A1(n6556), .A2(n862), .B1(n6560), .B2(n1083), .ZN(n1082)
         );
  OAI221_X1 U1343 ( .B1(n52), .B2(n232), .C1(\Mpath/the_alu/N21 ), .C2(
        net55854), .A(n1084), .ZN(n3910) );
  AOI22_X1 U1344 ( .A1(n6556), .A2(n1085), .B1(n6560), .B2(n1086), .ZN(n1084)
         );
  OAI221_X1 U1345 ( .B1(n167), .B2(n232), .C1(\Mpath/the_alu/N77 ), .C2(
        net55852), .A(n1087), .ZN(n3911) );
  AOI22_X1 U1346 ( .A1(n6556), .A2(n851), .B1(n6560), .B2(n1088), .ZN(n1087)
         );
  OAI221_X1 U1347 ( .B1(n163), .B2(n232), .C1(\Mpath/the_alu/N75 ), .C2(
        net55850), .A(n1089), .ZN(n3912) );
  AOI22_X1 U1348 ( .A1(n6556), .A2(n840), .B1(n6560), .B2(n1090), .ZN(n1089)
         );
  OAI221_X1 U1349 ( .B1(n147), .B2(n232), .C1(n7184), .C2(net55852), .A(n1091), 
        .ZN(n3913) );
  AOI22_X1 U1350 ( .A1(n6556), .A2(n829), .B1(n6560), .B2(n1092), .ZN(n1091)
         );
  OAI22_X1 U1351 ( .A1(n295), .A2(n1093), .B1(n147), .B2(n297), .ZN(n3914) );
  OAI22_X1 U1353 ( .A1(n295), .A2(n1094), .B1(n163), .B2(n297), .ZN(n3915) );
  OAI22_X1 U1355 ( .A1(n295), .A2(n1095), .B1(n167), .B2(n297), .ZN(n3916) );
  OAI22_X1 U1357 ( .A1(n295), .A2(n1096), .B1(n52), .B2(n297), .ZN(n3917) );
  OAI22_X1 U1359 ( .A1(n295), .A2(n1097), .B1(n59), .B2(n297), .ZN(n3918) );
  OAI22_X1 U1361 ( .A1(n295), .A2(n1098), .B1(n171), .B2(n297), .ZN(n3919) );
  OAI22_X1 U1363 ( .A1(n295), .A2(n1099), .B1(n63), .B2(n297), .ZN(n3920) );
  OAI22_X1 U1365 ( .A1(n295), .A2(n1100), .B1(n67), .B2(n297), .ZN(n3921) );
  OAI22_X1 U1367 ( .A1(n295), .A2(n1101), .B1(n71), .B2(n297), .ZN(n3922) );
  OAI22_X1 U1369 ( .A1(n295), .A2(n1102), .B1(n75), .B2(n297), .ZN(n3923) );
  OAI22_X1 U1371 ( .A1(n295), .A2(n1103), .B1(n87), .B2(n297), .ZN(n3924) );
  OAI22_X1 U1373 ( .A1(n295), .A2(n1104), .B1(n175), .B2(n297), .ZN(n3925) );
  OAI22_X1 U1375 ( .A1(n295), .A2(n1105), .B1(n123), .B2(n297), .ZN(n3926) );
  OAI22_X1 U1377 ( .A1(n295), .A2(n1106), .B1(n179), .B2(n297), .ZN(n3927) );
  OAI22_X1 U1381 ( .A1(n288), .A2(n4864), .B1(n147), .B2(n289), .ZN(n3928) );
  OAI22_X1 U1382 ( .A1(n288), .A2(n4868), .B1(n163), .B2(n289), .ZN(n3929) );
  OAI22_X1 U1383 ( .A1(n288), .A2(n4869), .B1(n167), .B2(n289), .ZN(n3930) );
  OAI22_X1 U1384 ( .A1(n288), .A2(n4870), .B1(n52), .B2(n289), .ZN(n3931) );
  OAI22_X1 U1385 ( .A1(n288), .A2(n4871), .B1(n59), .B2(n289), .ZN(n3932) );
  OAI22_X1 U1386 ( .A1(n288), .A2(n4872), .B1(n171), .B2(n289), .ZN(n3933) );
  OAI22_X1 U1387 ( .A1(n288), .A2(n4873), .B1(n63), .B2(n289), .ZN(n3934) );
  OAI22_X1 U1388 ( .A1(n288), .A2(n4874), .B1(n67), .B2(n289), .ZN(n3935) );
  OAI22_X1 U1389 ( .A1(n288), .A2(n4875), .B1(n71), .B2(n289), .ZN(n3936) );
  OAI22_X1 U1390 ( .A1(n288), .A2(n4876), .B1(n75), .B2(n289), .ZN(n3937) );
  OAI22_X1 U1391 ( .A1(n288), .A2(n4879), .B1(n87), .B2(n289), .ZN(n3938) );
  OAI22_X1 U1392 ( .A1(n288), .A2(n4883), .B1(n175), .B2(n289), .ZN(n3939) );
  OAI22_X1 U1393 ( .A1(n288), .A2(n4889), .B1(n123), .B2(n289), .ZN(n3940) );
  OAI22_X1 U1394 ( .A1(n288), .A2(n4894), .B1(n179), .B2(n289), .ZN(n3941) );
  OAI22_X1 U1397 ( .A1(n282), .A2(n1109), .B1(n147), .B2(n284), .ZN(n3942) );
  OAI22_X1 U1398 ( .A1(n282), .A2(n1110), .B1(n163), .B2(n284), .ZN(n3943) );
  OAI22_X1 U1399 ( .A1(n282), .A2(n1111), .B1(n167), .B2(n284), .ZN(n3944) );
  OAI22_X1 U1400 ( .A1(n282), .A2(n1112), .B1(n52), .B2(n284), .ZN(n3945) );
  OAI22_X1 U1401 ( .A1(n282), .A2(n1113), .B1(n59), .B2(n284), .ZN(n3946) );
  OAI22_X1 U1402 ( .A1(n282), .A2(n1114), .B1(n171), .B2(n284), .ZN(n3947) );
  OAI22_X1 U1403 ( .A1(n282), .A2(n1115), .B1(n63), .B2(n284), .ZN(n3948) );
  OAI22_X1 U1404 ( .A1(n282), .A2(n1116), .B1(n67), .B2(n284), .ZN(n3949) );
  OAI22_X1 U1405 ( .A1(n282), .A2(n1117), .B1(n71), .B2(n284), .ZN(n3950) );
  OAI22_X1 U1406 ( .A1(n282), .A2(n1118), .B1(n75), .B2(n284), .ZN(n3951) );
  OAI22_X1 U1407 ( .A1(n282), .A2(n1119), .B1(n87), .B2(n284), .ZN(n3952) );
  OAI22_X1 U1408 ( .A1(n282), .A2(n1120), .B1(n175), .B2(n284), .ZN(n3953) );
  OAI22_X1 U1409 ( .A1(n282), .A2(n1121), .B1(n123), .B2(n284), .ZN(n3954) );
  OAI22_X1 U1410 ( .A1(n282), .A2(n1122), .B1(n179), .B2(n284), .ZN(n3955) );
  OAI22_X1 U1413 ( .A1(n278), .A2(n4992), .B1(n147), .B2(n7276), .ZN(n3956) );
  OAI22_X1 U1414 ( .A1(n278), .A2(n4996), .B1(n163), .B2(n7276), .ZN(n3957) );
  OAI22_X1 U1415 ( .A1(n278), .A2(n4997), .B1(n167), .B2(n7276), .ZN(n3958) );
  OAI22_X1 U1416 ( .A1(n278), .A2(n4998), .B1(n52), .B2(n7276), .ZN(n3959) );
  OAI22_X1 U1417 ( .A1(n278), .A2(n4999), .B1(n59), .B2(n7276), .ZN(n3960) );
  OAI22_X1 U1418 ( .A1(n278), .A2(n5000), .B1(n171), .B2(n7276), .ZN(n3961) );
  OAI22_X1 U1419 ( .A1(n278), .A2(n5001), .B1(n63), .B2(n7276), .ZN(n3962) );
  OAI22_X1 U1420 ( .A1(n278), .A2(n5002), .B1(n67), .B2(n7276), .ZN(n3963) );
  OAI22_X1 U1421 ( .A1(n278), .A2(n5003), .B1(n71), .B2(n7276), .ZN(n3964) );
  OAI22_X1 U1422 ( .A1(n278), .A2(n5004), .B1(n75), .B2(n7276), .ZN(n3965) );
  OAI22_X1 U1423 ( .A1(n278), .A2(n5007), .B1(n87), .B2(n7276), .ZN(n3966) );
  OAI22_X1 U1424 ( .A1(n278), .A2(n5011), .B1(n175), .B2(n7276), .ZN(n3967) );
  OAI22_X1 U1425 ( .A1(n278), .A2(n5017), .B1(n123), .B2(n7276), .ZN(n3968) );
  OAI22_X1 U1426 ( .A1(n278), .A2(n5022), .B1(n179), .B2(n7276), .ZN(n3969) );
  OAI22_X1 U1429 ( .A1(n272), .A2(n1123), .B1(n147), .B2(n274), .ZN(n3970) );
  OAI22_X1 U1430 ( .A1(n272), .A2(n1124), .B1(n163), .B2(n274), .ZN(n3971) );
  OAI22_X1 U1431 ( .A1(n272), .A2(n1125), .B1(n167), .B2(n274), .ZN(n3972) );
  OAI22_X1 U1432 ( .A1(n272), .A2(n1126), .B1(n52), .B2(n274), .ZN(n3973) );
  OAI22_X1 U1433 ( .A1(n272), .A2(n1127), .B1(n59), .B2(n274), .ZN(n3974) );
  OAI22_X1 U1434 ( .A1(n272), .A2(n1128), .B1(n171), .B2(n274), .ZN(n3975) );
  OAI22_X1 U1435 ( .A1(n272), .A2(n1129), .B1(n63), .B2(n274), .ZN(n3976) );
  OAI22_X1 U1436 ( .A1(n272), .A2(n1130), .B1(n67), .B2(n274), .ZN(n3977) );
  OAI22_X1 U1437 ( .A1(n272), .A2(n1131), .B1(n71), .B2(n274), .ZN(n3978) );
  OAI22_X1 U1438 ( .A1(n272), .A2(n1132), .B1(n75), .B2(n274), .ZN(n3979) );
  OAI22_X1 U1439 ( .A1(n272), .A2(n1133), .B1(n87), .B2(n274), .ZN(n3980) );
  OAI22_X1 U1440 ( .A1(n272), .A2(n1134), .B1(n175), .B2(n274), .ZN(n3981) );
  OAI22_X1 U1441 ( .A1(n272), .A2(n1135), .B1(n123), .B2(n274), .ZN(n3982) );
  OAI22_X1 U1442 ( .A1(n272), .A2(n1136), .B1(n179), .B2(n274), .ZN(n3983) );
  OAI22_X1 U1445 ( .A1(n268), .A2(n5120), .B1(n147), .B2(n269), .ZN(n3984) );
  OAI22_X1 U1446 ( .A1(n268), .A2(n5124), .B1(n163), .B2(n269), .ZN(n3985) );
  OAI22_X1 U1447 ( .A1(n268), .A2(n5125), .B1(n167), .B2(n269), .ZN(n3986) );
  OAI22_X1 U1448 ( .A1(n268), .A2(n5126), .B1(n52), .B2(n269), .ZN(n3987) );
  OAI22_X1 U1449 ( .A1(n268), .A2(n5127), .B1(n59), .B2(n269), .ZN(n3988) );
  OAI22_X1 U1450 ( .A1(n268), .A2(n5128), .B1(n171), .B2(n269), .ZN(n3989) );
  OAI22_X1 U1451 ( .A1(n268), .A2(n5129), .B1(n63), .B2(n269), .ZN(n3990) );
  OAI22_X1 U1452 ( .A1(n268), .A2(n5130), .B1(n67), .B2(n269), .ZN(n3991) );
  OAI22_X1 U1453 ( .A1(n268), .A2(n5131), .B1(n71), .B2(n269), .ZN(n3992) );
  OAI22_X1 U1454 ( .A1(n268), .A2(n5132), .B1(n75), .B2(n269), .ZN(n3993) );
  OAI22_X1 U1455 ( .A1(n268), .A2(n5135), .B1(n87), .B2(n269), .ZN(n3994) );
  OAI22_X1 U1456 ( .A1(n268), .A2(n5139), .B1(n175), .B2(n269), .ZN(n3995) );
  OAI22_X1 U1457 ( .A1(n268), .A2(n5145), .B1(n123), .B2(n269), .ZN(n3996) );
  OAI22_X1 U1458 ( .A1(n268), .A2(n5150), .B1(n179), .B2(n269), .ZN(n3997) );
  OAI22_X1 U1461 ( .A1(n7115), .A2(n5216), .B1(n147), .B2(n262), .ZN(n3998) );
  OAI22_X1 U1462 ( .A1(n7115), .A2(n5220), .B1(n163), .B2(n262), .ZN(n3999) );
  OAI22_X1 U1463 ( .A1(n7115), .A2(n5221), .B1(n167), .B2(n262), .ZN(n4000) );
  OAI22_X1 U1464 ( .A1(n7115), .A2(n5222), .B1(n52), .B2(n262), .ZN(n4001) );
  OAI22_X1 U1465 ( .A1(n7115), .A2(n5223), .B1(n59), .B2(n262), .ZN(n4002) );
  OAI22_X1 U1466 ( .A1(n7115), .A2(n5224), .B1(n171), .B2(n262), .ZN(n4003) );
  OAI22_X1 U1467 ( .A1(n7115), .A2(n5225), .B1(n63), .B2(n262), .ZN(n4004) );
  OAI22_X1 U1468 ( .A1(n7115), .A2(n5226), .B1(n67), .B2(n262), .ZN(n4005) );
  OAI22_X1 U1469 ( .A1(n7115), .A2(n5227), .B1(n71), .B2(n262), .ZN(n4006) );
  OAI22_X1 U1470 ( .A1(n7115), .A2(n5228), .B1(n75), .B2(n262), .ZN(n4007) );
  OAI22_X1 U1471 ( .A1(n7115), .A2(n5231), .B1(n87), .B2(n262), .ZN(n4008) );
  OAI22_X1 U1472 ( .A1(n7115), .A2(n5235), .B1(n175), .B2(n262), .ZN(n4009) );
  OAI22_X1 U1473 ( .A1(n7115), .A2(n5241), .B1(n123), .B2(n262), .ZN(n4010) );
  OAI22_X1 U1474 ( .A1(n7115), .A2(n5246), .B1(n179), .B2(n262), .ZN(n4011) );
  OAI22_X1 U1477 ( .A1(n255), .A2(n1137), .B1(n147), .B2(n257), .ZN(n4012) );
  OAI22_X1 U1479 ( .A1(n255), .A2(n1138), .B1(n163), .B2(n257), .ZN(n4013) );
  OAI22_X1 U1481 ( .A1(n255), .A2(n1139), .B1(n167), .B2(n257), .ZN(n4014) );
  OAI22_X1 U1483 ( .A1(n255), .A2(n1140), .B1(n52), .B2(n257), .ZN(n4015) );
  OAI22_X1 U1485 ( .A1(n255), .A2(n1141), .B1(n59), .B2(n257), .ZN(n4016) );
  OAI22_X1 U1487 ( .A1(n255), .A2(n1142), .B1(n171), .B2(n257), .ZN(n4017) );
  OAI22_X1 U1489 ( .A1(n255), .A2(n1143), .B1(n63), .B2(n257), .ZN(n4018) );
  OAI22_X1 U1491 ( .A1(n255), .A2(n1144), .B1(n67), .B2(n257), .ZN(n4019) );
  OAI22_X1 U1493 ( .A1(n255), .A2(n1145), .B1(n71), .B2(n257), .ZN(n4020) );
  OAI22_X1 U1495 ( .A1(n255), .A2(n1146), .B1(n75), .B2(n257), .ZN(n4021) );
  OAI22_X1 U1497 ( .A1(n255), .A2(n1147), .B1(n87), .B2(n257), .ZN(n4022) );
  OAI22_X1 U1499 ( .A1(n255), .A2(n1148), .B1(n175), .B2(n257), .ZN(n4023) );
  OAI22_X1 U1501 ( .A1(n255), .A2(n1149), .B1(n123), .B2(n257), .ZN(n4024) );
  OAI22_X1 U1503 ( .A1(n255), .A2(n1150), .B1(n179), .B2(n257), .ZN(n4025) );
  OAI22_X1 U1507 ( .A1(n249), .A2(n1151), .B1(n147), .B2(n251), .ZN(n4026) );
  OAI22_X1 U1508 ( .A1(n249), .A2(n1152), .B1(n163), .B2(n251), .ZN(n4027) );
  OAI22_X1 U1509 ( .A1(n249), .A2(n1153), .B1(n167), .B2(n251), .ZN(n4028) );
  OAI22_X1 U1510 ( .A1(n249), .A2(n1154), .B1(n52), .B2(n251), .ZN(n4029) );
  OAI22_X1 U1511 ( .A1(n249), .A2(n1155), .B1(n59), .B2(n251), .ZN(n4030) );
  OAI22_X1 U1512 ( .A1(n249), .A2(n1156), .B1(n171), .B2(n251), .ZN(n4031) );
  OAI22_X1 U1513 ( .A1(n249), .A2(n1157), .B1(n63), .B2(n251), .ZN(n4032) );
  OAI22_X1 U1514 ( .A1(n249), .A2(n1158), .B1(n67), .B2(n251), .ZN(n4033) );
  OAI22_X1 U1515 ( .A1(n249), .A2(n1159), .B1(n71), .B2(n251), .ZN(n4034) );
  OAI22_X1 U1516 ( .A1(n249), .A2(n1160), .B1(n75), .B2(n251), .ZN(n4035) );
  OAI22_X1 U1517 ( .A1(n249), .A2(n1161), .B1(n87), .B2(n251), .ZN(n4036) );
  OAI22_X1 U1518 ( .A1(n249), .A2(n1162), .B1(n175), .B2(n251), .ZN(n4037) );
  OAI22_X1 U1519 ( .A1(n249), .A2(n1163), .B1(n123), .B2(n251), .ZN(n4038) );
  OAI22_X1 U1520 ( .A1(n249), .A2(n1164), .B1(n179), .B2(n251), .ZN(n4039) );
  OAI22_X1 U1523 ( .A1(n243), .A2(n1165), .B1(n147), .B2(n7370), .ZN(n4040) );
  OAI22_X1 U1525 ( .A1(n243), .A2(n1166), .B1(n163), .B2(n7370), .ZN(n4041) );
  OAI22_X1 U1527 ( .A1(n243), .A2(n1167), .B1(n167), .B2(n7370), .ZN(n4042) );
  OAI22_X1 U1529 ( .A1(n243), .A2(n1168), .B1(n52), .B2(n7370), .ZN(n4043) );
  OAI22_X1 U1531 ( .A1(n243), .A2(n1169), .B1(n59), .B2(n7370), .ZN(n4044) );
  OAI22_X1 U1533 ( .A1(n243), .A2(n1170), .B1(n171), .B2(n7370), .ZN(n4045) );
  OAI22_X1 U1535 ( .A1(n243), .A2(n1171), .B1(n63), .B2(n7370), .ZN(n4046) );
  OAI22_X1 U1537 ( .A1(n243), .A2(n1172), .B1(n67), .B2(n7370), .ZN(n4047) );
  OAI22_X1 U1539 ( .A1(n243), .A2(n1173), .B1(n71), .B2(n7370), .ZN(n4048) );
  OAI22_X1 U1541 ( .A1(n243), .A2(n1174), .B1(n75), .B2(n7370), .ZN(n4049) );
  OAI22_X1 U1543 ( .A1(n243), .A2(n1175), .B1(n87), .B2(n7370), .ZN(n4050) );
  OAI22_X1 U1545 ( .A1(n243), .A2(n1176), .B1(n175), .B2(n7370), .ZN(n4051) );
  OAI22_X1 U1547 ( .A1(n243), .A2(n1177), .B1(n123), .B2(n7370), .ZN(n4052) );
  OAI22_X1 U1549 ( .A1(n243), .A2(n1178), .B1(n179), .B2(n7370), .ZN(n4053) );
  OAI22_X1 U1553 ( .A1(n237), .A2(n1179), .B1(n147), .B2(n239), .ZN(n4054) );
  OAI22_X1 U1554 ( .A1(n237), .A2(n1180), .B1(n163), .B2(n239), .ZN(n4055) );
  OAI22_X1 U1555 ( .A1(n237), .A2(n1181), .B1(n167), .B2(n239), .ZN(n4056) );
  OAI22_X1 U1556 ( .A1(n237), .A2(n1182), .B1(n52), .B2(n239), .ZN(n4057) );
  OAI22_X1 U1557 ( .A1(n237), .A2(n1183), .B1(n59), .B2(n239), .ZN(n4058) );
  OAI22_X1 U1558 ( .A1(n237), .A2(n1184), .B1(n171), .B2(n239), .ZN(n4059) );
  OAI22_X1 U1559 ( .A1(n237), .A2(n1185), .B1(n63), .B2(n239), .ZN(n4060) );
  OAI22_X1 U1560 ( .A1(n237), .A2(n1186), .B1(n67), .B2(n239), .ZN(n4061) );
  OAI22_X1 U1561 ( .A1(n237), .A2(n1187), .B1(n71), .B2(n239), .ZN(n4062) );
  OAI22_X1 U1562 ( .A1(n237), .A2(n1188), .B1(n75), .B2(n239), .ZN(n4063) );
  OAI22_X1 U1563 ( .A1(n237), .A2(n1189), .B1(n87), .B2(n239), .ZN(n4064) );
  OAI22_X1 U1564 ( .A1(n237), .A2(n1190), .B1(n175), .B2(n239), .ZN(n4065) );
  OAI22_X1 U1565 ( .A1(n237), .A2(n1191), .B1(n123), .B2(n239), .ZN(n4066) );
  OAI22_X1 U1566 ( .A1(n237), .A2(n1192), .B1(n179), .B2(n239), .ZN(n4067) );
  OAI22_X1 U1569 ( .A1(n314), .A2(n1193), .B1(n147), .B2(n7210), .ZN(n4068) );
  OAI22_X1 U1570 ( .A1(n314), .A2(n1194), .B1(n163), .B2(n7210), .ZN(n4069) );
  OAI22_X1 U1571 ( .A1(n314), .A2(n1195), .B1(n167), .B2(n7210), .ZN(n4070) );
  OAI22_X1 U1572 ( .A1(n314), .A2(n1196), .B1(n52), .B2(n7210), .ZN(n4071) );
  OAI22_X1 U1573 ( .A1(n314), .A2(n1197), .B1(n59), .B2(n7210), .ZN(n4072) );
  OAI22_X1 U1574 ( .A1(n314), .A2(n1198), .B1(n171), .B2(n7210), .ZN(n4073) );
  OAI22_X1 U1575 ( .A1(n314), .A2(n1199), .B1(n63), .B2(n7210), .ZN(n4074) );
  OAI22_X1 U1576 ( .A1(n314), .A2(n1200), .B1(n67), .B2(n7210), .ZN(n4075) );
  OAI22_X1 U1577 ( .A1(n314), .A2(n1201), .B1(n71), .B2(n7210), .ZN(n4076) );
  OAI22_X1 U1578 ( .A1(n314), .A2(n1202), .B1(n75), .B2(n7210), .ZN(n4077) );
  OAI22_X1 U1579 ( .A1(n314), .A2(n1203), .B1(n87), .B2(n7210), .ZN(n4078) );
  OAI22_X1 U1580 ( .A1(n314), .A2(n1204), .B1(n175), .B2(n7210), .ZN(n4079) );
  OAI22_X1 U1581 ( .A1(n314), .A2(n1205), .B1(n123), .B2(n7210), .ZN(n4080) );
  OAI22_X1 U1582 ( .A1(n314), .A2(n1206), .B1(n179), .B2(n7210), .ZN(n4081) );
  OAI22_X1 U1585 ( .A1(n308), .A2(n1207), .B1(n147), .B2(n310), .ZN(n4082) );
  OAI22_X1 U1586 ( .A1(n308), .A2(n1208), .B1(n163), .B2(n310), .ZN(n4083) );
  OAI22_X1 U1587 ( .A1(n308), .A2(n1209), .B1(n167), .B2(n310), .ZN(n4084) );
  OAI22_X1 U1588 ( .A1(n308), .A2(n1210), .B1(n52), .B2(n310), .ZN(n4085) );
  OAI22_X1 U1589 ( .A1(n308), .A2(n1211), .B1(n59), .B2(n310), .ZN(n4086) );
  OAI22_X1 U1590 ( .A1(n308), .A2(n1212), .B1(n171), .B2(n310), .ZN(n4087) );
  OAI22_X1 U1591 ( .A1(n308), .A2(n1213), .B1(n63), .B2(n310), .ZN(n4088) );
  OAI22_X1 U1592 ( .A1(n308), .A2(n1214), .B1(n67), .B2(n310), .ZN(n4089) );
  OAI22_X1 U1593 ( .A1(n308), .A2(n1215), .B1(n71), .B2(n310), .ZN(n4090) );
  OAI22_X1 U1594 ( .A1(n308), .A2(n1216), .B1(n75), .B2(n310), .ZN(n4091) );
  OAI22_X1 U1595 ( .A1(n308), .A2(n1217), .B1(n87), .B2(n310), .ZN(n4092) );
  OAI22_X1 U1596 ( .A1(n308), .A2(n1218), .B1(n175), .B2(n310), .ZN(n4093) );
  OAI22_X1 U1597 ( .A1(n308), .A2(n1219), .B1(n123), .B2(n310), .ZN(n4094) );
  OAI22_X1 U1598 ( .A1(n308), .A2(n1220), .B1(n179), .B2(n310), .ZN(n4095) );
  OAI22_X1 U1601 ( .A1(n304), .A2(n4672), .B1(n147), .B2(n7113), .ZN(n4096) );
  OAI22_X1 U1602 ( .A1(n304), .A2(n4676), .B1(n163), .B2(n7113), .ZN(n4097) );
  OAI22_X1 U1603 ( .A1(n304), .A2(n4677), .B1(n167), .B2(n7113), .ZN(n4098) );
  OAI22_X1 U1604 ( .A1(n304), .A2(n4678), .B1(n52), .B2(n7113), .ZN(n4099) );
  OAI22_X1 U1605 ( .A1(n304), .A2(n4679), .B1(n59), .B2(n7113), .ZN(n4100) );
  OAI22_X1 U1606 ( .A1(n304), .A2(n4680), .B1(n171), .B2(n7113), .ZN(n4101) );
  OAI22_X1 U1607 ( .A1(n304), .A2(n4681), .B1(n63), .B2(n7113), .ZN(n4102) );
  OAI22_X1 U1608 ( .A1(n304), .A2(n4682), .B1(n67), .B2(n7113), .ZN(n4103) );
  OAI22_X1 U1609 ( .A1(n304), .A2(n4683), .B1(n71), .B2(n7113), .ZN(n4104) );
  OAI22_X1 U1610 ( .A1(n304), .A2(n4684), .B1(n75), .B2(n7113), .ZN(n4105) );
  OAI22_X1 U1611 ( .A1(n304), .A2(n4687), .B1(n87), .B2(n7113), .ZN(n4106) );
  OAI22_X1 U1612 ( .A1(n304), .A2(n4691), .B1(n175), .B2(n7113), .ZN(n4107) );
  OAI22_X1 U1613 ( .A1(n304), .A2(n4697), .B1(n123), .B2(n7113), .ZN(n4108) );
  OAI22_X1 U1614 ( .A1(n304), .A2(n4702), .B1(n179), .B2(n7113), .ZN(n4109) );
  OAI22_X1 U1618 ( .A1(n292), .A2(n1223), .B1(n147), .B2(n294), .ZN(n4110) );
  OAI22_X1 U1620 ( .A1(n292), .A2(n1224), .B1(n163), .B2(n294), .ZN(n4111) );
  OAI22_X1 U1622 ( .A1(n292), .A2(n1225), .B1(n167), .B2(n294), .ZN(n4112) );
  OAI22_X1 U1624 ( .A1(n292), .A2(n1226), .B1(n52), .B2(n294), .ZN(n4113) );
  OAI22_X1 U1626 ( .A1(n292), .A2(n1227), .B1(n59), .B2(n294), .ZN(n4114) );
  OAI22_X1 U1628 ( .A1(n292), .A2(n1228), .B1(n171), .B2(n294), .ZN(n4115) );
  OAI22_X1 U1630 ( .A1(n292), .A2(n1229), .B1(n63), .B2(n294), .ZN(n4116) );
  OAI22_X1 U1632 ( .A1(n292), .A2(n1230), .B1(n67), .B2(n294), .ZN(n4117) );
  OAI22_X1 U1634 ( .A1(n292), .A2(n1231), .B1(n71), .B2(n294), .ZN(n4118) );
  OAI22_X1 U1636 ( .A1(n292), .A2(n1232), .B1(n75), .B2(n294), .ZN(n4119) );
  OAI22_X1 U1638 ( .A1(n292), .A2(n1233), .B1(n87), .B2(n294), .ZN(n4120) );
  OAI22_X1 U1640 ( .A1(n292), .A2(n1234), .B1(n175), .B2(n294), .ZN(n4121) );
  OAI22_X1 U1642 ( .A1(n292), .A2(n1235), .B1(n123), .B2(n294), .ZN(n4122) );
  OAI22_X1 U1644 ( .A1(n292), .A2(n1236), .B1(n179), .B2(n294), .ZN(n4123) );
  OAI22_X1 U1649 ( .A1(n298), .A2(n1237), .B1(n147), .B2(n300), .ZN(n4124) );
  OAI22_X1 U1650 ( .A1(n298), .A2(n1238), .B1(n163), .B2(n300), .ZN(n4125) );
  OAI22_X1 U1651 ( .A1(n298), .A2(n1239), .B1(n167), .B2(n300), .ZN(n4126) );
  OAI22_X1 U1652 ( .A1(n298), .A2(n1240), .B1(n52), .B2(n300), .ZN(n4127) );
  OAI22_X1 U1653 ( .A1(n298), .A2(n1241), .B1(n59), .B2(n300), .ZN(n4128) );
  OAI22_X1 U1654 ( .A1(n298), .A2(n1242), .B1(n171), .B2(n300), .ZN(n4129) );
  OAI22_X1 U1655 ( .A1(n298), .A2(n1243), .B1(n63), .B2(n300), .ZN(n4130) );
  OAI22_X1 U1656 ( .A1(n298), .A2(n1244), .B1(n67), .B2(n300), .ZN(n4131) );
  OAI22_X1 U1657 ( .A1(n298), .A2(n1245), .B1(n71), .B2(n300), .ZN(n4132) );
  OAI22_X1 U1658 ( .A1(n298), .A2(n1246), .B1(n75), .B2(n300), .ZN(n4133) );
  OAI22_X1 U1659 ( .A1(n298), .A2(n1247), .B1(n87), .B2(n300), .ZN(n4134) );
  OAI22_X1 U1660 ( .A1(n298), .A2(n1248), .B1(n175), .B2(n300), .ZN(n4135) );
  OAI22_X1 U1661 ( .A1(n298), .A2(n1249), .B1(n123), .B2(n300), .ZN(n4136) );
  OAI22_X1 U1662 ( .A1(n298), .A2(n1250), .B1(n179), .B2(n300), .ZN(n4137) );
  OAI22_X1 U1665 ( .A1(n290), .A2(n4832), .B1(n147), .B2(n291), .ZN(n4138) );
  OAI22_X1 U1666 ( .A1(n290), .A2(n4836), .B1(n163), .B2(n291), .ZN(n4139) );
  OAI22_X1 U1667 ( .A1(n290), .A2(n4837), .B1(n167), .B2(n291), .ZN(n4140) );
  OAI22_X1 U1668 ( .A1(n290), .A2(n4838), .B1(n52), .B2(n291), .ZN(n4141) );
  OAI22_X1 U1669 ( .A1(n290), .A2(n4839), .B1(n59), .B2(n291), .ZN(n4142) );
  OAI22_X1 U1670 ( .A1(n290), .A2(n4840), .B1(n171), .B2(n291), .ZN(n4143) );
  OAI22_X1 U1671 ( .A1(n290), .A2(n4841), .B1(n63), .B2(n291), .ZN(n4144) );
  OAI22_X1 U1672 ( .A1(n290), .A2(n4842), .B1(n67), .B2(n291), .ZN(n4145) );
  OAI22_X1 U1673 ( .A1(n290), .A2(n4843), .B1(n71), .B2(n291), .ZN(n4146) );
  OAI22_X1 U1674 ( .A1(n290), .A2(n4844), .B1(n75), .B2(n291), .ZN(n4147) );
  OAI22_X1 U1675 ( .A1(n290), .A2(n4847), .B1(n87), .B2(n291), .ZN(n4148) );
  OAI22_X1 U1676 ( .A1(n290), .A2(n4851), .B1(n175), .B2(n291), .ZN(n4149) );
  OAI22_X1 U1677 ( .A1(n290), .A2(n4857), .B1(n123), .B2(n291), .ZN(n4150) );
  OAI22_X1 U1678 ( .A1(n290), .A2(n4862), .B1(n179), .B2(n291), .ZN(n4151) );
  OAI22_X1 U1681 ( .A1(n7119), .A2(n1253), .B1(n147), .B2(n287), .ZN(n4152) );
  OAI22_X1 U1682 ( .A1(n7119), .A2(n1254), .B1(n163), .B2(n287), .ZN(n4153) );
  OAI22_X1 U1683 ( .A1(n7119), .A2(n1255), .B1(n167), .B2(n287), .ZN(n4154) );
  OAI22_X1 U1684 ( .A1(n7119), .A2(n1256), .B1(n52), .B2(n287), .ZN(n4155) );
  OAI22_X1 U1685 ( .A1(n7119), .A2(n1257), .B1(n59), .B2(n287), .ZN(n4156) );
  OAI22_X1 U1686 ( .A1(n7119), .A2(n1258), .B1(n171), .B2(n287), .ZN(n4157) );
  OAI22_X1 U1687 ( .A1(n7119), .A2(n1259), .B1(n63), .B2(n287), .ZN(n4158) );
  OAI22_X1 U1688 ( .A1(n7119), .A2(n1260), .B1(n67), .B2(n287), .ZN(n4159) );
  OAI22_X1 U1689 ( .A1(n7119), .A2(n1261), .B1(n71), .B2(n287), .ZN(n4160) );
  OAI22_X1 U1690 ( .A1(n7119), .A2(n1262), .B1(n75), .B2(n287), .ZN(n4161) );
  OAI22_X1 U1691 ( .A1(n7119), .A2(n1263), .B1(n87), .B2(n287), .ZN(n4162) );
  OAI22_X1 U1692 ( .A1(n7119), .A2(n1264), .B1(n175), .B2(n287), .ZN(n4163) );
  OAI22_X1 U1693 ( .A1(n7119), .A2(n1265), .B1(n123), .B2(n287), .ZN(n4164) );
  OAI22_X1 U1694 ( .A1(n7119), .A2(n1266), .B1(n179), .B2(n287), .ZN(n4165) );
  OAI22_X1 U1697 ( .A1(n7122), .A2(n4960), .B1(n147), .B2(n281), .ZN(n4166) );
  OAI22_X1 U1698 ( .A1(n7122), .A2(n4964), .B1(n163), .B2(n281), .ZN(n4167) );
  OAI22_X1 U1699 ( .A1(n7122), .A2(n4965), .B1(n167), .B2(n281), .ZN(n4168) );
  OAI22_X1 U1700 ( .A1(n7122), .A2(n4966), .B1(n52), .B2(n281), .ZN(n4169) );
  OAI22_X1 U1701 ( .A1(n7122), .A2(n4967), .B1(n59), .B2(n281), .ZN(n4170) );
  OAI22_X1 U1702 ( .A1(n7122), .A2(n4968), .B1(n171), .B2(n281), .ZN(n4171) );
  OAI22_X1 U1703 ( .A1(n7122), .A2(n4969), .B1(n63), .B2(n281), .ZN(n4172) );
  OAI22_X1 U1704 ( .A1(n7122), .A2(n4970), .B1(n67), .B2(n281), .ZN(n4173) );
  OAI22_X1 U1705 ( .A1(n7122), .A2(n4971), .B1(n71), .B2(n281), .ZN(n4174) );
  OAI22_X1 U1706 ( .A1(n7122), .A2(n4972), .B1(n75), .B2(n281), .ZN(n4175) );
  OAI22_X1 U1707 ( .A1(n7122), .A2(n4975), .B1(n87), .B2(n281), .ZN(n4176) );
  OAI22_X1 U1708 ( .A1(n7122), .A2(n4979), .B1(n175), .B2(n281), .ZN(n4177) );
  OAI22_X1 U1709 ( .A1(n7122), .A2(n4985), .B1(n123), .B2(n281), .ZN(n4178) );
  OAI22_X1 U1710 ( .A1(n7122), .A2(n4990), .B1(n179), .B2(n281), .ZN(n4179) );
  OAI22_X1 U1713 ( .A1(n275), .A2(n1267), .B1(n147), .B2(n7363), .ZN(n4180) );
  OAI22_X1 U1714 ( .A1(n275), .A2(n1268), .B1(n163), .B2(n7363), .ZN(n4181) );
  OAI22_X1 U1715 ( .A1(n275), .A2(n1269), .B1(n167), .B2(n7363), .ZN(n4182) );
  OAI22_X1 U1716 ( .A1(n275), .A2(n1270), .B1(n52), .B2(n7363), .ZN(n4183) );
  OAI22_X1 U1717 ( .A1(n275), .A2(n1271), .B1(n59), .B2(n7363), .ZN(n4184) );
  OAI22_X1 U1718 ( .A1(n275), .A2(n1272), .B1(n171), .B2(n7363), .ZN(n4185) );
  OAI22_X1 U1719 ( .A1(n275), .A2(n1273), .B1(n63), .B2(n7363), .ZN(n4186) );
  OAI22_X1 U1720 ( .A1(n275), .A2(n1274), .B1(n67), .B2(n7363), .ZN(n4187) );
  OAI22_X1 U1721 ( .A1(n275), .A2(n1275), .B1(n71), .B2(n7363), .ZN(n4188) );
  OAI22_X1 U1722 ( .A1(n275), .A2(n1276), .B1(n75), .B2(n7363), .ZN(n4189) );
  OAI22_X1 U1723 ( .A1(n275), .A2(n1277), .B1(n87), .B2(n7363), .ZN(n4190) );
  OAI22_X1 U1724 ( .A1(n275), .A2(n1278), .B1(n175), .B2(n7363), .ZN(n4191) );
  OAI22_X1 U1725 ( .A1(n275), .A2(n1279), .B1(n123), .B2(n7363), .ZN(n4192) );
  OAI22_X1 U1726 ( .A1(n275), .A2(n1280), .B1(n179), .B2(n7363), .ZN(n4193) );
  OAI22_X1 U1729 ( .A1(n270), .A2(n5088), .B1(n147), .B2(n271), .ZN(n4194) );
  OAI22_X1 U1730 ( .A1(n270), .A2(n5092), .B1(n163), .B2(n271), .ZN(n4195) );
  OAI22_X1 U1731 ( .A1(n270), .A2(n5093), .B1(n167), .B2(n271), .ZN(n4196) );
  OAI22_X1 U1732 ( .A1(n270), .A2(n5094), .B1(n52), .B2(n271), .ZN(n4197) );
  OAI22_X1 U1733 ( .A1(n270), .A2(n5095), .B1(n59), .B2(n271), .ZN(n4198) );
  OAI22_X1 U1734 ( .A1(n270), .A2(n5096), .B1(n171), .B2(n271), .ZN(n4199) );
  OAI22_X1 U1735 ( .A1(n270), .A2(n5097), .B1(n63), .B2(n271), .ZN(n4200) );
  OAI22_X1 U1736 ( .A1(n270), .A2(n5098), .B1(n67), .B2(n271), .ZN(n4201) );
  OAI22_X1 U1737 ( .A1(n270), .A2(n5099), .B1(n71), .B2(n271), .ZN(n4202) );
  OAI22_X1 U1738 ( .A1(n270), .A2(n5100), .B1(n75), .B2(n271), .ZN(n4203) );
  OAI22_X1 U1739 ( .A1(n270), .A2(n5103), .B1(n87), .B2(n271), .ZN(n4204) );
  OAI22_X1 U1740 ( .A1(n270), .A2(n5107), .B1(n175), .B2(n271), .ZN(n4205) );
  OAI22_X1 U1741 ( .A1(n270), .A2(n5113), .B1(n123), .B2(n271), .ZN(n4206) );
  OAI22_X1 U1742 ( .A1(n270), .A2(n5118), .B1(n179), .B2(n271), .ZN(n4207) );
  OAI22_X1 U1745 ( .A1(n263), .A2(n5184), .B1(n147), .B2(n7158), .ZN(n4208) );
  OAI22_X1 U1746 ( .A1(n263), .A2(n5188), .B1(n163), .B2(n7158), .ZN(n4209) );
  OAI22_X1 U1747 ( .A1(n263), .A2(n5189), .B1(n167), .B2(n7158), .ZN(n4210) );
  OAI22_X1 U1748 ( .A1(n263), .A2(n5190), .B1(n52), .B2(n7158), .ZN(n4211) );
  OAI22_X1 U1749 ( .A1(n263), .A2(n5191), .B1(n59), .B2(n7158), .ZN(n4212) );
  OAI22_X1 U1750 ( .A1(n263), .A2(n5192), .B1(n171), .B2(n7158), .ZN(n4213) );
  OAI22_X1 U1751 ( .A1(n263), .A2(n5193), .B1(n63), .B2(n7158), .ZN(n4214) );
  OAI22_X1 U1752 ( .A1(n263), .A2(n5194), .B1(n67), .B2(n7158), .ZN(n4215) );
  OAI22_X1 U1753 ( .A1(n263), .A2(n5195), .B1(n71), .B2(n7158), .ZN(n4216) );
  OAI22_X1 U1754 ( .A1(n263), .A2(n5196), .B1(n75), .B2(n7158), .ZN(n4217) );
  OAI22_X1 U1755 ( .A1(n263), .A2(n5199), .B1(n87), .B2(n7158), .ZN(n4218) );
  OAI22_X1 U1756 ( .A1(n263), .A2(n5203), .B1(n175), .B2(n7158), .ZN(n4219) );
  OAI22_X1 U1757 ( .A1(n263), .A2(n5209), .B1(n123), .B2(n7158), .ZN(n4220) );
  OAI22_X1 U1758 ( .A1(n263), .A2(n5214), .B1(n179), .B2(n7158), .ZN(n4221) );
  OAI22_X1 U1761 ( .A1(n258), .A2(n1281), .B1(n147), .B2(n7117), .ZN(n4222) );
  OAI22_X1 U1762 ( .A1(n258), .A2(n1282), .B1(n163), .B2(n7117), .ZN(n4223) );
  OAI22_X1 U1763 ( .A1(n258), .A2(n1283), .B1(n167), .B2(n7117), .ZN(n4224) );
  OAI22_X1 U1764 ( .A1(n258), .A2(n1284), .B1(n52), .B2(n7117), .ZN(n4225) );
  OAI22_X1 U1765 ( .A1(n258), .A2(n1285), .B1(n59), .B2(n7117), .ZN(n4226) );
  OAI22_X1 U1766 ( .A1(n258), .A2(n1286), .B1(n171), .B2(n7117), .ZN(n4227) );
  OAI22_X1 U1767 ( .A1(n258), .A2(n1287), .B1(n63), .B2(n7117), .ZN(n4228) );
  OAI22_X1 U1768 ( .A1(n258), .A2(n1288), .B1(n67), .B2(n7117), .ZN(n4229) );
  OAI22_X1 U1769 ( .A1(n258), .A2(n1289), .B1(n71), .B2(n7117), .ZN(n4230) );
  OAI22_X1 U1770 ( .A1(n258), .A2(n1290), .B1(n75), .B2(n7117), .ZN(n4231) );
  OAI22_X1 U1771 ( .A1(n258), .A2(n1291), .B1(n87), .B2(n7117), .ZN(n4232) );
  OAI22_X1 U1772 ( .A1(n258), .A2(n1292), .B1(n175), .B2(n7117), .ZN(n4233) );
  OAI22_X1 U1773 ( .A1(n258), .A2(n1293), .B1(n123), .B2(n7117), .ZN(n4234) );
  OAI22_X1 U1774 ( .A1(n258), .A2(n1294), .B1(n179), .B2(n7117), .ZN(n4235) );
  OAI22_X1 U1777 ( .A1(n252), .A2(n1295), .B1(n147), .B2(n7271), .ZN(n4236) );
  OAI22_X1 U1778 ( .A1(n252), .A2(n1296), .B1(n163), .B2(n7271), .ZN(n4237) );
  OAI22_X1 U1779 ( .A1(n252), .A2(n1297), .B1(n167), .B2(n7271), .ZN(n4238) );
  OAI22_X1 U1780 ( .A1(n252), .A2(n1298), .B1(n52), .B2(n7271), .ZN(n4239) );
  OAI22_X1 U1781 ( .A1(n252), .A2(n1299), .B1(n59), .B2(n7271), .ZN(n4240) );
  OAI22_X1 U1782 ( .A1(n252), .A2(n1300), .B1(n171), .B2(n7271), .ZN(n4241) );
  OAI22_X1 U1783 ( .A1(n252), .A2(n1301), .B1(n63), .B2(n7271), .ZN(n4242) );
  OAI22_X1 U1784 ( .A1(n252), .A2(n1302), .B1(n67), .B2(n7271), .ZN(n4243) );
  OAI22_X1 U1785 ( .A1(n252), .A2(n1303), .B1(n71), .B2(n7271), .ZN(n4244) );
  OAI22_X1 U1786 ( .A1(n252), .A2(n1304), .B1(n75), .B2(n7271), .ZN(n4245) );
  OAI22_X1 U1787 ( .A1(n252), .A2(n1305), .B1(n87), .B2(n7271), .ZN(n4246) );
  OAI22_X1 U1788 ( .A1(n252), .A2(n1306), .B1(n175), .B2(n7271), .ZN(n4247) );
  OAI22_X1 U1789 ( .A1(n252), .A2(n1307), .B1(n123), .B2(n7271), .ZN(n4248) );
  OAI22_X1 U1790 ( .A1(n252), .A2(n1308), .B1(n179), .B2(n7271), .ZN(n4249) );
  OAI22_X1 U1793 ( .A1(n246), .A2(n1309), .B1(n147), .B2(n248), .ZN(n4250) );
  OAI22_X1 U1794 ( .A1(n246), .A2(n1310), .B1(n163), .B2(n248), .ZN(n4251) );
  OAI22_X1 U1795 ( .A1(n246), .A2(n1311), .B1(n167), .B2(n248), .ZN(n4252) );
  OAI22_X1 U1796 ( .A1(n246), .A2(n1312), .B1(n52), .B2(n248), .ZN(n4253) );
  OAI22_X1 U1797 ( .A1(n246), .A2(n1313), .B1(n59), .B2(n248), .ZN(n4254) );
  OAI22_X1 U1798 ( .A1(n246), .A2(n1314), .B1(n171), .B2(n248), .ZN(n4255) );
  OAI22_X1 U1799 ( .A1(n246), .A2(n1315), .B1(n63), .B2(n248), .ZN(n4256) );
  OAI22_X1 U1800 ( .A1(n246), .A2(n1316), .B1(n67), .B2(n248), .ZN(n4257) );
  OAI22_X1 U1801 ( .A1(n246), .A2(n1317), .B1(n71), .B2(n248), .ZN(n4258) );
  OAI22_X1 U1802 ( .A1(n246), .A2(n1318), .B1(n75), .B2(n248), .ZN(n4259) );
  OAI22_X1 U1803 ( .A1(n246), .A2(n1319), .B1(n87), .B2(n248), .ZN(n4260) );
  OAI22_X1 U1804 ( .A1(n246), .A2(n1320), .B1(n175), .B2(n248), .ZN(n4261) );
  OAI22_X1 U1805 ( .A1(n246), .A2(n1321), .B1(n123), .B2(n248), .ZN(n4262) );
  OAI22_X1 U1806 ( .A1(n246), .A2(n1322), .B1(n179), .B2(n248), .ZN(n4263) );
  OAI22_X1 U1809 ( .A1(n240), .A2(n1323), .B1(n147), .B2(n7318), .ZN(n4264) );
  OAI22_X1 U1810 ( .A1(n240), .A2(n1324), .B1(n163), .B2(n7318), .ZN(n4265) );
  OAI22_X1 U1811 ( .A1(n240), .A2(n1325), .B1(n167), .B2(n7318), .ZN(n4266) );
  OAI22_X1 U1812 ( .A1(n240), .A2(n1326), .B1(n52), .B2(n7318), .ZN(n4267) );
  OAI22_X1 U1813 ( .A1(n240), .A2(n1327), .B1(n59), .B2(n7318), .ZN(n4268) );
  OAI22_X1 U1814 ( .A1(n240), .A2(n1328), .B1(n171), .B2(n7318), .ZN(n4269) );
  OAI22_X1 U1815 ( .A1(n240), .A2(n1329), .B1(n63), .B2(n7318), .ZN(n4270) );
  OAI22_X1 U1816 ( .A1(n240), .A2(n1330), .B1(n67), .B2(n7318), .ZN(n4271) );
  OAI22_X1 U1817 ( .A1(n240), .A2(n1331), .B1(n71), .B2(n7318), .ZN(n4272) );
  OAI22_X1 U1818 ( .A1(n240), .A2(n1332), .B1(n75), .B2(n7318), .ZN(n4273) );
  OAI22_X1 U1819 ( .A1(n240), .A2(n1333), .B1(n87), .B2(n7318), .ZN(n4274) );
  OAI22_X1 U1820 ( .A1(n240), .A2(n1334), .B1(n175), .B2(n7318), .ZN(n4275) );
  OAI22_X1 U1821 ( .A1(n240), .A2(n1335), .B1(n123), .B2(n7318), .ZN(n4276) );
  OAI22_X1 U1822 ( .A1(n240), .A2(n1336), .B1(n179), .B2(n7318), .ZN(n4277) );
  OAI22_X1 U1825 ( .A1(n317), .A2(n1337), .B1(n147), .B2(n7209), .ZN(n4278) );
  OAI22_X1 U1826 ( .A1(n317), .A2(n1338), .B1(n163), .B2(n7209), .ZN(n4279) );
  OAI22_X1 U1827 ( .A1(n317), .A2(n1339), .B1(n167), .B2(n7209), .ZN(n4280) );
  OAI22_X1 U1828 ( .A1(n317), .A2(n1340), .B1(n52), .B2(n7209), .ZN(n4281) );
  OAI22_X1 U1829 ( .A1(n317), .A2(n1341), .B1(n59), .B2(n7209), .ZN(n4282) );
  OAI22_X1 U1830 ( .A1(n317), .A2(n1342), .B1(n171), .B2(n7209), .ZN(n4283) );
  OAI22_X1 U1831 ( .A1(n317), .A2(n1343), .B1(n63), .B2(n7209), .ZN(n4284) );
  OAI22_X1 U1832 ( .A1(n317), .A2(n1344), .B1(n67), .B2(n7209), .ZN(n4285) );
  OAI22_X1 U1833 ( .A1(n317), .A2(n1345), .B1(n71), .B2(n7209), .ZN(n4286) );
  OAI22_X1 U1834 ( .A1(n317), .A2(n1346), .B1(n75), .B2(n7209), .ZN(n4287) );
  OAI22_X1 U1835 ( .A1(n317), .A2(n1347), .B1(n87), .B2(n7209), .ZN(n4288) );
  OAI22_X1 U1836 ( .A1(n317), .A2(n1348), .B1(n175), .B2(n7209), .ZN(n4289) );
  OAI22_X1 U1837 ( .A1(n317), .A2(n1349), .B1(n123), .B2(n7209), .ZN(n4290) );
  OAI22_X1 U1838 ( .A1(n317), .A2(n1350), .B1(n179), .B2(n7209), .ZN(n4291) );
  OAI22_X1 U1841 ( .A1(n7074), .A2(n1351), .B1(n147), .B2(n313), .ZN(n4292) );
  OAI22_X1 U1842 ( .A1(n7074), .A2(n1352), .B1(n163), .B2(n313), .ZN(n4293) );
  OAI22_X1 U1843 ( .A1(n7074), .A2(n1353), .B1(n167), .B2(n313), .ZN(n4294) );
  OAI22_X1 U1844 ( .A1(n7074), .A2(n1354), .B1(n52), .B2(n313), .ZN(n4295) );
  OAI22_X1 U1845 ( .A1(n7074), .A2(n1355), .B1(n59), .B2(n313), .ZN(n4296) );
  OAI22_X1 U1846 ( .A1(n7074), .A2(n1356), .B1(n171), .B2(n313), .ZN(n4297) );
  OAI22_X1 U1847 ( .A1(n7074), .A2(n1357), .B1(n63), .B2(n313), .ZN(n4298) );
  OAI22_X1 U1848 ( .A1(n7074), .A2(n1358), .B1(n67), .B2(n313), .ZN(n4299) );
  OAI22_X1 U1849 ( .A1(n7074), .A2(n1359), .B1(n71), .B2(n313), .ZN(n4300) );
  OAI22_X1 U1850 ( .A1(n7074), .A2(n1360), .B1(n75), .B2(n313), .ZN(n4301) );
  OAI22_X1 U1851 ( .A1(n7074), .A2(n1361), .B1(n87), .B2(n313), .ZN(n4302) );
  OAI22_X1 U1852 ( .A1(n7074), .A2(n1362), .B1(n175), .B2(n313), .ZN(n4303) );
  OAI22_X1 U1853 ( .A1(n7074), .A2(n1363), .B1(n123), .B2(n313), .ZN(n4304) );
  OAI22_X1 U1854 ( .A1(n7074), .A2(n1364), .B1(n179), .B2(n313), .ZN(n4305) );
  OAI22_X1 U1857 ( .A1(n7112), .A2(n4640), .B1(n147), .B2(n307), .ZN(n4306) );
  OAI22_X1 U1858 ( .A1(n7112), .A2(n4644), .B1(n163), .B2(n307), .ZN(n4307) );
  OAI22_X1 U1859 ( .A1(n7112), .A2(n4645), .B1(n167), .B2(n307), .ZN(n4308) );
  OAI22_X1 U1860 ( .A1(n7112), .A2(n4646), .B1(n52), .B2(n307), .ZN(n4309) );
  OAI22_X1 U1861 ( .A1(n7112), .A2(n4647), .B1(n59), .B2(n307), .ZN(n4310) );
  OAI22_X1 U1862 ( .A1(n7112), .A2(n4648), .B1(n171), .B2(n307), .ZN(n4311) );
  OAI22_X1 U1863 ( .A1(n7112), .A2(n4649), .B1(n63), .B2(n307), .ZN(n4312) );
  OAI22_X1 U1864 ( .A1(n7112), .A2(n4650), .B1(n67), .B2(n307), .ZN(n4313) );
  OAI22_X1 U1865 ( .A1(n7112), .A2(n4651), .B1(n71), .B2(n307), .ZN(n4314) );
  OAI22_X1 U1866 ( .A1(n7112), .A2(n4652), .B1(n75), .B2(n307), .ZN(n4315) );
  OAI22_X1 U1867 ( .A1(n7112), .A2(n4655), .B1(n87), .B2(n307), .ZN(n4316) );
  OAI22_X1 U1868 ( .A1(n7112), .A2(n4659), .B1(n175), .B2(n307), .ZN(n4317) );
  OAI22_X1 U1869 ( .A1(n7112), .A2(n4665), .B1(n123), .B2(n307), .ZN(n4318) );
  OAI22_X1 U1870 ( .A1(n7112), .A2(n4670), .B1(n179), .B2(n307), .ZN(n4319) );
  OAI22_X1 U1873 ( .A1(n6558), .A2(n1365), .B1(n147), .B2(n7076), .ZN(n4320)
         );
  OAI22_X1 U1875 ( .A1(n6558), .A2(n1366), .B1(n163), .B2(n7076), .ZN(n4321)
         );
  OAI22_X1 U1877 ( .A1(n6559), .A2(n1367), .B1(n167), .B2(n7076), .ZN(n4322)
         );
  OAI22_X1 U1879 ( .A1(n6559), .A2(n1368), .B1(n52), .B2(n7076), .ZN(n4323) );
  OAI22_X1 U1881 ( .A1(n6559), .A2(n1369), .B1(n59), .B2(n7076), .ZN(n4324) );
  OAI22_X1 U1883 ( .A1(n6558), .A2(n1370), .B1(n171), .B2(n7076), .ZN(n4325)
         );
  OAI22_X1 U1885 ( .A1(n6558), .A2(n1371), .B1(n63), .B2(n7076), .ZN(n4326) );
  OAI22_X1 U1887 ( .A1(n6559), .A2(n1372), .B1(n67), .B2(n7076), .ZN(n4327) );
  OAI22_X1 U1889 ( .A1(n6559), .A2(n1373), .B1(n71), .B2(n7076), .ZN(n4328) );
  OAI22_X1 U1891 ( .A1(n6558), .A2(n1374), .B1(n75), .B2(n7076), .ZN(n4329) );
  OAI22_X1 U1893 ( .A1(n6558), .A2(n1375), .B1(n87), .B2(n7076), .ZN(n4330) );
  OAI22_X1 U1895 ( .A1(n6559), .A2(n1376), .B1(n175), .B2(n7076), .ZN(n4331)
         );
  OAI22_X1 U1897 ( .A1(n6559), .A2(n1377), .B1(n123), .B2(n7076), .ZN(n4332)
         );
  OAI22_X1 U1899 ( .A1(n6558), .A2(n1378), .B1(n179), .B2(n7076), .ZN(n4333)
         );
  OAI22_X1 U1904 ( .A1(n6895), .A2(n1380), .B1(n147), .B2(n6898), .ZN(n4334)
         );
  OAI211_X1 U1906 ( .C1(n6011), .C2(n653), .A(n654), .B(n1381), .ZN(n830) );
  AOI22_X1 U1907 ( .A1(n656), .A2(n6527), .B1(n1382), .B2(n658), .ZN(n1381) );
  INV_X1 U1908 ( .A(n5530), .ZN(n1382) );
  OAI22_X1 U1909 ( .A1(n6897), .A2(n1383), .B1(n163), .B2(n6898), .ZN(n4335)
         );
  OAI211_X1 U1911 ( .C1(n5745), .C2(n5542), .A(n1384), .B(n1385), .ZN(n841) );
  AOI222_X1 U1912 ( .A1(n913), .A2(n6535), .B1(n6518), .B2(n914), .C1(n915), 
        .C2(n6526), .ZN(n1385) );
  AOI22_X1 U1913 ( .A1(n5823), .A2(n916), .B1(n5820), .B2(n917), .ZN(n1384) );
  OAI22_X1 U1914 ( .A1(n6896), .A2(n1386), .B1(n167), .B2(n6898), .ZN(n4336)
         );
  OAI211_X1 U1916 ( .C1(n5745), .C2(n5545), .A(n1387), .B(n1388), .ZN(n852) );
  AOI222_X1 U1917 ( .A1(n913), .A2(n6533), .B1(n6520), .B2(n914), .C1(n915), 
        .C2(n6528), .ZN(n1388) );
  AOI22_X1 U1918 ( .A1(n5833), .A2(n916), .B1(n5830), .B2(n917), .ZN(n1387) );
  OAI22_X1 U1919 ( .A1(n6896), .A2(n1389), .B1(n52), .B2(n6898), .ZN(n4337) );
  OAI22_X1 U1921 ( .A1(n6895), .A2(n1391), .B1(n59), .B2(n6898), .ZN(n4338) );
  OAI22_X1 U1922 ( .A1(n6895), .A2(n1392), .B1(n171), .B2(n6898), .ZN(n4339)
         );
  OAI211_X1 U1924 ( .C1(n5745), .C2(n5554), .A(n1393), .B(n1394), .ZN(n863) );
  AOI222_X1 U1925 ( .A1(n913), .A2(n6531), .B1(n6522), .B2(n914), .C1(n915), 
        .C2(n6530), .ZN(n1394) );
  AND2_X1 U1926 ( .A1(n917), .A2(n5787), .ZN(n915) );
  AND2_X1 U1927 ( .A1(n5745), .A2(n1395), .ZN(n914) );
  OAI22_X1 U1928 ( .A1(n5938), .A2(n1396), .B1(\Mpath/the_memhandle/N34 ), 
        .B2(n1397), .ZN(n1395) );
  INV_X1 U1929 ( .A(n5786), .ZN(n1397) );
  NOR2_X1 U1930 ( .A1(n1398), .A2(n6000), .ZN(n913) );
  AOI22_X1 U1931 ( .A1(n5858), .A2(n916), .B1(n5855), .B2(n917), .ZN(n1393) );
  INV_X1 U1932 ( .A(n995), .ZN(n917) );
  INV_X1 U1933 ( .A(n1398), .ZN(n916) );
  OAI22_X1 U1934 ( .A1(n6897), .A2(n1399), .B1(n63), .B2(n6898), .ZN(n4340) );
  OAI22_X1 U1935 ( .A1(n6896), .A2(n1400), .B1(n67), .B2(n6898), .ZN(n4341) );
  OAI22_X1 U1936 ( .A1(n6897), .A2(n1401), .B1(n71), .B2(n6898), .ZN(n4342) );
  OAI22_X1 U1937 ( .A1(n6895), .A2(n1402), .B1(n75), .B2(n6898), .ZN(n4343) );
  OAI22_X1 U1938 ( .A1(n6897), .A2(n1403), .B1(n87), .B2(n6898), .ZN(n4344) );
  OAI22_X1 U1940 ( .A1(n6896), .A2(n1405), .B1(n175), .B2(n6898), .ZN(n4345)
         );
  OAI22_X1 U1942 ( .A1(n6896), .A2(n1407), .B1(n123), .B2(n6898), .ZN(n4346)
         );
  OAI211_X1 U1944 ( .C1(n5799), .C2(n653), .A(n654), .B(n1408), .ZN(n671) );
  AOI22_X1 U1945 ( .A1(n656), .A2(n6539), .B1(n1409), .B2(n658), .ZN(n1408) );
  INV_X1 U1946 ( .A(n5745), .ZN(n658) );
  INV_X1 U1947 ( .A(n5605), .ZN(n1409) );
  AND2_X1 U1948 ( .A1(n5746), .A2(n5745), .ZN(n656) );
  NAND2_X1 U1949 ( .A1(n5747), .A2(n5745), .ZN(n653) );
  OAI22_X1 U1950 ( .A1(n6895), .A2(n1410), .B1(n179), .B2(n6898), .ZN(n4347)
         );
  OAI22_X1 U1957 ( .A1(net55872), .A2(n1411), .B1(net55826), .B2(n1412), .ZN(
        n4348) );
  OAI221_X1 U1959 ( .B1(n6052), .B2(n1413), .C1(net55860), .C2(n1411), .A(
        n1414), .ZN(n4349) );
  AOI221_X1 U1960 ( .B1(n1415), .B2(n210), .C1(n1416), .C2(n1417), .A(n1418), 
        .ZN(n1414) );
  INV_X1 U1961 ( .A(n6051), .ZN(n210) );
  OAI22_X1 U1963 ( .A1(net55872), .A2(n1419), .B1(net55830), .B2(n3039), .ZN(
        n4350) );
  OAI221_X1 U1964 ( .B1(n5913), .B2(n1413), .C1(net55860), .C2(n1419), .A(
        n1420), .ZN(n4351) );
  AOI221_X1 U1965 ( .B1(n1415), .B2(n205), .C1(n1416), .C2(n6038), .A(n1418), 
        .ZN(n1420) );
  INV_X1 U1966 ( .A(n6050), .ZN(n205) );
  OAI22_X1 U1968 ( .A1(net55872), .A2(n1421), .B1(net55828), .B2(n3041), .ZN(
        n4352) );
  OAI221_X1 U1969 ( .B1(n5903), .B2(n1413), .C1(net55860), .C2(n1421), .A(
        n1422), .ZN(n4353) );
  AOI221_X1 U1970 ( .B1(n1415), .B2(n200), .C1(n1416), .C2(n1423), .A(n1418), 
        .ZN(n1422) );
  INV_X1 U1971 ( .A(n6048), .ZN(n200) );
  OAI22_X1 U1973 ( .A1(net55874), .A2(n1424), .B1(net55826), .B2(n3043), .ZN(
        n4354) );
  OAI221_X1 U1974 ( .B1(n5892), .B2(n1413), .C1(net55862), .C2(n1424), .A(
        n1425), .ZN(n4355) );
  AOI221_X1 U1975 ( .B1(n1415), .B2(n191), .C1(n1416), .C2(n6040), .A(n1418), 
        .ZN(n1425) );
  INV_X1 U1976 ( .A(n6047), .ZN(n191) );
  OAI22_X1 U1978 ( .A1(net55872), .A2(n1426), .B1(net55826), .B2(n3045), .ZN(
        n4356) );
  OAI221_X1 U1979 ( .B1(n5883), .B2(n1413), .C1(net55860), .C2(n1426), .A(
        n1427), .ZN(n4357) );
  AOI221_X1 U1980 ( .B1(n1415), .B2(n6045), .C1(n1416), .C2(n6041), .A(n1418), 
        .ZN(n1427) );
  NOR4_X1 U1981 ( .A1(n1428), .A2(n6054), .A3(n6053), .A4(
        \Mcontrol/Operation_decoding32/N1970 ), .ZN(n1418) );
  AND2_X1 U1982 ( .A1(net55862), .A2(n1429), .ZN(n1416) );
  OAI21_X1 U1983 ( .B1(n1430), .B2(n1431), .A(n1432), .ZN(n1429) );
  INV_X1 U1984 ( .A(n1433), .ZN(n1432) );
  AOI21_X1 U1985 ( .B1(n1434), .B2(n6076), .A(net57323), .ZN(n1433) );
  NAND3_X1 U1987 ( .A1(n7410), .A2(n7532), .A3(n6055), .ZN(n1437) );
  AOI21_X1 U1988 ( .B1(n1439), .B2(net57341), .A(net55910), .ZN(n1415) );
  OR3_X1 U1989 ( .A1(n1431), .A2(n7598), .A3(n7449), .ZN(n1439) );
  NAND3_X1 U1991 ( .A1(n1440), .A2(n1441), .A3(n6058), .ZN(n1413) );
  INV_X1 U1992 ( .A(n1428), .ZN(n1440) );
  NAND3_X1 U1993 ( .A1(n1436), .A2(net55834), .A3(n1442), .ZN(n1428) );
  NOR3_X1 U1994 ( .A1(n7432), .A2(n7226), .A3(n7449), .ZN(n1436) );
  OAI221_X1 U1995 ( .B1(n5520), .B2(n1443), .C1(\Mpath/the_alu/N468 ), .C2(
        net55852), .A(n1444), .ZN(n4358) );
  NAND3_X1 U1996 ( .A1(n1445), .A2(net57954), .A3(n1446), .ZN(n1444) );
  NAND3_X1 U1997 ( .A1(n1447), .A2(net57368), .A3(n1449), .ZN(n1445) );
  OAI21_X1 U1998 ( .B1(\Mcontrol/Operation_decoding32/N2071 ), .B2(net56922), 
        .A(n1450), .ZN(n1449) );
  OAI21_X1 U1999 ( .B1(n7402), .B2(n7229), .A(n7033), .ZN(n1450) );
  NAND3_X1 U2000 ( .A1(n1451), .A2(\Mcontrol/Operation_decoding32/N2060 ), 
        .A3(n6078), .ZN(n1447) );
  INV_X1 U2001 ( .A(n1452), .ZN(n1451) );
  AOI21_X1 U2002 ( .B1(\Mcontrol/Operation_decoding32/N2047 ), .B2(
        \Mcontrol/Operation_decoding32/N2071 ), .A(net58533), .ZN(n1452) );
  NOR2_X1 U2003 ( .A1(n1453), .A2(n1454), .ZN(n4359) );
  AOI22_X1 U2004 ( .A1(shift_op[0]), .A2(net55870), .B1(net55840), .B2(n1455), 
        .ZN(n1453) );
  INV_X1 U2005 ( .A(n5520), .ZN(n1455) );
  OAI221_X1 U2006 ( .B1(net55834), .B2(\Mcontrol/st_logic/N34 ), .C1(n5520), 
        .C2(net55916), .A(n1456), .ZN(n4360) );
  INV_X1 U2007 ( .A(n1457), .ZN(n4361) );
  AOI22_X1 U2008 ( .A1(n7189), .A2(I_DATA_INBUS[0]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [0]), .ZN(n1457) );
  OAI221_X1 U2009 ( .B1(n5519), .B2(n1443), .C1(\Mpath/the_alu/N467 ), .C2(
        net55852), .A(n1458), .ZN(n4362) );
  NAND4_X1 U2010 ( .A1(n1442), .A2(net55834), .A3(n7402), .A4(n1459), .ZN(
        n1458) );
  OAI21_X1 U2011 ( .B1(\Mcontrol/Operation_decoding32/N2047 ), .B2(
        \Mcontrol/Operation_decoding32/N1922 ), .A(n1460), .ZN(n1459) );
  INV_X1 U2012 ( .A(n1461), .ZN(n1460) );
  INV_X1 U2013 ( .A(n1431), .ZN(n1442) );
  NAND3_X1 U2014 ( .A1(n1434), .A2(net57341), .A3(n6076), .ZN(n1431) );
  NOR2_X1 U2015 ( .A1(n1462), .A2(n1454), .ZN(n4363) );
  AOI22_X1 U2016 ( .A1(shift_op[1]), .A2(net55870), .B1(net55840), .B2(n1463), 
        .ZN(n1462) );
  INV_X1 U2017 ( .A(n5519), .ZN(n1463) );
  OAI221_X1 U2018 ( .B1(net55834), .B2(\Mcontrol/st_logic/N27 ), .C1(n5519), 
        .C2(net55918), .A(n1456), .ZN(n4364) );
  INV_X1 U2019 ( .A(n1464), .ZN(n4365) );
  AOI22_X1 U2020 ( .A1(n7189), .A2(I_DATA_INBUS[1]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [1]), .ZN(n1464) );
  OAI221_X1 U2021 ( .B1(n5518), .B2(n1443), .C1(net55862), .C2(n3049), .A(
        n1465), .ZN(n4366) );
  NOR2_X1 U2022 ( .A1(n1466), .A2(n1454), .ZN(n4367) );
  OAI21_X1 U2023 ( .B1(n1467), .B2(net55918), .A(n1468), .ZN(n1454) );
  INV_X1 U2024 ( .A(n1469), .ZN(n1468) );
  AOI21_X1 U2025 ( .B1(n7415), .B2(n7552), .A(n1471), .ZN(n1467) );
  AOI22_X1 U2026 ( .A1(shift_op[2]), .A2(net55870), .B1(net55840), .B2(n1472), 
        .ZN(n1466) );
  INV_X1 U2027 ( .A(n5518), .ZN(n1472) );
  INV_X1 U2029 ( .A(n1473), .ZN(n4369) );
  AOI22_X1 U2030 ( .A1(n7189), .A2(I_DATA_INBUS[2]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [2]), .ZN(n1473) );
  OAI221_X1 U2031 ( .B1(n5517), .B2(n1443), .C1(net55862), .C2(n3051), .A(
        n1465), .ZN(n4370) );
  NAND3_X1 U2032 ( .A1(n6960), .A2(n1461), .A3(n1446), .ZN(n1465) );
  AOI21_X1 U2034 ( .B1(n7236), .B2(net55824), .A(n1469), .ZN(n1456) );
  OAI21_X1 U2035 ( .B1(n6960), .B2(net55918), .A(n1443), .ZN(n1469) );
  INV_X1 U2036 ( .A(n1475), .ZN(n4372) );
  AOI22_X1 U2037 ( .A1(n7189), .A2(I_DATA_INBUS[3]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [3]), .ZN(n1475) );
  NAND3_X1 U2039 ( .A1(n1434), .A2(n1477), .A3(n1446), .ZN(n1476) );
  NAND3_X1 U2040 ( .A1(n6075), .A2(n7598), .A3(n7420), .ZN(n1477) );
  OAI22_X1 U2041 ( .A1(net55824), .A2(n3054), .B1(n5516), .B2(n1479), .ZN(
        n4374) );
  INV_X1 U2042 ( .A(n1480), .ZN(n4375) );
  AOI22_X1 U2043 ( .A1(n7189), .A2(I_DATA_INBUS[4]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [4]), .ZN(n1480) );
  OAI221_X1 U2044 ( .B1(n5515), .B2(n1443), .C1(\Mpath/the_alu/N466 ), .C2(
        net55856), .A(n1481), .ZN(n4376) );
  OAI211_X1 U2045 ( .C1(n7587), .C2(n1461), .A(net55834), .B(net56982), .ZN(
        n1481) );
  OAI21_X1 U2046 ( .B1(n6077), .B2(n6075), .A(n7598), .ZN(n1461) );
  NAND2_X1 U2047 ( .A1(net55840), .A2(net56846), .ZN(n1443) );
  OAI22_X1 U2048 ( .A1(net55822), .A2(n3056), .B1(n5515), .B2(n1479), .ZN(
        n4377) );
  NAND3_X1 U2049 ( .A1(n6960), .A2(n1471), .A3(n1446), .ZN(n1479) );
  NOR2_X1 U2050 ( .A1(net55870), .A2(net56846), .ZN(n1446) );
  INV_X1 U2051 ( .A(n1483), .ZN(n4378) );
  AOI22_X1 U2052 ( .A1(n7189), .A2(I_DATA_INBUS[5]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [5]), .ZN(n1483) );
  INV_X1 U2053 ( .A(n1484), .ZN(n4379) );
  AOI22_X1 U2054 ( .A1(n7189), .A2(I_DATA_INBUS[6]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [6]), .ZN(n1484) );
  INV_X1 U2055 ( .A(n1485), .ZN(n4380) );
  AOI22_X1 U2056 ( .A1(n7189), .A2(I_DATA_INBUS[7]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [7]), .ZN(n1485) );
  INV_X1 U2057 ( .A(n1486), .ZN(n4381) );
  AOI22_X1 U2058 ( .A1(n7189), .A2(I_DATA_INBUS[8]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [8]), .ZN(n1486) );
  INV_X1 U2059 ( .A(n1487), .ZN(n4382) );
  AOI22_X1 U2060 ( .A1(n7189), .A2(I_DATA_INBUS[9]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [9]), .ZN(n1487) );
  INV_X1 U2061 ( .A(n1488), .ZN(n4383) );
  AOI22_X1 U2062 ( .A1(n7189), .A2(I_DATA_INBUS[10]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [10]), .ZN(n1488) );
  INV_X1 U2063 ( .A(n1489), .ZN(n4384) );
  AOI22_X1 U2064 ( .A1(n7189), .A2(I_DATA_INBUS[11]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [11]), .ZN(n1489) );
  INV_X1 U2065 ( .A(n1490), .ZN(n4385) );
  AOI22_X1 U2066 ( .A1(n7189), .A2(I_DATA_INBUS[12]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [12]), .ZN(n1490) );
  INV_X1 U2067 ( .A(n1491), .ZN(n4386) );
  AOI22_X1 U2068 ( .A1(n7189), .A2(I_DATA_INBUS[13]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [13]), .ZN(n1491) );
  INV_X1 U2069 ( .A(n1492), .ZN(n4387) );
  AOI22_X1 U2070 ( .A1(n7189), .A2(I_DATA_INBUS[14]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [14]), .ZN(n1492) );
  INV_X1 U2071 ( .A(n1493), .ZN(n4388) );
  AOI22_X1 U2072 ( .A1(n7189), .A2(I_DATA_INBUS[15]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [15]), .ZN(n1493) );
  INV_X1 U2073 ( .A(n1494), .ZN(n4389) );
  AOI22_X1 U2074 ( .A1(n7189), .A2(I_DATA_INBUS[16]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [16]), .ZN(n1494) );
  OAI22_X1 U2075 ( .A1(n1495), .A2(net55912), .B1(net55826), .B2(
        \Mcontrol/bvgen/N4 ), .ZN(n4390) );
  INV_X1 U2076 ( .A(n6953), .ZN(n1495) );
  INV_X1 U2077 ( .A(n1496), .ZN(n4391) );
  AOI22_X1 U2078 ( .A1(n7189), .A2(I_DATA_INBUS[17]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [17]), .ZN(n1496) );
  INV_X1 U2079 ( .A(n1497), .ZN(n4392) );
  AOI22_X1 U2080 ( .A1(n7189), .A2(I_DATA_INBUS[18]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [18]), .ZN(n1497) );
  INV_X1 U2083 ( .A(n1499), .ZN(n4394) );
  AOI22_X1 U2084 ( .A1(n7189), .A2(I_DATA_INBUS[19]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [19]), .ZN(n1499) );
  OAI22_X1 U2085 ( .A1(net55872), .A2(n1500), .B1(net55826), .B2(n3072), .ZN(
        n4395) );
  INV_X1 U2086 ( .A(n1501), .ZN(n4396) );
  AOI22_X1 U2087 ( .A1(n7189), .A2(I_DATA_INBUS[20]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [20]), .ZN(n1501) );
  INV_X1 U2088 ( .A(n1502), .ZN(n4397) );
  AOI22_X1 U2089 ( .A1(n7189), .A2(I_DATA_INBUS[21]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [21]), .ZN(n1502) );
  INV_X1 U2090 ( .A(n1503), .ZN(n4398) );
  AOI22_X1 U2091 ( .A1(n7189), .A2(I_DATA_INBUS[22]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [22]), .ZN(n1503) );
  INV_X1 U2092 ( .A(n1504), .ZN(n4399) );
  AOI22_X1 U2093 ( .A1(n7189), .A2(I_DATA_INBUS[23]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [23]), .ZN(n1504) );
  INV_X1 U2094 ( .A(n1505), .ZN(n4400) );
  AOI22_X1 U2095 ( .A1(n7189), .A2(I_DATA_INBUS[24]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [24]), .ZN(n1505) );
  INV_X1 U2096 ( .A(n1506), .ZN(n4401) );
  AOI22_X1 U2097 ( .A1(n7189), .A2(I_DATA_INBUS[25]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [25]), .ZN(n1506) );
  NOR2_X1 U2098 ( .A1(n1507), .A2(n1508), .ZN(n4402) );
  AOI22_X1 U2099 ( .A1(exe_outsel[0]), .A2(net55870), .B1(net55840), .B2(n7160), .ZN(n1508) );
  NOR2_X1 U2101 ( .A1(n1507), .A2(n1510), .ZN(n4403) );
  AOI22_X1 U2102 ( .A1(exe_outsel[1]), .A2(net55872), .B1(net55840), .B2(n7042), .ZN(n1510) );
  NOR2_X1 U2104 ( .A1(n1507), .A2(n1512), .ZN(n4404) );
  AOI22_X1 U2105 ( .A1(exe_outsel[2]), .A2(net55872), .B1(net55840), .B2(n7427), .ZN(n1512) );
  AND3_X1 U2107 ( .A1(net56982), .A2(n7159), .A3(n1514), .ZN(n1507) );
  NOR3_X1 U2108 ( .A1(net55864), .A2(n7587), .A3(n7432), .ZN(n1514) );
  OAI22_X1 U2109 ( .A1(net55874), .A2(n1515), .B1(net55826), .B2(
        \Mcontrol/N17 ), .ZN(n4405) );
  OAI22_X1 U2110 ( .A1(net55824), .A2(n1515), .B1(n1516), .B2(net55900), .ZN(
        n4406) );
  NOR2_X1 U2111 ( .A1(n1517), .A2(n1518), .ZN(n1516) );
  OAI22_X1 U2113 ( .A1(n5505), .A2(net55914), .B1(net55828), .B2(
        \Mpath/the_memhandle/N236 ), .ZN(n4407) );
  OAI22_X1 U2114 ( .A1(net55822), .A2(n1519), .B1(n1520), .B2(net55900), .ZN(
        n4408) );
  NOR3_X1 U2115 ( .A1(n1521), .A2(n1522), .A3(n1523), .ZN(n1520) );
  NOR3_X1 U2116 ( .A1(n1524), .A2(n7530), .A3(n7531), .ZN(n1522) );
  OR3_X1 U2117 ( .A1(n7529), .A2(n7226), .A3(n7456), .ZN(n1521) );
  OAI22_X1 U2118 ( .A1(n4508), .A2(net55912), .B1(net55828), .B2(
        \Mpath/the_memhandle/N238 ), .ZN(n4409) );
  OAI22_X1 U2119 ( .A1(net55822), .A2(n1526), .B1(n1527), .B2(net55900), .ZN(
        n4410) );
  NOR4_X1 U2120 ( .A1(n7226), .A2(n1528), .A3(n1523), .A4(n7530), .ZN(n1527)
         );
  NOR3_X1 U2121 ( .A1(n1529), .A2(n7529), .A3(n7456), .ZN(n1528) );
  NOR3_X1 U2122 ( .A1(n1524), .A2(n7510), .A3(n7531), .ZN(n1529) );
  INV_X1 U2123 ( .A(\Mcontrol/Operation_decoding32/N1987 ), .ZN(n1524) );
  OAI22_X1 U2124 ( .A1(n4507), .A2(net55914), .B1(n5745), .B2(net55836), .ZN(
        n4411) );
  OAI22_X1 U2125 ( .A1(net55824), .A2(n1530), .B1(n1531), .B2(net55902), .ZN(
        n4412) );
  NOR2_X1 U2126 ( .A1(n1532), .A2(n7174), .ZN(n1531) );
  INV_X1 U2127 ( .A(n1533), .ZN(n1532) );
  OAI22_X1 U2128 ( .A1(net55822), .A2(n3083), .B1(n187), .B2(net55898), .ZN(
        n4413) );
  AND3_X1 U2129 ( .A1(n7174), .A2(n1534), .A3(n1533), .ZN(n187) );
  NAND3_X1 U2130 ( .A1(\Mcontrol/Operation_decoding32/N1975 ), .A2(n7510), 
        .A3(n7378), .ZN(n1534) );
  OAI22_X1 U2131 ( .A1(net55824), .A2(\Mpath/the_memhandle/N235 ), .B1(n1535), 
        .B2(net55902), .ZN(n4414) );
  NOR2_X1 U2132 ( .A1(\Mcontrol/x_sampled_dmem_command[SIGN] ), .A2(
        \Mcontrol/x_sampled_dwe ), .ZN(n1535) );
  INV_X1 U2133 ( .A(n1536), .ZN(n4415) );
  AOI22_X1 U2134 ( .A1(net55864), .A2(\Mcontrol/x_sampled_dmem_command[SIGN] ), 
        .B1(n1537), .B2(net55834), .ZN(n1536) );
  OAI21_X1 U2135 ( .B1(n1538), .B2(n7456), .A(n1533), .ZN(n1537) );
  AOI21_X1 U2136 ( .B1(\Mcontrol/Operation_decoding32/N2005 ), .B2(net57379), 
        .A(n7522), .ZN(n1538) );
  OAI22_X1 U2137 ( .A1(n7030), .A2(n1539), .B1(n7189), .B2(n3085), .ZN(n4416)
         );
  INV_X1 U2138 ( .A(I_DATA_INBUS[26]), .ZN(n1539) );
  OAI22_X1 U2139 ( .A1(n7030), .A2(n1540), .B1(n7189), .B2(n3086), .ZN(n4417)
         );
  INV_X1 U2140 ( .A(I_DATA_INBUS[27]), .ZN(n1540) );
  OAI22_X1 U2141 ( .A1(n7030), .A2(n1541), .B1(n7189), .B2(n3087), .ZN(n4418)
         );
  INV_X1 U2142 ( .A(I_DATA_INBUS[28]), .ZN(n1541) );
  INV_X1 U2143 ( .A(n1542), .ZN(n4419) );
  AOI22_X1 U2144 ( .A1(n7189), .A2(I_DATA_INBUS[29]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [29]), .ZN(n1542) );
  INV_X1 U2145 ( .A(n1543), .ZN(n4420) );
  AOI22_X1 U2146 ( .A1(n7189), .A2(I_DATA_INBUS[30]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [30]), .ZN(n1543) );
  INV_X1 U2147 ( .A(n1544), .ZN(n4421) );
  AOI22_X1 U2148 ( .A1(n7189), .A2(I_DATA_INBUS[31]), .B1(n7030), .B2(
        \Mcontrol/d_sampled_finstr [31]), .ZN(n1544) );
  OAI22_X1 U2149 ( .A1(net55822), .A2(\Mcontrol/bp_logicA/N14 ), .B1(n1545), 
        .B2(net55900), .ZN(n4422) );
  NOR2_X1 U2150 ( .A1(n7110), .A2(\Mcontrol/x_sampled_dwe ), .ZN(n1545) );
  OAI22_X1 U2151 ( .A1(net55822), .A2(n1546), .B1(n1547), .B2(net55904), .ZN(
        n4423) );
  AND3_X1 U2152 ( .A1(n1548), .A2(n7207), .A3(\Mcontrol/stall_decode ), .ZN(
        n1547) );
  INV_X1 U2153 ( .A(n1549), .ZN(n1548) );
  OAI22_X1 U2154 ( .A1(n7207), .A2(n7189), .B1(n1550), .B2(n7030), .ZN(n4424)
         );
  NOR2_X1 U2155 ( .A1(n6102), .A2(n1549), .ZN(n1550) );
  NAND2_X1 U2156 ( .A1(n6545), .A2(serve_exception), .ZN(n1549) );
  OAI22_X1 U2157 ( .A1(n7110), .A2(net55914), .B1(n6102), .B2(net55836), .ZN(
        n4425) );
  OAI22_X1 U2158 ( .A1(net55822), .A2(n1551), .B1(n1552), .B2(n1553), .ZN(
        n4426) );
  OAI21_X1 U2159 ( .B1(n1554), .B2(n1060), .A(net55824), .ZN(n1553) );
  OR4_X1 U2160 ( .A1(n1517), .A2(\Mcontrol/Operation_decoding32/N89 ), .A3(
        n5743), .A4(net57730), .ZN(n1060) );
  INV_X1 U2161 ( .A(\Scc_coproc/N562 ), .ZN(n1554) );
  OAI21_X1 U2162 ( .B1(n7189), .B2(n1552), .A(n1063), .ZN(n4427) );
  NAND3_X1 U2163 ( .A1(n1043), .A2(n7189), .A3(n1555), .ZN(n1063) );
  INV_X1 U2164 ( .A(n871), .ZN(n1555) );
  AOI22_X1 U2167 ( .A1(epc[1]), .A2(n1562), .B1(n1563), .B2(n7586), .ZN(n1558)
         );
  INV_X1 U2168 ( .A(branch_rega[1]), .ZN(n1556) );
  INV_X1 U2170 ( .A(n1566), .ZN(n1565) );
  OAI221_X1 U2175 ( .B1(n1567), .B2(n214), .C1(\Mpath/the_alu/N82 ), .C2(
        net55852), .A(n1568), .ZN(n4428) );
  AOI222_X1 U2176 ( .A1(n197), .A2(n177), .B1(n192), .B2(n1077), .C1(n195), 
        .C2(n1406), .ZN(n1568) );
  OAI222_X1 U2177 ( .A1(n1569), .A2(n995), .B1(n1570), .B2(n1398), .C1(n5745), 
        .C2(n5587), .ZN(n1406) );
  AOI221_X1 U2178 ( .B1(n6536), .B2(n1571), .C1(n6529), .C2(n1572), .A(n5937), 
        .ZN(n1570) );
  AOI221_X1 U2179 ( .B1(n5786), .B2(n6542), .C1(n5787), .C2(n6532), .A(n5935), 
        .ZN(n1569) );
  INV_X1 U2180 ( .A(n7586), .ZN(n1567) );
  OAI22_X1 U2181 ( .A1(n5587), .A2(net55842), .B1(n174), .B2(net55904), .ZN(
        n4429) );
  INV_X1 U2182 ( .A(n1077), .ZN(n174) );
  OAI222_X1 U2183 ( .A1(n1573), .A2(n323), .B1(n6087), .B2(n402), .C1(n1574), 
        .C2(n322), .ZN(n1077) );
  INV_X1 U2184 ( .A(n6092), .ZN(n1574) );
  OAI22_X1 U2185 ( .A1(n5735), .A2(net55914), .B1(net55826), .B2(n1575), .ZN(
        n4430) );
  OAI22_X1 U2186 ( .A1(n5736), .A2(n626), .B1(n5735), .B2(n627), .ZN(n4431) );
  OAI222_X1 U2187 ( .A1(n628), .A2(n1575), .B1(n5735), .B2(n629), .C1(n5736), 
        .C2(n359), .ZN(n4432) );
  OAI22_X1 U2189 ( .A1(n5554), .A2(net55842), .B1(n170), .B2(net55906), .ZN(
        n4433) );
  INV_X1 U2190 ( .A(n862), .ZN(n170) );
  OAI222_X1 U2191 ( .A1(n1576), .A2(n323), .B1(n6209), .B2(n402), .C1(n1577), 
        .C2(n322), .ZN(n862) );
  INV_X1 U2192 ( .A(n6213), .ZN(n1577) );
  INV_X1 U2193 ( .A(n6212), .ZN(n1576) );
  OAI22_X1 U2194 ( .A1(n6484), .A2(n7110), .B1(serve_exception), .B2(n47), 
        .ZN(n4434) );
  AOI22_X1 U2195 ( .A1(\Scc_coproc/x_exc_word[2] ), .A2(n883), .B1(n1578), 
        .B2(n885), .ZN(n47) );
  NOR3_X1 U2196 ( .A1(\Scc_coproc/interrupt[8] ), .A2(
        \Scc_coproc/interrupt[9] ), .A3(n1579), .ZN(n885) );
  OAI21_X1 U2197 ( .B1(n1580), .B2(\Scc_coproc/interrupt[3] ), .A(n1581), .ZN(
        n1578) );
  OAI22_X1 U2198 ( .A1(n5733), .A2(net55914), .B1(net55828), .B2(n1582), .ZN(
        n4435) );
  OAI22_X1 U2199 ( .A1(n5734), .A2(n626), .B1(n5733), .B2(n627), .ZN(n4436) );
  OAI222_X1 U2200 ( .A1(n628), .A2(n1582), .B1(n5733), .B2(n629), .C1(n5734), 
        .C2(n359), .ZN(n4437) );
  OAI22_X1 U2202 ( .A1(n5545), .A2(net55842), .B1(n166), .B2(net55906), .ZN(
        n4438) );
  INV_X1 U2203 ( .A(n851), .ZN(n166) );
  OAI222_X1 U2204 ( .A1(n1583), .A2(n323), .B1(n6194), .B2(n402), .C1(n1584), 
        .C2(n322), .ZN(n851) );
  INV_X1 U2205 ( .A(n6198), .ZN(n1584) );
  INV_X1 U2206 ( .A(n6197), .ZN(n1583) );
  OAI22_X1 U2207 ( .A1(n6482), .A2(n7110), .B1(serve_exception), .B2(n46), 
        .ZN(n4439) );
  AOI21_X1 U2208 ( .B1(n1585), .B2(n1586), .A(n1587), .ZN(n46) );
  INV_X1 U2209 ( .A(n1588), .ZN(n1586) );
  AOI21_X1 U2210 ( .B1(n883), .B2(\Scc_coproc/x_exc_word[3] ), .A(n1589), .ZN(
        n1588) );
  AOI21_X1 U2211 ( .B1(n1590), .B2(n1591), .A(n1579), .ZN(n1589) );
  OAI22_X1 U2212 ( .A1(n5731), .A2(net55912), .B1(net55826), .B2(n1592), .ZN(
        n4440) );
  OAI22_X1 U2213 ( .A1(n5732), .A2(n626), .B1(n5731), .B2(n627), .ZN(n4441) );
  OAI222_X1 U2214 ( .A1(n628), .A2(n1592), .B1(n5731), .B2(n629), .C1(n5732), 
        .C2(n359), .ZN(n4442) );
  OAI22_X1 U2216 ( .A1(n5542), .A2(net55842), .B1(n162), .B2(net55906), .ZN(
        n4443) );
  INV_X1 U2217 ( .A(n840), .ZN(n162) );
  OAI222_X1 U2218 ( .A1(n1593), .A2(n323), .B1(n6180), .B2(n402), .C1(n1594), 
        .C2(n322), .ZN(n840) );
  INV_X1 U2219 ( .A(n6184), .ZN(n1594) );
  INV_X1 U2220 ( .A(n6183), .ZN(n1593) );
  INV_X1 U2221 ( .A(n1595), .ZN(n4444) );
  AOI22_X1 U2222 ( .A1(serve_exception), .A2(\Scc_coproc/cause[4] ), .B1(n7109), .B2(n1596), .ZN(n1595) );
  OAI22_X1 U2223 ( .A1(n5723), .A2(net55916), .B1(net55828), .B2(n1597), .ZN(
        n4445) );
  OAI22_X1 U2224 ( .A1(n5724), .A2(n626), .B1(n5723), .B2(n627), .ZN(n4446) );
  AND2_X1 U2225 ( .A1(D_BUSY), .A2(n1598), .ZN(n627) );
  OR4_X1 U2226 ( .A1(n1599), .A2(n1600), .A3(n7110), .A4(n373), .ZN(n626) );
  OAI222_X1 U2227 ( .A1(n628), .A2(n1597), .B1(n5723), .B2(n629), .C1(n5724), 
        .C2(n359), .ZN(n4447) );
  OAI21_X1 U2228 ( .B1(n1601), .B2(n1602), .A(D_BUSY), .ZN(n629) );
  NOR3_X1 U2229 ( .A1(n1579), .A2(\Scc_coproc/x_status[14] ), .A3(
        serve_exception), .ZN(n1601) );
  OR2_X1 U2231 ( .A1(n1603), .A2(n357), .ZN(n628) );
  OAI22_X1 U2232 ( .A1(n5530), .A2(net55844), .B1(n146), .B2(net55898), .ZN(
        n4448) );
  INV_X1 U2233 ( .A(n829), .ZN(n146) );
  OAI222_X1 U2234 ( .A1(n1604), .A2(n323), .B1(n6127), .B2(n402), .C1(n1605), 
        .C2(n322), .ZN(n829) );
  INV_X1 U2235 ( .A(n6131), .ZN(n1605) );
  INV_X1 U2236 ( .A(n6130), .ZN(n1604) );
  OAI22_X1 U2237 ( .A1(n5740), .A2(net55914), .B1(net55826), .B2(n1603), .ZN(
        n4449) );
  OAI21_X1 U2239 ( .B1(n5740), .B2(n1606), .A(n1607), .ZN(n4450) );
  OR4_X1 U2240 ( .A1(n1598), .A2(n1600), .A3(\Scc_coproc/N601 ), .A4(n5739), 
        .ZN(n1607) );
  NAND3_X1 U2241 ( .A1(n1599), .A2(n6547), .A3(serve_exception), .ZN(n1598) );
  NOR2_X1 U2242 ( .A1(n1608), .A2(n1600), .ZN(n1606) );
  AOI211_X1 U2243 ( .C1(n1609), .C2(n1599), .A(n373), .B(n7110), .ZN(n1608) );
  NAND3_X1 U2244 ( .A1(n6545), .A2(n7207), .A3(\Mcontrol/stall_decode ), .ZN(
        n1599) );
  INV_X1 U2245 ( .A(\Scc_coproc/N601 ), .ZN(n1609) );
  OAI211_X1 U2246 ( .C1(n5739), .C2(n359), .A(n357), .B(n1049), .ZN(n4451) );
  NAND2_X1 U2247 ( .A1(n1602), .A2(D_BUSY), .ZN(n1049) );
  NOR2_X1 U2248 ( .A1(n1610), .A2(serve_exception), .ZN(n1602) );
  INV_X1 U2251 ( .A(D_BUSY), .ZN(n1600) );
  OAI22_X1 U2252 ( .A1(n5605), .A2(net55844), .B1(n122), .B2(net55900), .ZN(
        n4452) );
  INV_X1 U2253 ( .A(n670), .ZN(n122) );
  OAI222_X1 U2254 ( .A1(n1611), .A2(n323), .B1(n6341), .B2(n402), .C1(n1612), 
        .C2(n322), .ZN(n670) );
  INV_X1 U2255 ( .A(n6345), .ZN(n1612) );
  INV_X1 U2256 ( .A(n6344), .ZN(n1611) );
  OAI221_X1 U2257 ( .B1(n75), .B2(n232), .C1(\Mpath/the_alu/N31 ), .C2(
        net55850), .A(n1613), .ZN(n4453) );
  AOI22_X1 U2258 ( .A1(n6556), .A2(n225), .B1(n6560), .B2(n1614), .ZN(n1613)
         );
  OAI221_X1 U2260 ( .B1(n5857), .B2(n320), .C1(n5745), .C2(n5566), .A(n321), 
        .ZN(n222) );
  OAI22_X1 U2261 ( .A1(n5566), .A2(net55842), .B1(n74), .B2(net55904), .ZN(
        n4454) );
  INV_X1 U2262 ( .A(n225), .ZN(n74) );
  OAI22_X1 U2263 ( .A1(n5690), .A2(n322), .B1(n5691), .B2(n323), .ZN(n225) );
  OAI221_X1 U2264 ( .B1(n71), .B2(n6554), .C1(\Mpath/the_alu/N29 ), .C2(
        net55850), .A(n1615), .ZN(n4455) );
  AOI22_X1 U2265 ( .A1(n6556), .A2(n211), .B1(n6560), .B2(n1616), .ZN(n1615)
         );
  OAI221_X1 U2267 ( .B1(n5832), .B2(n320), .C1(n5745), .C2(n5563), .A(n321), 
        .ZN(n216) );
  OAI22_X1 U2268 ( .A1(n5563), .A2(net55842), .B1(n70), .B2(net55908), .ZN(
        n4456) );
  INV_X1 U2269 ( .A(n211), .ZN(n70) );
  OAI22_X1 U2270 ( .A1(n5682), .A2(n322), .B1(n5683), .B2(n323), .ZN(n211) );
  OAI221_X1 U2271 ( .B1(n67), .B2(n6554), .C1(\Mpath/the_alu/N27 ), .C2(
        net55856), .A(n1617), .ZN(n4457) );
  AOI22_X1 U2272 ( .A1(n6556), .A2(n206), .B1(n6560), .B2(n1618), .ZN(n1617)
         );
  OAI221_X1 U2274 ( .B1(n5822), .B2(n320), .C1(n5745), .C2(n5560), .A(n321), 
        .ZN(n207) );
  OAI22_X1 U2275 ( .A1(n5560), .A2(net55844), .B1(n66), .B2(net55908), .ZN(
        n4458) );
  INV_X1 U2276 ( .A(n206), .ZN(n66) );
  OAI22_X1 U2277 ( .A1(n5674), .A2(n322), .B1(n5675), .B2(n323), .ZN(n206) );
  OAI221_X1 U2278 ( .B1(n63), .B2(n6554), .C1(\Mpath/the_alu/N25 ), .C2(
        net55852), .A(n1619), .ZN(n4459) );
  AOI22_X1 U2279 ( .A1(n6556), .A2(n201), .B1(n6560), .B2(n1620), .ZN(n1619)
         );
  OAI221_X1 U2281 ( .B1(n5812), .B2(n320), .C1(n5745), .C2(n5557), .A(n321), 
        .ZN(n202) );
  OAI22_X1 U2282 ( .A1(n5557), .A2(net55844), .B1(n62), .B2(net55908), .ZN(
        n4460) );
  INV_X1 U2283 ( .A(n201), .ZN(n62) );
  OAI22_X1 U2284 ( .A1(n5666), .A2(n322), .B1(n5667), .B2(n323), .ZN(n201) );
  OAI221_X1 U2285 ( .B1(n59), .B2(n6554), .C1(\Mpath/the_alu/N23 ), .C2(
        net55852), .A(n1621), .ZN(n4461) );
  AOI22_X1 U2286 ( .A1(n6556), .A2(n193), .B1(n6560), .B2(n1622), .ZN(n1621)
         );
  OAI221_X1 U2288 ( .B1(n5800), .B2(n320), .C1(n5745), .C2(n5551), .A(n321), 
        .ZN(n196) );
  OAI22_X1 U2289 ( .A1(n5551), .A2(net55844), .B1(n58), .B2(net55910), .ZN(
        n4462) );
  INV_X1 U2290 ( .A(n193), .ZN(n58) );
  OAI22_X1 U2291 ( .A1(n5656), .A2(n322), .B1(n5658), .B2(n323), .ZN(n193) );
  OAI221_X1 U2292 ( .B1(n1623), .B2(n214), .C1(\Mpath/the_alu/N38 ), .C2(
        net55854), .A(n1624), .ZN(n4463) );
  AOI222_X1 U2293 ( .A1(n197), .A2(n89), .B1(n192), .B2(n1080), .C1(n195), 
        .C2(n1404), .ZN(n1624) );
  OAI221_X1 U2294 ( .B1(n320), .B2(n1625), .C1(n5745), .C2(n5575), .A(n321), 
        .ZN(n1404) );
  INV_X1 U2295 ( .A(n6544), .ZN(n1625) );
  OAI22_X1 U2296 ( .A1(n5575), .A2(net55842), .B1(n86), .B2(net55910), .ZN(
        n4464) );
  INV_X1 U2297 ( .A(n1080), .ZN(n86) );
  OAI222_X1 U2298 ( .A1(n1626), .A2(n323), .B1(n6223), .B2(n402), .C1(n1627), 
        .C2(n322), .ZN(n1080) );
  INV_X1 U2299 ( .A(n6226), .ZN(n1627) );
  INV_X1 U2300 ( .A(n6225), .ZN(n1626) );
  OAI22_X1 U2301 ( .A1(net55880), .A2(n1628), .B1(n6223), .B2(net55838), .ZN(
        n4465) );
  INV_X1 U2302 ( .A(jar_in[23]), .ZN(n1628) );
  OAI22_X1 U2303 ( .A1(net55880), .A2(n1629), .B1(n6235), .B2(net55840), .ZN(
        n4466) );
  INV_X1 U2304 ( .A(jar_in[22]), .ZN(n1629) );
  OAI22_X1 U2305 ( .A1(net55880), .A2(n1630), .B1(n6247), .B2(net55840), .ZN(
        n4467) );
  INV_X1 U2306 ( .A(jar_in[21]), .ZN(n1630) );
  OAI22_X1 U2307 ( .A1(net55880), .A2(n1631), .B1(n6263), .B2(net55838), .ZN(
        n4468) );
  INV_X1 U2308 ( .A(jar_in[20]), .ZN(n1631) );
  OAI22_X1 U2309 ( .A1(net55880), .A2(n1632), .B1(n6276), .B2(net55838), .ZN(
        n4469) );
  INV_X1 U2310 ( .A(jar_in[19]), .ZN(n1632) );
  OAI22_X1 U2311 ( .A1(net55880), .A2(n1633), .B1(n6291), .B2(net55838), .ZN(
        n4470) );
  INV_X1 U2312 ( .A(jar_in[18]), .ZN(n1633) );
  OAI22_X1 U2313 ( .A1(net55882), .A2(n1634), .B1(n6305), .B2(net55838), .ZN(
        n4471) );
  INV_X1 U2314 ( .A(jar_in[17]), .ZN(n1634) );
  OAI22_X1 U2315 ( .A1(net55882), .A2(n1635), .B1(n6317), .B2(net55838), .ZN(
        n4472) );
  INV_X1 U2316 ( .A(jar_in[16]), .ZN(n1635) );
  OAI22_X1 U2317 ( .A1(net55882), .A2(n1636), .B1(n6329), .B2(net55836), .ZN(
        n4473) );
  INV_X1 U2318 ( .A(jar_in[15]), .ZN(n1636) );
  OAI22_X1 U2319 ( .A1(net55882), .A2(n1637), .B1(n6341), .B2(net55836), .ZN(
        n4474) );
  INV_X1 U2320 ( .A(jar_in[14]), .ZN(n1637) );
  OAI22_X1 U2321 ( .A1(net55882), .A2(n1638), .B1(n6353), .B2(net55836), .ZN(
        n4475) );
  INV_X1 U2322 ( .A(jar_in[13]), .ZN(n1638) );
  OAI22_X1 U2323 ( .A1(net55882), .A2(n1639), .B1(n6365), .B2(net55838), .ZN(
        n4476) );
  INV_X1 U2324 ( .A(jar_in[12]), .ZN(n1639) );
  OAI22_X1 U2325 ( .A1(net55882), .A2(n1640), .B1(n6377), .B2(net55838), .ZN(
        n4477) );
  INV_X1 U2326 ( .A(jar_in[11]), .ZN(n1640) );
  OAI22_X1 U2327 ( .A1(net55884), .A2(n1641), .B1(n6391), .B2(net55838), .ZN(
        n4478) );
  INV_X1 U2328 ( .A(jar_in[10]), .ZN(n1641) );
  OAI22_X1 U2329 ( .A1(net55884), .A2(n1642), .B1(n6114), .B2(net55836), .ZN(
        n4479) );
  INV_X1 U2330 ( .A(jar_in[9]), .ZN(n1642) );
  OAI22_X1 U2331 ( .A1(net55884), .A2(n1643), .B1(n6127), .B2(net55838), .ZN(
        n4480) );
  INV_X1 U2332 ( .A(jar_in[8]), .ZN(n1643) );
  OAI22_X1 U2333 ( .A1(net55884), .A2(n1644), .B1(n6139), .B2(net55838), .ZN(
        n4481) );
  INV_X1 U2334 ( .A(jar_in[7]), .ZN(n1644) );
  OAI22_X1 U2335 ( .A1(net55884), .A2(n1645), .B1(n6151), .B2(net55836), .ZN(
        n4482) );
  INV_X1 U2336 ( .A(jar_in[6]), .ZN(n1645) );
  OAI22_X1 U2337 ( .A1(net55884), .A2(n1646), .B1(n6163), .B2(net55836), .ZN(
        n4483) );
  INV_X1 U2338 ( .A(jar_in[5]), .ZN(n1646) );
  OAI22_X1 U2339 ( .A1(net55884), .A2(n1647), .B1(n6180), .B2(net55838), .ZN(
        n4484) );
  INV_X1 U2340 ( .A(jar_in[4]), .ZN(n1647) );
  OAI22_X1 U2341 ( .A1(net55886), .A2(n1648), .B1(n6194), .B2(net55836), .ZN(
        n4485) );
  INV_X1 U2342 ( .A(jar_in[3]), .ZN(n1648) );
  OAI22_X1 U2343 ( .A1(net55886), .A2(n1649), .B1(n6209), .B2(net55836), .ZN(
        n4486) );
  INV_X1 U2344 ( .A(jar_in[2]), .ZN(n1649) );
  OAI22_X1 U2345 ( .A1(net55886), .A2(n1650), .B1(n6087), .B2(net55836), .ZN(
        n4487) );
  INV_X1 U2346 ( .A(jar_in[1]), .ZN(n1650) );
  OAI22_X1 U2347 ( .A1(net55888), .A2(n1651), .B1(net55832), .B2(n1652), .ZN(
        n4488) );
  INV_X1 U2348 ( .A(jar_in[0]), .ZN(n1651) );
  INV_X1 U2351 ( .A(n1654), .ZN(n4490) );
  AOI221_X1 U2352 ( .B1(n371), .B2(\Mcontrol/f_currpc[10] ), .C1(n372), .C2(
        n7881), .A(n373), .ZN(n1654) );
  INV_X1 U2353 ( .A(n6547), .ZN(n373) );
  OAI22_X1 U2357 ( .A1(n6489), .A2(n7110), .B1(serve_exception), .B2(n49), 
        .ZN(n4491) );
  AOI22_X1 U2358 ( .A1(\Scc_coproc/x_exc_word[0] ), .A2(n883), .B1(n1656), 
        .B2(\Scc_coproc/N551 ), .ZN(n49) );
  NAND2_X1 U2359 ( .A1(n1590), .A2(n1657), .ZN(n1656) );
  OAI21_X1 U2360 ( .B1(\Scc_coproc/interrupt[7] ), .B2(n6490), .A(n1591), .ZN(
        n1657) );
  OAI221_X1 U2361 ( .B1(n5547), .B2(n1658), .C1(\Mpath/the_alu/N22 ), .C2(
        net55856), .A(n1659), .ZN(n4492) );
  AOI21_X1 U2362 ( .B1(n195), .B2(n1390), .A(n1660), .ZN(n1659) );
  OAI22_X1 U2363 ( .A1(n50), .A2(n1661), .B1(n1662), .B2(n214), .ZN(n1660) );
  AOI21_X1 U2364 ( .B1(n5845), .B2(n215), .A(n1663), .ZN(n1662) );
  OAI221_X1 U2365 ( .B1(n5791), .B2(n320), .C1(n5745), .C2(n5548), .A(n321), 
        .ZN(n1390) );
  AND2_X1 U2366 ( .A1(n654), .A2(n1664), .ZN(n321) );
  NAND2_X1 U2367 ( .A1(n5962), .A2(n5745), .ZN(n1664) );
  NAND2_X1 U2368 ( .A1(n5748), .A2(n5745), .ZN(n654) );
  NAND3_X1 U2369 ( .A1(n5967), .A2(n5745), .A3(n5968), .ZN(n320) );
  OAI22_X1 U2370 ( .A1(n5548), .A2(net55846), .B1(n50), .B2(net55910), .ZN(
        n4493) );
  INV_X1 U2371 ( .A(n1085), .ZN(n50) );
  OAI22_X1 U2372 ( .A1(n6436), .A2(n322), .B1(n6437), .B2(n323), .ZN(n1085) );
  OAI221_X1 U2373 ( .B1(n179), .B2(n6554), .C1(\Mpath/the_alu/N83 ), .C2(
        net55858), .A(n1665), .ZN(n4494) );
  AOI22_X1 U2374 ( .A1(n6556), .A2(n1666), .B1(n6560), .B2(n1667), .ZN(n1665)
         );
  NOR3_X1 U2375 ( .A1(\regfile/N264 ), .A2(byp_controlA[2]), .A3(net55910), 
        .ZN(n235) );
  NOR2_X1 U2376 ( .A1(rs1_addr[0]), .A2(\regfile/N262 ), .ZN(\regfile/N264 )
         );
  NAND3_X1 U2378 ( .A1(net55840), .A2(n7324), .A3(byp_controlA[2]), .ZN(n232)
         );
  OAI22_X1 U2380 ( .A1(n5620), .A2(net55844), .B1(n178), .B2(net55910), .ZN(
        n4495) );
  INV_X1 U2381 ( .A(n1666), .ZN(n178) );
  OAI22_X1 U2382 ( .A1(n5714), .A2(net55916), .B1(\Mpath/the_memhandle/N240 ), 
        .B2(net55836), .ZN(n4496) );
  OAI211_X1 U2383 ( .C1(\Mpath/the_alu/N84 ), .C2(net55862), .A(n1669), .B(
        n1670), .ZN(n4497) );
  AOI221_X1 U2384 ( .B1(n195), .B2(n1668), .C1(n192), .C2(n1666), .A(n1671), 
        .ZN(n1670) );
  NOR4_X1 U2385 ( .A1(n1672), .A2(net55888), .A3(n1517), .A4(n1518), .ZN(n1671) );
  INV_X1 U2386 ( .A(n1673), .ZN(n1517) );
  OAI222_X1 U2387 ( .A1(n5714), .A2(n323), .B1(n402), .B2(n1652), .C1(n5715), 
        .C2(n322), .ZN(n1666) );
  NAND2_X1 U2389 ( .A1(n322), .A2(n1674), .ZN(n402) );
  INV_X1 U2390 ( .A(\Mpath/N197 ), .ZN(n1674) );
  NAND3_X1 U2393 ( .A1(exe_outsel[1]), .A2(exe_outsel[0]), .A3(exe_outsel[2]), 
        .ZN(n1675) );
  NAND2_X1 U2395 ( .A1(n1676), .A2(n185), .ZN(n1661) );
  NOR2_X1 U2396 ( .A1(n1677), .A2(byp_controlB[0]), .ZN(n185) );
  OAI222_X1 U2397 ( .A1(n1678), .A2(n995), .B1(n1679), .B2(n1398), .C1(n5745), 
        .C2(n5620), .ZN(n1668) );
  NAND2_X1 U2398 ( .A1(\Mpath/the_memhandle/N34 ), .A2(n5745), .ZN(n1398) );
  AOI221_X1 U2399 ( .B1(n6538), .B2(n1571), .C1(n6527), .C2(n1572), .A(n6014), 
        .ZN(n1679) );
  INV_X1 U2400 ( .A(n6000), .ZN(n1572) );
  INV_X1 U2401 ( .A(n5804), .ZN(n1571) );
  NAND2_X1 U2402 ( .A1(n5745), .A2(n1396), .ZN(n995) );
  INV_X1 U2403 ( .A(\Mpath/the_memhandle/N34 ), .ZN(n1396) );
  AOI221_X1 U2404 ( .B1(n5786), .B2(n1564), .C1(n5787), .C2(n6534), .A(n6010), 
        .ZN(n1678) );
  INV_X1 U2405 ( .A(n6015), .ZN(n1564) );
  NOR2_X1 U2407 ( .A1(n1677), .A2(\Mcontrol/st_logic/N42 ), .ZN(n184) );
  INV_X1 U2408 ( .A(byp_controlB[2]), .ZN(n1677) );
  AOI22_X1 U2409 ( .A1(n197), .A2(n181), .B1(n329), .B2(net56595), .ZN(n1669)
         );
  INV_X1 U2410 ( .A(n214), .ZN(n329) );
  NAND2_X1 U2411 ( .A1(n1672), .A2(net55824), .ZN(n214) );
  NAND2_X1 U2413 ( .A1(n1676), .A2(n182), .ZN(n1658) );
  NOR2_X1 U2414 ( .A1(byp_controlB[2]), .A2(\regfile/N269 ), .ZN(n182) );
  NOR2_X1 U2415 ( .A1(rs2_addr[0]), .A2(\regfile/N267 ), .ZN(\regfile/N269 )
         );
  AOI21_X1 U2417 ( .B1(n1680), .B2(n6960), .A(net57323), .ZN(n1672) );
  OAI21_X1 U2418 ( .B1(n1681), .B2(\Mcontrol/Operation_decoding32/N2037 ), .A(
        n7225), .ZN(n1680) );
  INV_X1 U2419 ( .A(n6510), .ZN(n1681) );
  OAI22_X1 U2420 ( .A1(n1573), .A2(net55916), .B1(net55832), .B2(
        \Mpath/the_memhandle/N239 ), .ZN(n4498) );
  INV_X1 U2421 ( .A(daddr_out[1]), .ZN(n1573) );
  OAI22_X1 U2422 ( .A1(net55886), .A2(n1682), .B1(net55834), .B2(n3102), .ZN(
        n4499) );
  OAI22_X1 U2423 ( .A1(net55886), .A2(n1683), .B1(net55832), .B2(n3103), .ZN(
        n4500) );
  OAI22_X1 U2424 ( .A1(n3107), .A2(net55914), .B1(net55832), .B2(n3104), .ZN(
        n4501) );
  NOR2_X1 U2425 ( .A1(net55822), .A2(n1682), .ZN(n4502) );
  NOR2_X1 U2427 ( .A1(net55822), .A2(n1683), .ZN(n4503) );
  NOR2_X1 U2429 ( .A1(n3107), .A2(net55834), .ZN(n4504) );
  NOR3_X1 U2435 ( .A1(n7187), .A2(n1690), .A3(n1688), .ZN(n1691) );
  INV_X1 U2436 ( .A(\Mpath/the_alu/N22 ), .ZN(n1690) );
  OAI21_X1 U2437 ( .B1(\Mpath/the_alu/N21 ), .B2(n1693), .A(n1694), .ZN(n1689)
         );
  INV_X1 U2438 ( .A(\Mpath/the_alu/N21 ), .ZN(n1688) );
  INV_X1 U2439 ( .A(n1695), .ZN(n1687) );
  XOR2_X1 U2441 ( .A(\Mpath/the_alu/N21 ), .B(\Mpath/the_alu/N22 ), .Z(n6512)
         );
  AND2_X1 U2442 ( .A1(n1699), .A2(n1700), .ZN(n6436) );
  AOI222_X1 U2443 ( .A1(\Mpath/the_shift/sh_rol [31]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [31]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [31]), .C2(n1703), .ZN(n1700) );
  AOI22_X1 U2444 ( .A1(\Mpath/the_shift/sh_sra [31]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [31]), .B2(\Mpath/the_shift/N118 ), .ZN(n1699)
         );
  NAND2_X1 U2445 ( .A1(n1705), .A2(n1706), .ZN(n6395) );
  AOI222_X1 U2446 ( .A1(\Mpath/the_shift/sh_rol [10]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [10]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [10]), .C2(n1703), .ZN(n1706) );
  AOI22_X1 U2447 ( .A1(\Mpath/the_shift/sh_sra [10]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [10]), .B2(\Mpath/the_shift/N118 ), .ZN(n1705)
         );
  NAND3_X1 U2448 ( .A1(n1707), .A2(n1708), .A3(n1709), .ZN(n6394) );
  AOI222_X1 U2449 ( .A1(\Mpath/the_alu/sum[10] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[10] ), .B2(n1698), .C1(n7293), .C2(n1711), .ZN(
        n1709) );
  INV_X1 U2450 ( .A(\Mpath/the_alu/N63 ), .ZN(n1711) );
  AOI22_X1 U2451 ( .A1(\Mpath/the_alu/N115 ), .A2(n1712), .B1(
        \Mpath/the_alu/N179 ), .B2(n1697), .ZN(n1708) );
  AOI22_X1 U2452 ( .A1(\Mpath/the_alu/N211 ), .A2(n1713), .B1(
        \Mpath/the_alu/N147 ), .B2(n1714), .ZN(n1707) );
  NAND2_X1 U2454 ( .A1(n1715), .A2(n1716), .ZN(n6381) );
  AOI222_X1 U2455 ( .A1(\Mpath/the_shift/sh_rol [11]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [11]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [11]), .C2(n1703), .ZN(n1716) );
  AOI22_X1 U2456 ( .A1(\Mpath/the_shift/sh_sra [11]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [11]), .B2(\Mpath/the_shift/N118 ), .ZN(n1715)
         );
  NAND3_X1 U2457 ( .A1(n1717), .A2(n1718), .A3(n1719), .ZN(n6380) );
  AOI222_X1 U2458 ( .A1(\Mpath/the_alu/sum[11] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[11] ), .B2(n1698), .C1(n7293), .C2(n1720), .ZN(
        n1719) );
  INV_X1 U2459 ( .A(\Mpath/the_alu/N61 ), .ZN(n1720) );
  AOI22_X1 U2460 ( .A1(\Mpath/the_alu/N114 ), .A2(n1712), .B1(
        \Mpath/the_alu/N178 ), .B2(n1697), .ZN(n1718) );
  AOI22_X1 U2461 ( .A1(\Mpath/the_alu/N210 ), .A2(n1713), .B1(
        \Mpath/the_alu/N146 ), .B2(n1714), .ZN(n1717) );
  NAND2_X1 U2462 ( .A1(n1721), .A2(n1722), .ZN(n6369) );
  AOI222_X1 U2463 ( .A1(\Mpath/the_shift/sh_rol [12]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [12]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [12]), .C2(n1703), .ZN(n1722) );
  AOI22_X1 U2464 ( .A1(\Mpath/the_shift/sh_sra [12]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [12]), .B2(\Mpath/the_shift/N118 ), .ZN(n1721)
         );
  NAND3_X1 U2465 ( .A1(n1723), .A2(n1724), .A3(n1725), .ZN(n6368) );
  AOI222_X1 U2466 ( .A1(\Mpath/the_alu/sum[12] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[12] ), .B2(n1698), .C1(n7293), .C2(n1726), .ZN(
        n1725) );
  INV_X1 U2467 ( .A(\Mpath/the_alu/N59 ), .ZN(n1726) );
  AOI22_X1 U2468 ( .A1(\Mpath/the_alu/N113 ), .A2(n1712), .B1(
        \Mpath/the_alu/N177 ), .B2(n1697), .ZN(n1724) );
  AOI22_X1 U2469 ( .A1(\Mpath/the_alu/N209 ), .A2(n1713), .B1(
        \Mpath/the_alu/N145 ), .B2(n1714), .ZN(n1723) );
  NAND2_X1 U2470 ( .A1(n1727), .A2(n1728), .ZN(n6357) );
  AOI222_X1 U2471 ( .A1(\Mpath/the_shift/sh_rol [13]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [13]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [13]), .C2(n1703), .ZN(n1728) );
  AOI22_X1 U2472 ( .A1(\Mpath/the_shift/sh_sra [13]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [13]), .B2(\Mpath/the_shift/N118 ), .ZN(n1727)
         );
  NAND3_X1 U2473 ( .A1(n1729), .A2(n1730), .A3(n1731), .ZN(n6356) );
  AOI222_X1 U2474 ( .A1(\Mpath/the_alu/sum[13] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[13] ), .B2(n1698), .C1(n7293), .C2(n1732), .ZN(
        n1731) );
  INV_X1 U2475 ( .A(\Mpath/the_alu/N57 ), .ZN(n1732) );
  AOI22_X1 U2476 ( .A1(\Mpath/the_alu/N112 ), .A2(n1712), .B1(
        \Mpath/the_alu/N176 ), .B2(n1697), .ZN(n1730) );
  AOI22_X1 U2477 ( .A1(\Mpath/the_alu/N208 ), .A2(n1713), .B1(
        \Mpath/the_alu/N144 ), .B2(n1714), .ZN(n1729) );
  AOI222_X1 U2479 ( .A1(\Mpath/the_shift/sh_rol [14]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [14]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [14]), .C2(n1703), .ZN(n1734) );
  AOI22_X1 U2480 ( .A1(\Mpath/the_shift/sh_sra [14]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [14]), .B2(\Mpath/the_shift/N118 ), .ZN(n1733)
         );
  NAND3_X1 U2481 ( .A1(n1735), .A2(n1736), .A3(n1737), .ZN(n6344) );
  AOI222_X1 U2482 ( .A1(\Mpath/the_alu/sum[14] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[14] ), .B2(n1698), .C1(n7293), .C2(n1738), .ZN(
        n1737) );
  INV_X1 U2483 ( .A(\Mpath/the_alu/N55 ), .ZN(n1738) );
  AOI22_X1 U2484 ( .A1(\Mpath/the_alu/N111 ), .A2(n1712), .B1(
        \Mpath/the_alu/N175 ), .B2(n1697), .ZN(n1736) );
  AOI22_X1 U2485 ( .A1(\Mpath/the_alu/N207 ), .A2(n1713), .B1(
        \Mpath/the_alu/N143 ), .B2(n1714), .ZN(n1735) );
  NAND2_X1 U2486 ( .A1(n1739), .A2(n1740), .ZN(n6333) );
  AOI222_X1 U2487 ( .A1(\Mpath/the_shift/sh_rol [15]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [15]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [15]), .C2(n1703), .ZN(n1740) );
  AOI22_X1 U2488 ( .A1(\Mpath/the_shift/sh_sra [15]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [15]), .B2(\Mpath/the_shift/N118 ), .ZN(n1739)
         );
  NAND3_X1 U2489 ( .A1(n1741), .A2(n1742), .A3(n1743), .ZN(n6332) );
  AOI222_X1 U2490 ( .A1(\Mpath/the_alu/sum[15] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[15] ), .B2(n1698), .C1(n7293), .C2(n1744), .ZN(
        n1743) );
  INV_X1 U2491 ( .A(\Mpath/the_alu/N53 ), .ZN(n1744) );
  AOI22_X1 U2492 ( .A1(\Mpath/the_alu/N110 ), .A2(n1712), .B1(
        \Mpath/the_alu/N174 ), .B2(n1697), .ZN(n1742) );
  AOI22_X1 U2493 ( .A1(\Mpath/the_alu/N206 ), .A2(n1713), .B1(
        \Mpath/the_alu/N142 ), .B2(n1714), .ZN(n1741) );
  NAND3_X1 U2494 ( .A1(n1474), .A2(n7598), .A3(n7436), .ZN(n6321) );
  NAND2_X1 U2495 ( .A1(n1745), .A2(n1746), .ZN(n6320) );
  AOI222_X1 U2496 ( .A1(\Mpath/the_shift/sh_rol [16]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [16]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [16]), .C2(n1703), .ZN(n1746) );
  AOI22_X1 U2497 ( .A1(\Mpath/the_shift/sh_sra [16]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [16]), .B2(\Mpath/the_shift/N118 ), .ZN(n1745)
         );
  NAND3_X1 U2498 ( .A1(n1747), .A2(n1748), .A3(n1749), .ZN(n6319) );
  AOI222_X1 U2499 ( .A1(\Mpath/the_alu/sum[16] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[16] ), .B2(n1698), .C1(n7293), .C2(n1750), .ZN(
        n1749) );
  INV_X1 U2500 ( .A(\Mpath/the_alu/N51 ), .ZN(n1750) );
  AOI22_X1 U2501 ( .A1(\Mpath/the_alu/N109 ), .A2(n1712), .B1(
        \Mpath/the_alu/N173 ), .B2(n1697), .ZN(n1748) );
  AOI22_X1 U2502 ( .A1(\Mpath/the_alu/N205 ), .A2(n1713), .B1(
        \Mpath/the_alu/N141 ), .B2(n1714), .ZN(n1747) );
  NAND2_X1 U2503 ( .A1(n1751), .A2(n1752), .ZN(n6308) );
  AOI222_X1 U2504 ( .A1(\Mpath/the_shift/sh_rol [17]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [17]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [17]), .C2(n1703), .ZN(n1752) );
  AOI22_X1 U2505 ( .A1(\Mpath/the_shift/sh_sra [17]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [17]), .B2(\Mpath/the_shift/N118 ), .ZN(n1751)
         );
  NAND3_X1 U2506 ( .A1(n1753), .A2(n1754), .A3(n1755), .ZN(n6307) );
  AOI222_X1 U2507 ( .A1(\Mpath/the_alu/sum[17] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[17] ), .B2(n1698), .C1(n7293), .C2(n1756), .ZN(
        n1755) );
  INV_X1 U2508 ( .A(\Mpath/the_alu/N49 ), .ZN(n1756) );
  AOI22_X1 U2509 ( .A1(\Mpath/the_alu/N108 ), .A2(n1712), .B1(
        \Mpath/the_alu/N172 ), .B2(n1697), .ZN(n1754) );
  AOI22_X1 U2510 ( .A1(\Mpath/the_alu/N204 ), .A2(n1713), .B1(
        \Mpath/the_alu/N140 ), .B2(n1714), .ZN(n1753) );
  NAND2_X1 U2511 ( .A1(n1757), .A2(n1758), .ZN(n6294) );
  AOI222_X1 U2512 ( .A1(\Mpath/the_shift/sh_rol [18]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [18]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [18]), .C2(n1703), .ZN(n1758) );
  AOI22_X1 U2513 ( .A1(\Mpath/the_shift/sh_sra [18]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [18]), .B2(\Mpath/the_shift/N118 ), .ZN(n1757)
         );
  NAND3_X1 U2514 ( .A1(n1759), .A2(n1760), .A3(n1761), .ZN(n6293) );
  AOI222_X1 U2515 ( .A1(\Mpath/the_alu/sum[18] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[18] ), .B2(n1698), .C1(n7293), .C2(n1762), .ZN(
        n1761) );
  INV_X1 U2516 ( .A(\Mpath/the_alu/N47 ), .ZN(n1762) );
  AOI22_X1 U2517 ( .A1(\Mpath/the_alu/N107 ), .A2(n1712), .B1(
        \Mpath/the_alu/N171 ), .B2(n1697), .ZN(n1760) );
  AOI22_X1 U2518 ( .A1(\Mpath/the_alu/N203 ), .A2(n1713), .B1(
        \Mpath/the_alu/N139 ), .B2(n1714), .ZN(n1759) );
  NAND2_X1 U2519 ( .A1(n1763), .A2(n1764), .ZN(n6279) );
  AOI222_X1 U2520 ( .A1(\Mpath/the_shift/sh_rol [19]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [19]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [19]), .C2(n1703), .ZN(n1764) );
  AOI22_X1 U2521 ( .A1(\Mpath/the_shift/sh_sra [19]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [19]), .B2(\Mpath/the_shift/N118 ), .ZN(n1763)
         );
  NAND3_X1 U2522 ( .A1(n1765), .A2(n1766), .A3(n1767), .ZN(n6278) );
  AOI222_X1 U2523 ( .A1(\Mpath/the_alu/sum[19] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[19] ), .B2(n1698), .C1(n7293), .C2(n1768), .ZN(
        n1767) );
  INV_X1 U2524 ( .A(\Mpath/the_alu/N45 ), .ZN(n1768) );
  AOI22_X1 U2525 ( .A1(\Mpath/the_alu/N106 ), .A2(n1712), .B1(
        \Mpath/the_alu/N170 ), .B2(n1697), .ZN(n1766) );
  AOI22_X1 U2526 ( .A1(\Mpath/the_alu/N202 ), .A2(n1713), .B1(
        \Mpath/the_alu/N138 ), .B2(n1714), .ZN(n1765) );
  NAND2_X1 U2527 ( .A1(n1769), .A2(n1770), .ZN(n6266) );
  AOI222_X1 U2528 ( .A1(\Mpath/the_shift/sh_rol [20]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [20]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [20]), .C2(n1703), .ZN(n1770) );
  AOI22_X1 U2529 ( .A1(\Mpath/the_shift/sh_sra [20]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [20]), .B2(\Mpath/the_shift/N118 ), .ZN(n1769)
         );
  NAND3_X1 U2530 ( .A1(n1771), .A2(n1772), .A3(n1773), .ZN(n6265) );
  AOI222_X1 U2531 ( .A1(\Mpath/the_alu/sum[20] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[20] ), .B2(n1698), .C1(n7293), .C2(n1774), .ZN(
        n1773) );
  INV_X1 U2532 ( .A(\Mpath/the_alu/N43 ), .ZN(n1774) );
  AOI22_X1 U2533 ( .A1(\Mpath/the_alu/N105 ), .A2(n1712), .B1(
        \Mpath/the_alu/N169 ), .B2(n1697), .ZN(n1772) );
  AOI22_X1 U2534 ( .A1(\Mpath/the_alu/N201 ), .A2(n1713), .B1(
        \Mpath/the_alu/N137 ), .B2(n1714), .ZN(n1771) );
  NAND2_X1 U2535 ( .A1(n1775), .A2(n1776), .ZN(n6250) );
  AOI222_X1 U2536 ( .A1(\Mpath/the_shift/sh_rol [21]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [21]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [21]), .C2(n1703), .ZN(n1776) );
  AOI22_X1 U2537 ( .A1(\Mpath/the_shift/sh_sra [21]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [21]), .B2(\Mpath/the_shift/N118 ), .ZN(n1775)
         );
  NAND3_X1 U2538 ( .A1(n1777), .A2(n1778), .A3(n1779), .ZN(n6249) );
  AOI222_X1 U2539 ( .A1(\Mpath/the_alu/sum[21] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[21] ), .B2(n1698), .C1(n7293), .C2(n1780), .ZN(
        n1779) );
  INV_X1 U2540 ( .A(\Mpath/the_alu/N41 ), .ZN(n1780) );
  AOI22_X1 U2541 ( .A1(\Mpath/the_alu/N104 ), .A2(n1712), .B1(
        \Mpath/the_alu/N168 ), .B2(n1697), .ZN(n1778) );
  AOI22_X1 U2542 ( .A1(\Mpath/the_alu/N200 ), .A2(n1713), .B1(
        \Mpath/the_alu/N136 ), .B2(n1714), .ZN(n1777) );
  NAND2_X1 U2543 ( .A1(n1781), .A2(n1782), .ZN(n6238) );
  AOI222_X1 U2544 ( .A1(\Mpath/the_shift/sh_rol [22]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [22]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [22]), .C2(n1703), .ZN(n1782) );
  AOI22_X1 U2545 ( .A1(\Mpath/the_shift/sh_sra [22]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [22]), .B2(\Mpath/the_shift/N118 ), .ZN(n1781)
         );
  NAND3_X1 U2546 ( .A1(n1783), .A2(n1784), .A3(n1785), .ZN(n6237) );
  AOI222_X1 U2547 ( .A1(\Mpath/the_alu/sum[22] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[22] ), .B2(n1698), .C1(n7293), .C2(n1786), .ZN(
        n1785) );
  INV_X1 U2548 ( .A(\Mpath/the_alu/N39 ), .ZN(n1786) );
  AOI22_X1 U2549 ( .A1(\Mpath/the_alu/N103 ), .A2(n1712), .B1(
        \Mpath/the_alu/N167 ), .B2(n1697), .ZN(n1784) );
  AOI22_X1 U2550 ( .A1(\Mpath/the_alu/N199 ), .A2(n1713), .B1(
        \Mpath/the_alu/N135 ), .B2(n1714), .ZN(n1783) );
  NAND2_X1 U2551 ( .A1(n1787), .A2(n1788), .ZN(n6226) );
  AOI222_X1 U2552 ( .A1(\Mpath/the_shift/sh_rol [23]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [23]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [23]), .C2(n1703), .ZN(n1788) );
  AOI22_X1 U2553 ( .A1(\Mpath/the_shift/sh_sra [23]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [23]), .B2(\Mpath/the_shift/N118 ), .ZN(n1787)
         );
  NAND3_X1 U2554 ( .A1(n1789), .A2(n1790), .A3(n1791), .ZN(n6225) );
  AOI222_X1 U2555 ( .A1(\Mpath/the_alu/sum[23] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[23] ), .B2(n1698), .C1(n7293), .C2(n1792), .ZN(
        n1791) );
  INV_X1 U2556 ( .A(\Mpath/the_alu/N37 ), .ZN(n1792) );
  AOI22_X1 U2557 ( .A1(\Mpath/the_alu/N102 ), .A2(n1712), .B1(
        \Mpath/the_alu/N166 ), .B2(n1697), .ZN(n1790) );
  AOI22_X1 U2558 ( .A1(\Mpath/the_alu/N198 ), .A2(n1713), .B1(
        \Mpath/the_alu/N134 ), .B2(n1714), .ZN(n1789) );
  NAND2_X1 U2559 ( .A1(n1793), .A2(n1794), .ZN(n6213) );
  AOI222_X1 U2560 ( .A1(\Mpath/the_shift/sh_rol [2]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [2]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [2]), .C2(n1703), .ZN(n1794) );
  AOI22_X1 U2561 ( .A1(\Mpath/the_shift/sh_sra [2]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [2]), .B2(\Mpath/the_shift/N118 ), .ZN(n1793)
         );
  NAND3_X1 U2562 ( .A1(n1795), .A2(n1796), .A3(n1797), .ZN(n6212) );
  AOI222_X1 U2563 ( .A1(\Mpath/the_alu/sum[2] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[2] ), .B2(n1698), .C1(n7293), .C2(n1798), .ZN(
        n1797) );
  INV_X1 U2564 ( .A(\Mpath/the_alu/N79 ), .ZN(n1798) );
  AOI22_X1 U2565 ( .A1(\Mpath/the_alu/N123 ), .A2(n1712), .B1(
        \Mpath/the_alu/N187 ), .B2(n1697), .ZN(n1796) );
  AOI22_X1 U2566 ( .A1(\Mpath/the_alu/N219 ), .A2(n1713), .B1(
        \Mpath/the_alu/N155 ), .B2(n1714), .ZN(n1795) );
  NAND2_X1 U2567 ( .A1(n1799), .A2(n1800), .ZN(n6198) );
  AOI222_X1 U2568 ( .A1(\Mpath/the_shift/sh_rol [3]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [3]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [3]), .C2(n1703), .ZN(n1800) );
  AOI22_X1 U2569 ( .A1(\Mpath/the_shift/sh_sra [3]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [3]), .B2(\Mpath/the_shift/N118 ), .ZN(n1799)
         );
  NAND3_X1 U2570 ( .A1(n1801), .A2(n1802), .A3(n1803), .ZN(n6197) );
  AOI222_X1 U2571 ( .A1(\Mpath/the_alu/sum[3] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[3] ), .B2(n1698), .C1(n7293), .C2(n1804), .ZN(
        n1803) );
  INV_X1 U2572 ( .A(\Mpath/the_alu/N77 ), .ZN(n1804) );
  AOI22_X1 U2573 ( .A1(\Mpath/the_alu/N122 ), .A2(n1712), .B1(
        \Mpath/the_alu/N186 ), .B2(n1697), .ZN(n1802) );
  AOI22_X1 U2574 ( .A1(\Mpath/the_alu/N218 ), .A2(n1713), .B1(
        \Mpath/the_alu/N154 ), .B2(n1714), .ZN(n1801) );
  NAND2_X1 U2575 ( .A1(n1805), .A2(n1806), .ZN(n6184) );
  AOI222_X1 U2576 ( .A1(\Mpath/the_shift/sh_rol [4]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [4]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [4]), .C2(n1703), .ZN(n1806) );
  AOI22_X1 U2577 ( .A1(\Mpath/the_shift/sh_sra [4]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [4]), .B2(\Mpath/the_shift/N118 ), .ZN(n1805)
         );
  NAND3_X1 U2578 ( .A1(n1807), .A2(n1808), .A3(n1809), .ZN(n6183) );
  AOI222_X1 U2579 ( .A1(\Mpath/the_alu/sum[4] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[4] ), .B2(n1698), .C1(n7293), .C2(n1810), .ZN(
        n1809) );
  INV_X1 U2580 ( .A(\Mpath/the_alu/N75 ), .ZN(n1810) );
  AOI22_X1 U2581 ( .A1(\Mpath/the_alu/N121 ), .A2(n1712), .B1(
        \Mpath/the_alu/N185 ), .B2(n1697), .ZN(n1808) );
  AOI22_X1 U2582 ( .A1(\Mpath/the_alu/N217 ), .A2(n1713), .B1(
        \Mpath/the_alu/N153 ), .B2(n1714), .ZN(n1807) );
  NAND2_X1 U2583 ( .A1(n1811), .A2(n1812), .ZN(n6167) );
  AOI222_X1 U2584 ( .A1(\Mpath/the_shift/sh_rol [5]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [5]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [5]), .C2(n1703), .ZN(n1812) );
  AOI22_X1 U2585 ( .A1(\Mpath/the_shift/sh_sra [5]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [5]), .B2(\Mpath/the_shift/N118 ), .ZN(n1811)
         );
  NAND3_X1 U2586 ( .A1(n1813), .A2(n1814), .A3(n1815), .ZN(n6166) );
  AOI222_X1 U2587 ( .A1(\Mpath/the_alu/sum[5] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[5] ), .B2(n1698), .C1(n7293), .C2(n1816), .ZN(
        n1815) );
  INV_X1 U2588 ( .A(\Mpath/the_alu/N73 ), .ZN(n1816) );
  AOI22_X1 U2589 ( .A1(\Mpath/the_alu/N120 ), .A2(n1712), .B1(
        \Mpath/the_alu/N184 ), .B2(n1697), .ZN(n1814) );
  AOI22_X1 U2590 ( .A1(\Mpath/the_alu/N216 ), .A2(n1713), .B1(
        \Mpath/the_alu/N152 ), .B2(n1714), .ZN(n1813) );
  AOI222_X1 U2592 ( .A1(\Mpath/the_shift/sh_rol [6]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [6]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [6]), .C2(n1703), .ZN(n1818) );
  AOI22_X1 U2593 ( .A1(\Mpath/the_shift/sh_sra [6]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [6]), .B2(\Mpath/the_shift/N118 ), .ZN(n1817)
         );
  NAND3_X1 U2594 ( .A1(n1819), .A2(n1820), .A3(n1821), .ZN(n6154) );
  AOI222_X1 U2595 ( .A1(\Mpath/the_alu/sum[6] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[6] ), .B2(n1698), .C1(n7293), .C2(n1822), .ZN(
        n1821) );
  INV_X1 U2596 ( .A(\Mpath/the_alu/N71 ), .ZN(n1822) );
  AOI22_X1 U2597 ( .A1(\Mpath/the_alu/N119 ), .A2(n1712), .B1(
        \Mpath/the_alu/N183 ), .B2(n1697), .ZN(n1820) );
  AOI22_X1 U2598 ( .A1(\Mpath/the_alu/N215 ), .A2(n1713), .B1(
        \Mpath/the_alu/N151 ), .B2(n1714), .ZN(n1819) );
  NAND2_X1 U2599 ( .A1(n1823), .A2(n1824), .ZN(n6143) );
  AOI222_X1 U2600 ( .A1(\Mpath/the_shift/sh_rol [7]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [7]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [7]), .C2(n1703), .ZN(n1824) );
  AOI22_X1 U2601 ( .A1(\Mpath/the_shift/sh_sra [7]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [7]), .B2(\Mpath/the_shift/N118 ), .ZN(n1823)
         );
  NAND3_X1 U2602 ( .A1(n1825), .A2(n1826), .A3(n1827), .ZN(n6142) );
  AOI222_X1 U2603 ( .A1(\Mpath/the_alu/sum[7] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[7] ), .B2(n1698), .C1(n7293), .C2(n1828), .ZN(
        n1827) );
  INV_X1 U2604 ( .A(\Mpath/the_alu/N69 ), .ZN(n1828) );
  AOI22_X1 U2605 ( .A1(\Mpath/the_alu/N118 ), .A2(n1712), .B1(
        \Mpath/the_alu/N182 ), .B2(n1697), .ZN(n1826) );
  AOI22_X1 U2606 ( .A1(\Mpath/the_alu/N214 ), .A2(n1713), .B1(
        \Mpath/the_alu/N150 ), .B2(n1714), .ZN(n1825) );
  NAND2_X1 U2607 ( .A1(n1829), .A2(n1830), .ZN(n6131) );
  AOI222_X1 U2608 ( .A1(\Mpath/the_shift/sh_rol [8]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [8]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [8]), .C2(n1703), .ZN(n1830) );
  AOI22_X1 U2609 ( .A1(\Mpath/the_shift/sh_sra [8]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [8]), .B2(\Mpath/the_shift/N118 ), .ZN(n1829)
         );
  NAND3_X1 U2610 ( .A1(n1831), .A2(n1832), .A3(n1833), .ZN(n6130) );
  AOI222_X1 U2611 ( .A1(\Mpath/the_alu/sum[8] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[8] ), .B2(n1698), .C1(n7293), .C2(n1834), .ZN(
        n1833) );
  AOI22_X1 U2613 ( .A1(\Mpath/the_alu/N117 ), .A2(n1712), .B1(
        \Mpath/the_alu/N181 ), .B2(n1697), .ZN(n1832) );
  AOI22_X1 U2614 ( .A1(\Mpath/the_alu/N213 ), .A2(n1713), .B1(
        \Mpath/the_alu/N149 ), .B2(n1714), .ZN(n1831) );
  NAND2_X1 U2615 ( .A1(n1835), .A2(n1836), .ZN(n6118) );
  AOI222_X1 U2616 ( .A1(\Mpath/the_shift/sh_rol [9]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [9]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [9]), .C2(n1703), .ZN(n1836) );
  AOI22_X1 U2617 ( .A1(\Mpath/the_shift/sh_sra [9]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [9]), .B2(\Mpath/the_shift/N118 ), .ZN(n1835)
         );
  NAND3_X1 U2618 ( .A1(n1837), .A2(n1838), .A3(n1839), .ZN(n6117) );
  AOI222_X1 U2619 ( .A1(\Mpath/the_alu/sum[9] ), .A2(n7634), .B1(
        \Mpath/the_alu/diff[9] ), .B2(n1698), .C1(n7293), .C2(n1840), .ZN(
        n1839) );
  INV_X1 U2620 ( .A(\Mpath/the_alu/N65 ), .ZN(n1840) );
  AOI22_X1 U2621 ( .A1(\Mpath/the_alu/N116 ), .A2(n1712), .B1(
        \Mpath/the_alu/N180 ), .B2(n1697), .ZN(n1838) );
  INV_X1 U2623 ( .A(n1693), .ZN(n1712) );
  AOI22_X1 U2624 ( .A1(\Mpath/the_alu/N212 ), .A2(n1713), .B1(
        \Mpath/the_alu/N148 ), .B2(n1714), .ZN(n1837) );
  NAND2_X1 U2626 ( .A1(n1842), .A2(n1843), .ZN(n6092) );
  AOI222_X1 U2627 ( .A1(\Mpath/the_shift/sh_rol [1]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [1]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [1]), .C2(n1703), .ZN(n1843) );
  AOI22_X1 U2628 ( .A1(\Mpath/the_shift/sh_sra [1]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [1]), .B2(\Mpath/the_shift/N118 ), .ZN(n1842)
         );
  INV_X1 U2629 ( .A(n1518), .ZN(n6077) );
  NAND2_X1 U2630 ( .A1(n1441), .A2(net56319), .ZN(n1518) );
  NOR2_X1 U2631 ( .A1(n7571), .A2(n7534), .ZN(n1441) );
  NAND3_X1 U2632 ( .A1(\Mcontrol/Operation_decoding32/N1975 ), .A2(n7434), 
        .A3(n7436), .ZN(n6075) );
  OAI21_X1 U2639 ( .B1(net56922), .B2(n7059), .A(n1851), .ZN(n1849) );
  NAND3_X1 U2640 ( .A1(\Mcontrol/Operation_decoding32/N2017 ), .A2(
        \Mcontrol/Operation_decoding32/N1922 ), .A3(
        \Mcontrol/Operation_decoding32/N2005 ), .ZN(n1851) );
  NAND2_X1 U2646 ( .A1(\Mcontrol/d_sampled_finstr [21]), .A2(n7278), .ZN(n6052) );
  INV_X1 U2647 ( .A(n5846), .ZN(n6045) );
  INV_X1 U2648 ( .A(n6538), .ZN(n6011) );
  INV_X1 U2649 ( .A(n6540), .ZN(n6001) );
  INV_X1 U2650 ( .A(n6534), .ZN(n5961) );
  INV_X1 U2651 ( .A(n6532), .ZN(n5940) );
  INV_X1 U2652 ( .A(n6542), .ZN(n5939) );
  INV_X1 U2653 ( .A(n6536), .ZN(n5936) );
  NAND2_X1 U2654 ( .A1(\Mcontrol/d_sampled_finstr [22]), .A2(n7207), .ZN(n5913) );
  INV_X1 U2655 ( .A(n6527), .ZN(n5905) );
  NAND2_X1 U2656 ( .A1(\Mcontrol/d_sampled_finstr [23]), .A2(n7207), .ZN(n5903) );
  INV_X1 U2657 ( .A(n6529), .ZN(n5895) );
  NAND2_X1 U2658 ( .A1(\Mcontrol/d_sampled_finstr [24]), .A2(n7207), .ZN(n5892) );
  NAND2_X1 U2659 ( .A1(\Mcontrol/d_sampled_finstr [25]), .A2(n7207), .ZN(n5883) );
  INV_X1 U2660 ( .A(n6530), .ZN(n5859) );
  INV_X1 U2661 ( .A(n6531), .ZN(n5857) );
  INV_X1 U2662 ( .A(D_DATA_INBUS[10]), .ZN(n5856) );
  INV_X1 U2663 ( .A(n6528), .ZN(n5834) );
  INV_X1 U2664 ( .A(n6533), .ZN(n5832) );
  INV_X1 U2665 ( .A(D_DATA_INBUS[11]), .ZN(n5831) );
  INV_X1 U2666 ( .A(n6526), .ZN(n5824) );
  INV_X1 U2667 ( .A(n6535), .ZN(n5822) );
  INV_X1 U2668 ( .A(D_DATA_INBUS[12]), .ZN(n5821) );
  INV_X1 U2669 ( .A(n6524), .ZN(n5814) );
  INV_X1 U2670 ( .A(n6537), .ZN(n5812) );
  INV_X1 U2671 ( .A(D_DATA_INBUS[13]), .ZN(n5811) );
  INV_X1 U2672 ( .A(n6525), .ZN(n5803) );
  INV_X1 U2673 ( .A(n6539), .ZN(n5800) );
  INV_X1 U2674 ( .A(D_DATA_INBUS[14]), .ZN(n5799) );
  INV_X1 U2675 ( .A(n6541), .ZN(n5791) );
  INV_X1 U2676 ( .A(n6546), .ZN(n5789) );
  NAND2_X1 U2677 ( .A1(n5999), .A2(\Mpath/the_memhandle/N34 ), .ZN(n5785) );
  AND2_X1 U2678 ( .A1(n1852), .A2(n1853), .ZN(n5715) );
  AOI222_X1 U2679 ( .A1(\Mpath/the_shift/sh_rol [0]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [0]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [0]), .C2(n1703), .ZN(n1853) );
  AOI22_X1 U2680 ( .A1(\Mpath/the_shift/sh_sra [0]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [0]), .B2(\Mpath/the_shift/N118 ), .ZN(n1852)
         );
  INV_X1 U2681 ( .A(n6977), .ZN(n5714) );
  INV_X1 U2682 ( .A(n1854), .ZN(n5707) );
  OAI211_X1 U2683 ( .C1(\Mpath/the_alu/N35 ), .C2(n7315), .A(n1855), .B(n1856), 
        .ZN(n1854) );
  AOI22_X1 U2684 ( .A1(\Mpath/the_alu/diff[24] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[24] ), .B2(n7634), .ZN(n1856) );
  AOI22_X1 U2685 ( .A1(\Mpath/the_alu/N36 ), .A2(n1857), .B1(n1858), .B2(n327), 
        .ZN(n1855) );
  INV_X1 U2686 ( .A(\Mpath/the_alu/N36 ), .ZN(n327) );
  OAI22_X1 U2688 ( .A1(n1692), .A2(n1859), .B1(\Mpath/the_alu/N35 ), .B2(n1841), .ZN(n1857) );
  INV_X1 U2689 ( .A(\Mpath/the_alu/N35 ), .ZN(n1859) );
  AND2_X1 U2690 ( .A1(n1860), .A2(n1861), .ZN(n5706) );
  AOI222_X1 U2691 ( .A1(\Mpath/the_shift/sh_rol [24]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [24]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [24]), .C2(n1703), .ZN(n1861) );
  AOI22_X1 U2692 ( .A1(\Mpath/the_shift/sh_sra [24]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [24]), .B2(\Mpath/the_shift/N118 ), .ZN(n1860)
         );
  INV_X1 U2693 ( .A(n1862), .ZN(n5699) );
  OAI211_X1 U2694 ( .C1(\Mpath/the_alu/N33 ), .C2(n1695), .A(n1863), .B(n1864), 
        .ZN(n1862) );
  AOI22_X1 U2695 ( .A1(\Mpath/the_alu/diff[25] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[25] ), .B2(n7634), .ZN(n1864) );
  AOI22_X1 U2696 ( .A1(\Mpath/the_alu/N34 ), .A2(n1865), .B1(n1866), .B2(n229), 
        .ZN(n1863) );
  INV_X1 U2697 ( .A(\Mpath/the_alu/N34 ), .ZN(n229) );
  OAI22_X1 U2699 ( .A1(n7187), .A2(n1867), .B1(\Mpath/the_alu/N33 ), .B2(n1841), .ZN(n1865) );
  INV_X1 U2700 ( .A(\Mpath/the_alu/N33 ), .ZN(n1867) );
  AND2_X1 U2701 ( .A1(n1868), .A2(n1869), .ZN(n5698) );
  AOI222_X1 U2702 ( .A1(\Mpath/the_shift/sh_rol [25]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [25]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [25]), .C2(n1703), .ZN(n1869) );
  AOI22_X1 U2703 ( .A1(\Mpath/the_shift/sh_sra [25]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [25]), .B2(\Mpath/the_shift/N118 ), .ZN(n1868)
         );
  INV_X1 U2704 ( .A(n1870), .ZN(n5691) );
  OAI211_X1 U2705 ( .C1(\Mpath/the_alu/N31 ), .C2(n7315), .A(n1871), .B(n1872), 
        .ZN(n1870) );
  AOI22_X1 U2706 ( .A1(\Mpath/the_alu/diff[26] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[26] ), .B2(n7634), .ZN(n1872) );
  AOI22_X1 U2707 ( .A1(\Mpath/the_alu/N32 ), .A2(n1873), .B1(n1874), .B2(n221), 
        .ZN(n1871) );
  INV_X1 U2708 ( .A(\Mpath/the_alu/N32 ), .ZN(n221) );
  OAI22_X1 U2710 ( .A1(n7187), .A2(n1875), .B1(\Mpath/the_alu/N31 ), .B2(n1841), .ZN(n1873) );
  INV_X1 U2711 ( .A(\Mpath/the_alu/N31 ), .ZN(n1875) );
  AND2_X1 U2712 ( .A1(n1876), .A2(n1877), .ZN(n5690) );
  AOI222_X1 U2713 ( .A1(\Mpath/the_shift/sh_rol [26]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [26]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [26]), .C2(n1703), .ZN(n1877) );
  AOI22_X1 U2714 ( .A1(\Mpath/the_shift/sh_sra [26]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [26]), .B2(\Mpath/the_shift/N118 ), .ZN(n1876)
         );
  INV_X1 U2715 ( .A(n1878), .ZN(n5683) );
  OAI211_X1 U2716 ( .C1(\Mpath/the_alu/N29 ), .C2(n7315), .A(n1879), .B(n1880), 
        .ZN(n1878) );
  AOI22_X1 U2717 ( .A1(\Mpath/the_alu/diff[27] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[27] ), .B2(n7634), .ZN(n1880) );
  AOI22_X1 U2718 ( .A1(\Mpath/the_alu/N30 ), .A2(n1881), .B1(n1882), .B2(n1883), .ZN(n1879) );
  INV_X1 U2719 ( .A(\Mpath/the_alu/N30 ), .ZN(n1883) );
  OAI22_X1 U2721 ( .A1(n1692), .A2(n1884), .B1(\Mpath/the_alu/N29 ), .B2(n1841), .ZN(n1881) );
  INV_X1 U2722 ( .A(\Mpath/the_alu/N29 ), .ZN(n1884) );
  AND2_X1 U2723 ( .A1(n1885), .A2(n1886), .ZN(n5682) );
  AOI222_X1 U2724 ( .A1(\Mpath/the_shift/sh_rol [27]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [27]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [27]), .C2(n1703), .ZN(n1886) );
  AOI22_X1 U2725 ( .A1(\Mpath/the_shift/sh_sra [27]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [27]), .B2(\Mpath/the_shift/N118 ), .ZN(n1885)
         );
  INV_X1 U2726 ( .A(n1887), .ZN(n5675) );
  OAI211_X1 U2727 ( .C1(\Mpath/the_alu/N27 ), .C2(n7315), .A(n1888), .B(n1889), 
        .ZN(n1887) );
  AOI22_X1 U2728 ( .A1(\Mpath/the_alu/diff[28] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[28] ), .B2(n7634), .ZN(n1889) );
  AOI22_X1 U2729 ( .A1(\Mpath/the_alu/N28 ), .A2(n1890), .B1(n1891), .B2(n1892), .ZN(n1888) );
  INV_X1 U2730 ( .A(\Mpath/the_alu/N28 ), .ZN(n1892) );
  OAI22_X1 U2732 ( .A1(n1692), .A2(n1893), .B1(\Mpath/the_alu/N27 ), .B2(n1841), .ZN(n1890) );
  INV_X1 U2733 ( .A(\Mpath/the_alu/N27 ), .ZN(n1893) );
  AND2_X1 U2734 ( .A1(n1894), .A2(n1895), .ZN(n5674) );
  AOI222_X1 U2735 ( .A1(\Mpath/the_shift/sh_rol [28]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [28]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [28]), .C2(n1703), .ZN(n1895) );
  AOI22_X1 U2736 ( .A1(\Mpath/the_shift/sh_sra [28]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [28]), .B2(\Mpath/the_shift/N118 ), .ZN(n1894)
         );
  INV_X1 U2737 ( .A(n1896), .ZN(n5667) );
  OAI211_X1 U2738 ( .C1(\Mpath/the_alu/N25 ), .C2(n7315), .A(n1897), .B(n1898), 
        .ZN(n1896) );
  AOI22_X1 U2739 ( .A1(\Mpath/the_alu/diff[29] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[29] ), .B2(n7634), .ZN(n1898) );
  AOI22_X1 U2740 ( .A1(\Mpath/the_alu/N26 ), .A2(n1899), .B1(n1900), .B2(n1901), .ZN(n1897) );
  INV_X1 U2741 ( .A(\Mpath/the_alu/N26 ), .ZN(n1901) );
  OAI22_X1 U2743 ( .A1(n1692), .A2(n1902), .B1(\Mpath/the_alu/N25 ), .B2(n1841), .ZN(n1899) );
  INV_X1 U2744 ( .A(\Mpath/the_alu/N25 ), .ZN(n1902) );
  AND2_X1 U2745 ( .A1(n1903), .A2(n1904), .ZN(n5666) );
  AOI222_X1 U2746 ( .A1(\Mpath/the_shift/sh_rol [29]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [29]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [29]), .C2(n1703), .ZN(n1904) );
  AOI22_X1 U2747 ( .A1(\Mpath/the_shift/sh_sra [29]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [29]), .B2(\Mpath/the_shift/N118 ), .ZN(n1903)
         );
  OAI211_X1 U2749 ( .C1(\Mpath/the_alu/N23 ), .C2(n1695), .A(n1906), .B(n1907), 
        .ZN(n1905) );
  AOI22_X1 U2751 ( .A1(\Mpath/the_alu/N24 ), .A2(n1908), .B1(n1909), .B2(n1910), .ZN(n1906) );
  INV_X1 U2752 ( .A(\Mpath/the_alu/N24 ), .ZN(n1910) );
  OAI22_X1 U2754 ( .A1(n1692), .A2(n1911), .B1(\Mpath/the_alu/N23 ), .B2(n1841), .ZN(n1908) );
  INV_X1 U2755 ( .A(\Mpath/the_alu/N23 ), .ZN(n1911) );
  AND2_X1 U2756 ( .A1(n1912), .A2(n1913), .ZN(n5656) );
  AOI222_X1 U2757 ( .A1(\Mpath/the_shift/sh_rol [30]), .A2(n1701), .B1(
        \Mpath/the_shift/sh_ror [30]), .B2(n6553), .C1(
        \Mpath/the_shift/sh_sll [30]), .C2(n1703), .ZN(n1913) );
  INV_X1 U2760 ( .A(\Mpath/the_shift/N111 ), .ZN(n1914) );
  INV_X1 U2762 ( .A(n6503), .ZN(n1915) );
  AOI22_X1 U2763 ( .A1(\Mpath/the_shift/sh_sra [30]), .A2(n1704), .B1(
        \Mpath/the_shift/sh_srl [30]), .B2(\Mpath/the_shift/N118 ), .ZN(n1912)
         );
  INV_X1 U2765 ( .A(\Mpath/the_shift/N115 ), .ZN(n1916) );
  INV_X1 U2766 ( .A(n181), .ZN(n5619) );
  NAND4_X1 U2767 ( .A1(n1917), .A2(n1918), .A3(n1919), .A4(n1920), .ZN(n181)
         );
  NOR4_X1 U2768 ( .A1(n1921), .A2(n1922), .A3(n1923), .A4(n1924), .ZN(n1920)
         );
  NAND3_X1 U2769 ( .A1(n6031), .A2(n6027), .A3(n6036), .ZN(n1924) );
  OAI211_X1 U2770 ( .C1(n5779), .C2(n1336), .A(n6016), .B(n6023), .ZN(n1923)
         );
  OAI222_X1 U2771 ( .A1(n5777), .A2(n1308), .B1(n7025), .B2(n1164), .C1(n5778), 
        .C2(n1192), .ZN(n1922) );
  OAI221_X1 U2772 ( .B1(n7492), .B2(n1364), .C1(n5772), .C2(n1220), .A(n1925), 
        .ZN(n1921) );
  AOI22_X1 U2773 ( .A1(\regfile/reg_out[2][0] ), .A2(n1926), .B1(
        \regfile/reg_out[3][0] ), .B2(n1927), .ZN(n1925) );
  AOI211_X1 U2774 ( .C1(\regfile/reg_out[30][0] ), .C2(n1928), .A(n1929), .B(
        n1930), .ZN(n1919) );
  OAI22_X1 U2775 ( .A1(n7026), .A2(n1250), .B1(n5760), .B2(n1122), .ZN(n1930)
         );
  OAI222_X1 U2778 ( .A1(n5755), .A2(n1136), .B1(n6906), .B2(n1280), .C1(n5759), 
        .C2(n1266), .ZN(n1929) );
  AOI221_X1 U2782 ( .B1(\regfile/reg_out[1][0] ), .B2(n1931), .C1(
        \regfile/reg_out[12][0] ), .C2(n1932), .A(n1933), .ZN(n1918) );
  OAI22_X1 U2783 ( .A1(n1934), .A2(n1206), .B1(n7017), .B2(n1322), .ZN(n1933)
         );
  AOI222_X1 U2785 ( .A1(\regfile/reg_out[16][0] ), .A2(n1936), .B1(
        \regfile/reg_out[9][0] ), .B2(n1937), .C1(\regfile/reg_out[17][0] ), 
        .C2(n1938), .ZN(n1917) );
  INV_X1 U2786 ( .A(n141), .ZN(n5616) );
  NAND4_X1 U2787 ( .A1(n1939), .A2(n1940), .A3(n1941), .A4(n1942), .ZN(n141)
         );
  NOR4_X1 U2788 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(n1942)
         );
  NAND3_X1 U2789 ( .A1(n6008), .A2(n6007), .A3(n6009), .ZN(n1946) );
  OAI211_X1 U2790 ( .C1(n5779), .C2(n682), .A(n6005), .B(n6006), .ZN(n1945) );
  OAI222_X1 U2791 ( .A1(n5777), .A2(n686), .B1(n7025), .B2(n685), .C1(n5778), 
        .C2(n681), .ZN(n1944) );
  OAI221_X1 U2792 ( .B1(n7491), .B2(n699), .C1(n5772), .C2(n698), .A(n1947), 
        .ZN(n1943) );
  AOI22_X1 U2793 ( .A1(\regfile/reg_out[2][10] ), .A2(n1926), .B1(
        \regfile/reg_out[3][10] ), .B2(n1927), .ZN(n1947) );
  AOI211_X1 U2794 ( .C1(\regfile/reg_out[30][10] ), .C2(n1928), .A(n1948), .B(
        n1949), .ZN(n1941) );
  OAI22_X1 U2795 ( .A1(n7026), .A2(n696), .B1(n5760), .B2(n692), .ZN(n1949) );
  OAI222_X1 U2798 ( .A1(n5755), .A2(n690), .B1(n6906), .B2(n691), .C1(n5759), 
        .C2(n693), .ZN(n1948) );
  AOI221_X1 U2802 ( .B1(\regfile/reg_out[1][10] ), .B2(n1931), .C1(
        \regfile/reg_out[12][10] ), .C2(n1932), .A(n1950), .ZN(n1940) );
  OAI22_X1 U2803 ( .A1(n1934), .A2(n700), .B1(n7017), .B2(n684), .ZN(n1950) );
  AOI222_X1 U2805 ( .A1(\regfile/reg_out[16][10] ), .A2(n1936), .B1(
        \regfile/reg_out[9][10] ), .B2(n1937), .C1(\regfile/reg_out[17][10] ), 
        .C2(n1938), .ZN(n1939) );
  INV_X1 U2806 ( .A(n137), .ZN(n5613) );
  NAND4_X1 U2807 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(n1954), .ZN(n137)
         );
  NOR4_X1 U2808 ( .A1(n1955), .A2(n1956), .A3(n1957), .A4(n1958), .ZN(n1954)
         );
  NAND3_X1 U2809 ( .A1(n5997), .A2(n5996), .A3(n5998), .ZN(n1958) );
  OAI211_X1 U2810 ( .C1(n5779), .C2(n720), .A(n5994), .B(n5995), .ZN(n1957) );
  OAI222_X1 U2811 ( .A1(n5777), .A2(n724), .B1(n7025), .B2(n723), .C1(n5778), 
        .C2(n719), .ZN(n1956) );
  OAI221_X1 U2812 ( .B1(n7492), .B2(n737), .C1(n5772), .C2(n736), .A(n1959), 
        .ZN(n1955) );
  AOI22_X1 U2813 ( .A1(\regfile/reg_out[2][11] ), .A2(n1926), .B1(
        \regfile/reg_out[3][11] ), .B2(n1927), .ZN(n1959) );
  AOI211_X1 U2814 ( .C1(\regfile/reg_out[30][11] ), .C2(n6892), .A(n1960), .B(
        n1961), .ZN(n1953) );
  OAI22_X1 U2815 ( .A1(n7026), .A2(n734), .B1(n5760), .B2(n730), .ZN(n1961) );
  OAI222_X1 U2818 ( .A1(n5755), .A2(n728), .B1(n6906), .B2(n729), .C1(n5759), 
        .C2(n731), .ZN(n1960) );
  AOI221_X1 U2822 ( .B1(\regfile/reg_out[1][11] ), .B2(n1931), .C1(
        \regfile/reg_out[12][11] ), .C2(n1932), .A(n1962), .ZN(n1952) );
  OAI22_X1 U2823 ( .A1(n1934), .A2(n738), .B1(n7017), .B2(n722), .ZN(n1962) );
  AOI222_X1 U2825 ( .A1(\regfile/reg_out[16][11] ), .A2(n1936), .B1(
        \regfile/reg_out[9][11] ), .B2(n1937), .C1(\regfile/reg_out[17][11] ), 
        .C2(n1938), .ZN(n1951) );
  INV_X1 U2826 ( .A(n133), .ZN(n5610) );
  NAND4_X1 U2827 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(n133)
         );
  NOR4_X1 U2828 ( .A1(n1967), .A2(n1968), .A3(n1969), .A4(n1970), .ZN(n1966)
         );
  NAND3_X1 U2829 ( .A1(n5992), .A2(n5991), .A3(n5993), .ZN(n1970) );
  OAI211_X1 U2830 ( .C1(n5779), .C2(n758), .A(n5989), .B(n5990), .ZN(n1969) );
  OAI222_X1 U2831 ( .A1(n5777), .A2(n762), .B1(n7025), .B2(n761), .C1(n5778), 
        .C2(n757), .ZN(n1968) );
  OAI221_X1 U2832 ( .B1(n7493), .B2(n775), .C1(n5772), .C2(n774), .A(n1971), 
        .ZN(n1967) );
  AOI22_X1 U2833 ( .A1(\regfile/reg_out[2][12] ), .A2(n1926), .B1(
        \regfile/reg_out[3][12] ), .B2(n1927), .ZN(n1971) );
  AOI211_X1 U2834 ( .C1(\regfile/reg_out[30][12] ), .C2(n1928), .A(n1972), .B(
        n1973), .ZN(n1965) );
  OAI22_X1 U2835 ( .A1(n7026), .A2(n772), .B1(n5760), .B2(n768), .ZN(n1973) );
  OAI222_X1 U2838 ( .A1(n5755), .A2(n766), .B1(n6906), .B2(n767), .C1(n5759), 
        .C2(n769), .ZN(n1972) );
  AOI221_X1 U2842 ( .B1(\regfile/reg_out[1][12] ), .B2(n1931), .C1(
        \regfile/reg_out[12][12] ), .C2(n1932), .A(n1974), .ZN(n1964) );
  OAI22_X1 U2843 ( .A1(n1934), .A2(n776), .B1(n7017), .B2(n760), .ZN(n1974) );
  AOI222_X1 U2845 ( .A1(\regfile/reg_out[16][12] ), .A2(n1936), .B1(
        \regfile/reg_out[9][12] ), .B2(n1937), .C1(\regfile/reg_out[17][12] ), 
        .C2(n1938), .ZN(n1963) );
  INV_X1 U2846 ( .A(n129), .ZN(n5607) );
  NAND4_X1 U2847 ( .A1(n1975), .A2(n1976), .A3(n1977), .A4(n1978), .ZN(n129)
         );
  NOR4_X1 U2848 ( .A1(n1979), .A2(n1980), .A3(n1981), .A4(n1982), .ZN(n1978)
         );
  NAND3_X1 U2849 ( .A1(n5987), .A2(n5986), .A3(n5988), .ZN(n1982) );
  OAI211_X1 U2850 ( .C1(n5779), .C2(n796), .A(n5984), .B(n5985), .ZN(n1981) );
  OAI222_X1 U2851 ( .A1(n5777), .A2(n800), .B1(n7025), .B2(n799), .C1(n5778), 
        .C2(n795), .ZN(n1980) );
  OAI221_X1 U2852 ( .B1(n7491), .B2(n813), .C1(n5772), .C2(n812), .A(n1983), 
        .ZN(n1979) );
  AOI22_X1 U2853 ( .A1(\regfile/reg_out[2][13] ), .A2(n1926), .B1(
        \regfile/reg_out[3][13] ), .B2(n1927), .ZN(n1983) );
  AOI211_X1 U2854 ( .C1(\regfile/reg_out[30][13] ), .C2(n6892), .A(n1984), .B(
        n1985), .ZN(n1977) );
  OAI22_X1 U2855 ( .A1(n7026), .A2(n810), .B1(n5760), .B2(n806), .ZN(n1985) );
  OAI222_X1 U2858 ( .A1(n5755), .A2(n804), .B1(n6906), .B2(n805), .C1(n5759), 
        .C2(n807), .ZN(n1984) );
  AOI221_X1 U2862 ( .B1(\regfile/reg_out[1][13] ), .B2(n1931), .C1(
        \regfile/reg_out[12][13] ), .C2(n1932), .A(n1986), .ZN(n1976) );
  OAI22_X1 U2863 ( .A1(n1934), .A2(n814), .B1(n7017), .B2(n798), .ZN(n1986) );
  AOI222_X1 U2865 ( .A1(\regfile/reg_out[16][13] ), .A2(n1936), .B1(
        \regfile/reg_out[9][13] ), .B2(n1937), .C1(\regfile/reg_out[17][13] ), 
        .C2(n1938), .ZN(n1975) );
  INV_X1 U2866 ( .A(n125), .ZN(n5604) );
  NAND4_X1 U2867 ( .A1(n1987), .A2(n1988), .A3(n1989), .A4(n1990), .ZN(n125)
         );
  NOR4_X1 U2868 ( .A1(n1991), .A2(n1992), .A3(n1993), .A4(n1994), .ZN(n1990)
         );
  NAND3_X1 U2869 ( .A1(n5982), .A2(n5981), .A3(n5983), .ZN(n1994) );
  OAI211_X1 U2870 ( .C1(n5779), .C2(n1335), .A(n5979), .B(n5980), .ZN(n1993)
         );
  OAI222_X1 U2871 ( .A1(n5777), .A2(n1307), .B1(n7025), .B2(n1163), .C1(n5778), 
        .C2(n1191), .ZN(n1992) );
  OAI221_X1 U2872 ( .B1(n7493), .B2(n1363), .C1(n5772), .C2(n1219), .A(n1995), 
        .ZN(n1991) );
  AOI22_X1 U2873 ( .A1(\regfile/reg_out[2][14] ), .A2(n1926), .B1(
        \regfile/reg_out[3][14] ), .B2(n1927), .ZN(n1995) );
  AOI211_X1 U2874 ( .C1(\regfile/reg_out[30][14] ), .C2(n6892), .A(n1996), .B(
        n1997), .ZN(n1989) );
  OAI22_X1 U2875 ( .A1(n7026), .A2(n1249), .B1(n5760), .B2(n1121), .ZN(n1997)
         );
  OAI222_X1 U2878 ( .A1(n5755), .A2(n1135), .B1(n6906), .B2(n1279), .C1(n5759), 
        .C2(n1265), .ZN(n1996) );
  AOI221_X1 U2882 ( .B1(\regfile/reg_out[1][14] ), .B2(n1931), .C1(
        \regfile/reg_out[12][14] ), .C2(n1932), .A(n1998), .ZN(n1988) );
  OAI22_X1 U2883 ( .A1(n1934), .A2(n1205), .B1(n7017), .B2(n1321), .ZN(n1998)
         );
  AOI222_X1 U2885 ( .A1(\regfile/reg_out[16][14] ), .A2(n1936), .B1(
        \regfile/reg_out[9][14] ), .B2(n1937), .C1(\regfile/reg_out[17][14] ), 
        .C2(n1938), .ZN(n1987) );
  INV_X1 U2886 ( .A(n121), .ZN(n5601) );
  NAND4_X1 U2887 ( .A1(n1999), .A2(n2000), .A3(n2001), .A4(n2002), .ZN(n121)
         );
  NOR4_X1 U2888 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .ZN(n2002)
         );
  NAND3_X1 U2889 ( .A1(n5977), .A2(n5976), .A3(n5978), .ZN(n2006) );
  OAI211_X1 U2890 ( .C1(n5779), .C2(n633), .A(n5974), .B(n5975), .ZN(n2005) );
  OAI222_X1 U2891 ( .A1(n5777), .A2(n637), .B1(n7025), .B2(n636), .C1(n5778), 
        .C2(n632), .ZN(n2004) );
  OAI221_X1 U2892 ( .B1(n7492), .B2(n650), .C1(n5772), .C2(n649), .A(n2007), 
        .ZN(n2003) );
  AOI22_X1 U2893 ( .A1(\regfile/reg_out[2][15] ), .A2(n1926), .B1(
        \regfile/reg_out[3][15] ), .B2(n1927), .ZN(n2007) );
  AOI211_X1 U2894 ( .C1(\regfile/reg_out[30][15] ), .C2(n1928), .A(n2008), .B(
        n2009), .ZN(n2001) );
  OAI22_X1 U2895 ( .A1(n7026), .A2(n647), .B1(n5760), .B2(n643), .ZN(n2009) );
  OAI222_X1 U2898 ( .A1(n5755), .A2(n641), .B1(n6906), .B2(n642), .C1(n5759), 
        .C2(n644), .ZN(n2008) );
  AOI221_X1 U2902 ( .B1(\regfile/reg_out[1][15] ), .B2(n1931), .C1(
        \regfile/reg_out[12][15] ), .C2(n1932), .A(n2010), .ZN(n2000) );
  OAI22_X1 U2903 ( .A1(n1934), .A2(n651), .B1(n7017), .B2(n635), .ZN(n2010) );
  AOI222_X1 U2905 ( .A1(\regfile/reg_out[16][15] ), .A2(n1936), .B1(
        \regfile/reg_out[9][15] ), .B2(n1937), .C1(\regfile/reg_out[17][15] ), 
        .C2(n1938), .ZN(n1999) );
  INV_X1 U2906 ( .A(n117), .ZN(n5598) );
  NAND4_X1 U2907 ( .A1(n2011), .A2(n2012), .A3(n2013), .A4(n2014), .ZN(n117)
         );
  NOR4_X1 U2908 ( .A1(n2015), .A2(n2016), .A3(n2017), .A4(n2018), .ZN(n2014)
         );
  NAND3_X1 U2909 ( .A1(n5972), .A2(n5971), .A3(n5973), .ZN(n2018) );
  OAI211_X1 U2910 ( .C1(n5779), .C2(n592), .A(n5969), .B(n5970), .ZN(n2017) );
  OAI222_X1 U2911 ( .A1(n5777), .A2(n596), .B1(n7025), .B2(n595), .C1(n5778), 
        .C2(n591), .ZN(n2016) );
  OAI221_X1 U2912 ( .B1(n7491), .B2(n609), .C1(n5772), .C2(n608), .A(n2019), 
        .ZN(n2015) );
  AOI22_X1 U2913 ( .A1(\regfile/reg_out[2][16] ), .A2(n1926), .B1(
        \regfile/reg_out[3][16] ), .B2(n1927), .ZN(n2019) );
  AOI211_X1 U2914 ( .C1(\regfile/reg_out[30][16] ), .C2(n6892), .A(n2020), .B(
        n2021), .ZN(n2013) );
  OAI22_X1 U2915 ( .A1(n7026), .A2(n606), .B1(n5760), .B2(n602), .ZN(n2021) );
  OAI222_X1 U2918 ( .A1(n5755), .A2(n600), .B1(n6906), .B2(n601), .C1(n5759), 
        .C2(n603), .ZN(n2020) );
  AOI221_X1 U2922 ( .B1(\regfile/reg_out[1][16] ), .B2(n1931), .C1(
        \regfile/reg_out[12][16] ), .C2(n1932), .A(n2022), .ZN(n2012) );
  OAI22_X1 U2923 ( .A1(n1934), .A2(n610), .B1(n7017), .B2(n594), .ZN(n2022) );
  AOI222_X1 U2925 ( .A1(\regfile/reg_out[16][16] ), .A2(n1936), .B1(
        \regfile/reg_out[9][16] ), .B2(n1937), .C1(\regfile/reg_out[17][16] ), 
        .C2(n1938), .ZN(n2011) );
  INV_X1 U2926 ( .A(n113), .ZN(n5595) );
  NAND4_X1 U2927 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .ZN(n113)
         );
  NOR4_X1 U2928 ( .A1(n2027), .A2(n2028), .A3(n2029), .A4(n2030), .ZN(n2026)
         );
  NAND3_X1 U2929 ( .A1(n5959), .A2(n5958), .A3(n5960), .ZN(n2030) );
  OAI211_X1 U2930 ( .C1(n5779), .C2(n557), .A(n5956), .B(n5957), .ZN(n2029) );
  OAI222_X1 U2931 ( .A1(n5777), .A2(n561), .B1(n7025), .B2(n560), .C1(n5778), 
        .C2(n556), .ZN(n2028) );
  OAI221_X1 U2932 ( .B1(n7492), .B2(n574), .C1(n5772), .C2(n573), .A(n2031), 
        .ZN(n2027) );
  AOI22_X1 U2933 ( .A1(\regfile/reg_out[2][17] ), .A2(n1926), .B1(
        \regfile/reg_out[3][17] ), .B2(n1927), .ZN(n2031) );
  AOI211_X1 U2934 ( .C1(\regfile/reg_out[30][17] ), .C2(n6892), .A(n2032), .B(
        n2033), .ZN(n2025) );
  OAI22_X1 U2935 ( .A1(n7026), .A2(n571), .B1(n5760), .B2(n567), .ZN(n2033) );
  OAI222_X1 U2938 ( .A1(n5755), .A2(n565), .B1(n6906), .B2(n566), .C1(n5759), 
        .C2(n568), .ZN(n2032) );
  AOI221_X1 U2942 ( .B1(\regfile/reg_out[1][17] ), .B2(n1931), .C1(
        \regfile/reg_out[12][17] ), .C2(n1932), .A(n2034), .ZN(n2024) );
  OAI22_X1 U2943 ( .A1(n1934), .A2(n575), .B1(n7017), .B2(n559), .ZN(n2034) );
  AOI222_X1 U2945 ( .A1(\regfile/reg_out[16][17] ), .A2(n1936), .B1(
        \regfile/reg_out[9][17] ), .B2(n1937), .C1(\regfile/reg_out[17][17] ), 
        .C2(n1938), .ZN(n2023) );
  INV_X1 U2946 ( .A(n109), .ZN(n5592) );
  NAND4_X1 U2947 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n109)
         );
  NOR4_X1 U2948 ( .A1(n2039), .A2(n2040), .A3(n2041), .A4(n2042), .ZN(n2038)
         );
  NAND3_X1 U2949 ( .A1(n5954), .A2(n5953), .A3(n5955), .ZN(n2042) );
  OAI211_X1 U2950 ( .C1(n5779), .C2(n522), .A(n5951), .B(n5952), .ZN(n2041) );
  OAI222_X1 U2951 ( .A1(n5777), .A2(n526), .B1(n7024), .B2(n525), .C1(n5778), 
        .C2(n521), .ZN(n2040) );
  OAI221_X1 U2952 ( .B1(n7492), .B2(n539), .C1(n5772), .C2(n538), .A(n2043), 
        .ZN(n2039) );
  AOI22_X1 U2953 ( .A1(\regfile/reg_out[2][18] ), .A2(n1926), .B1(
        \regfile/reg_out[3][18] ), .B2(n1927), .ZN(n2043) );
  AOI211_X1 U2954 ( .C1(\regfile/reg_out[30][18] ), .C2(n1928), .A(n2044), .B(
        n2045), .ZN(n2037) );
  OAI22_X1 U2955 ( .A1(n7026), .A2(n536), .B1(n5760), .B2(n532), .ZN(n2045) );
  OAI222_X1 U2958 ( .A1(n5755), .A2(n530), .B1(n6906), .B2(n531), .C1(n5759), 
        .C2(n533), .ZN(n2044) );
  AOI221_X1 U2962 ( .B1(\regfile/reg_out[1][18] ), .B2(n1931), .C1(
        \regfile/reg_out[12][18] ), .C2(n1932), .A(n2046), .ZN(n2036) );
  OAI22_X1 U2963 ( .A1(n1934), .A2(n540), .B1(n7017), .B2(n524), .ZN(n2046) );
  AOI222_X1 U2965 ( .A1(\regfile/reg_out[16][18] ), .A2(n1936), .B1(
        \regfile/reg_out[9][18] ), .B2(n1937), .C1(\regfile/reg_out[17][18] ), 
        .C2(n1938), .ZN(n2035) );
  INV_X1 U2966 ( .A(n105), .ZN(n5589) );
  NAND4_X1 U2967 ( .A1(n2047), .A2(n2048), .A3(n2049), .A4(n2050), .ZN(n105)
         );
  NOR4_X1 U2968 ( .A1(n2051), .A2(n2052), .A3(n2053), .A4(n2054), .ZN(n2050)
         );
  NAND3_X1 U2969 ( .A1(n5949), .A2(n5948), .A3(n5950), .ZN(n2054) );
  OAI211_X1 U2970 ( .C1(n5779), .C2(n487), .A(n5946), .B(n5947), .ZN(n2053) );
  OAI222_X1 U2971 ( .A1(n5777), .A2(n491), .B1(n7024), .B2(n490), .C1(n5778), 
        .C2(n486), .ZN(n2052) );
  OAI221_X1 U2972 ( .B1(n7491), .B2(n504), .C1(n5772), .C2(n503), .A(n2055), 
        .ZN(n2051) );
  AOI22_X1 U2973 ( .A1(\regfile/reg_out[2][19] ), .A2(n1926), .B1(
        \regfile/reg_out[3][19] ), .B2(n1927), .ZN(n2055) );
  AOI211_X1 U2974 ( .C1(\regfile/reg_out[30][19] ), .C2(n1928), .A(n2056), .B(
        n2057), .ZN(n2049) );
  OAI22_X1 U2975 ( .A1(n7026), .A2(n501), .B1(n5760), .B2(n497), .ZN(n2057) );
  OAI222_X1 U2978 ( .A1(n5755), .A2(n495), .B1(n6906), .B2(n496), .C1(n5759), 
        .C2(n498), .ZN(n2056) );
  AOI221_X1 U2982 ( .B1(\regfile/reg_out[1][19] ), .B2(n1931), .C1(
        \regfile/reg_out[12][19] ), .C2(n1932), .A(n2058), .ZN(n2048) );
  OAI22_X1 U2983 ( .A1(n1934), .A2(n505), .B1(n7017), .B2(n489), .ZN(n2058) );
  AOI222_X1 U2985 ( .A1(\regfile/reg_out[16][19] ), .A2(n1936), .B1(
        \regfile/reg_out[9][19] ), .B2(n1937), .C1(\regfile/reg_out[17][19] ), 
        .C2(n1938), .ZN(n2047) );
  INV_X1 U2986 ( .A(n177), .ZN(n5586) );
  NAND4_X1 U2987 ( .A1(n2059), .A2(n2060), .A3(n2061), .A4(n2062), .ZN(n177)
         );
  NOR4_X1 U2988 ( .A1(n2063), .A2(n2064), .A3(n2065), .A4(n2066), .ZN(n2062)
         );
  NAND3_X1 U2989 ( .A1(n5944), .A2(n5943), .A3(n5945), .ZN(n2066) );
  OAI211_X1 U2990 ( .C1(n5779), .C2(n1334), .A(n5941), .B(n5942), .ZN(n2065)
         );
  OAI222_X1 U2991 ( .A1(n5777), .A2(n1306), .B1(n7025), .B2(n1162), .C1(n5778), 
        .C2(n1190), .ZN(n2064) );
  OAI221_X1 U2992 ( .B1(n7492), .B2(n1362), .C1(n5772), .C2(n1218), .A(n2067), 
        .ZN(n2063) );
  AOI22_X1 U2993 ( .A1(\regfile/reg_out[2][1] ), .A2(n1926), .B1(
        \regfile/reg_out[3][1] ), .B2(n1927), .ZN(n2067) );
  AOI211_X1 U2994 ( .C1(\regfile/reg_out[30][1] ), .C2(n6892), .A(n2068), .B(
        n2069), .ZN(n2061) );
  OAI22_X1 U2995 ( .A1(n7026), .A2(n1248), .B1(n5760), .B2(n1120), .ZN(n2069)
         );
  OAI222_X1 U2998 ( .A1(n5755), .A2(n1134), .B1(n6906), .B2(n1278), .C1(n5759), 
        .C2(n1264), .ZN(n2068) );
  AOI221_X1 U3002 ( .B1(\regfile/reg_out[1][1] ), .B2(n1931), .C1(
        \regfile/reg_out[12][1] ), .C2(n1932), .A(n2070), .ZN(n2060) );
  OAI22_X1 U3003 ( .A1(n1934), .A2(n1204), .B1(n7017), .B2(n1320), .ZN(n2070)
         );
  AOI222_X1 U3005 ( .A1(\regfile/reg_out[16][1] ), .A2(n1936), .B1(
        \regfile/reg_out[9][1] ), .B2(n1937), .C1(\regfile/reg_out[17][1] ), 
        .C2(n1938), .ZN(n2059) );
  INV_X1 U3006 ( .A(n101), .ZN(n5583) );
  NAND4_X1 U3007 ( .A1(n2071), .A2(n2072), .A3(n2073), .A4(n2074), .ZN(n101)
         );
  NOR4_X1 U3008 ( .A1(n2075), .A2(n2076), .A3(n2077), .A4(n2078), .ZN(n2074)
         );
  NAND3_X1 U3009 ( .A1(n5933), .A2(n5932), .A3(n5934), .ZN(n2078) );
  OAI211_X1 U3010 ( .C1(n5779), .C2(n452), .A(n5930), .B(n5931), .ZN(n2077) );
  OAI222_X1 U3011 ( .A1(n5777), .A2(n456), .B1(n7025), .B2(n455), .C1(n5778), 
        .C2(n451), .ZN(n2076) );
  OAI221_X1 U3012 ( .B1(n7492), .B2(n469), .C1(n5772), .C2(n468), .A(n2079), 
        .ZN(n2075) );
  AOI22_X1 U3013 ( .A1(\regfile/reg_out[2][20] ), .A2(n1926), .B1(
        \regfile/reg_out[3][20] ), .B2(n1927), .ZN(n2079) );
  AOI211_X1 U3014 ( .C1(\regfile/reg_out[30][20] ), .C2(n1928), .A(n2080), .B(
        n2081), .ZN(n2073) );
  OAI22_X1 U3015 ( .A1(n7026), .A2(n466), .B1(n5760), .B2(n462), .ZN(n2081) );
  OAI222_X1 U3018 ( .A1(n5755), .A2(n460), .B1(n6906), .B2(n461), .C1(n5759), 
        .C2(n463), .ZN(n2080) );
  AOI221_X1 U3022 ( .B1(\regfile/reg_out[1][20] ), .B2(n1931), .C1(
        \regfile/reg_out[12][20] ), .C2(n1932), .A(n2082), .ZN(n2072) );
  OAI22_X1 U3023 ( .A1(n1934), .A2(n470), .B1(n7017), .B2(n454), .ZN(n2082) );
  AOI222_X1 U3025 ( .A1(\regfile/reg_out[16][20] ), .A2(n1936), .B1(
        \regfile/reg_out[9][20] ), .B2(n1937), .C1(\regfile/reg_out[17][20] ), 
        .C2(n1938), .ZN(n2071) );
  INV_X1 U3026 ( .A(n97), .ZN(n5580) );
  NAND4_X1 U3027 ( .A1(n2083), .A2(n2084), .A3(n2085), .A4(n2086), .ZN(n97) );
  NOR4_X1 U3028 ( .A1(n2087), .A2(n2088), .A3(n2089), .A4(n2090), .ZN(n2086)
         );
  NAND3_X1 U3029 ( .A1(n5928), .A2(n5927), .A3(n5929), .ZN(n2090) );
  OAI211_X1 U3030 ( .C1(n5779), .C2(n417), .A(n5925), .B(n5926), .ZN(n2089) );
  OAI222_X1 U3031 ( .A1(n5777), .A2(n421), .B1(n7024), .B2(n420), .C1(n5778), 
        .C2(n416), .ZN(n2088) );
  OAI221_X1 U3032 ( .B1(n7491), .B2(n434), .C1(n5772), .C2(n433), .A(n2091), 
        .ZN(n2087) );
  AOI22_X1 U3033 ( .A1(\regfile/reg_out[2][21] ), .A2(n1926), .B1(
        \regfile/reg_out[3][21] ), .B2(n1927), .ZN(n2091) );
  AOI211_X1 U3034 ( .C1(\regfile/reg_out[30][21] ), .C2(n6892), .A(n2092), .B(
        n2093), .ZN(n2085) );
  OAI22_X1 U3035 ( .A1(n7026), .A2(n431), .B1(n5760), .B2(n427), .ZN(n2093) );
  OAI222_X1 U3038 ( .A1(n5755), .A2(n425), .B1(n6906), .B2(n426), .C1(n5759), 
        .C2(n428), .ZN(n2092) );
  AOI221_X1 U3042 ( .B1(\regfile/reg_out[1][21] ), .B2(n1931), .C1(
        \regfile/reg_out[12][21] ), .C2(n1932), .A(n2094), .ZN(n2084) );
  OAI22_X1 U3043 ( .A1(n1934), .A2(n435), .B1(n7017), .B2(n419), .ZN(n2094) );
  AOI222_X1 U3045 ( .A1(\regfile/reg_out[16][21] ), .A2(n1936), .B1(
        \regfile/reg_out[9][21] ), .B2(n1937), .C1(\regfile/reg_out[17][21] ), 
        .C2(n1938), .ZN(n2083) );
  NOR4_X1 U3048 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .ZN(n2098)
         );
  NAND3_X1 U3049 ( .A1(n5923), .A2(n5922), .A3(n5924), .ZN(n2102) );
  OAI211_X1 U3050 ( .C1(n5779), .C2(n381), .A(n5920), .B(n5921), .ZN(n2101) );
  OAI222_X1 U3051 ( .A1(n5777), .A2(n385), .B1(n7024), .B2(n384), .C1(n5778), 
        .C2(n380), .ZN(n2100) );
  OAI221_X1 U3052 ( .B1(n7492), .B2(n398), .C1(n5772), .C2(n397), .A(n2103), 
        .ZN(n2099) );
  AOI22_X1 U3053 ( .A1(\regfile/reg_out[2][22] ), .A2(n1926), .B1(
        \regfile/reg_out[3][22] ), .B2(n1927), .ZN(n2103) );
  AOI211_X1 U3054 ( .C1(\regfile/reg_out[30][22] ), .C2(n6892), .A(n2104), .B(
        n2105), .ZN(n2097) );
  OAI22_X1 U3055 ( .A1(n7026), .A2(n395), .B1(n5760), .B2(n391), .ZN(n2105) );
  OAI222_X1 U3058 ( .A1(n5755), .A2(n389), .B1(n6906), .B2(n390), .C1(n5759), 
        .C2(n392), .ZN(n2104) );
  AOI221_X1 U3062 ( .B1(\regfile/reg_out[1][22] ), .B2(n1931), .C1(
        \regfile/reg_out[12][22] ), .C2(n1932), .A(n2106), .ZN(n2096) );
  OAI22_X1 U3063 ( .A1(n1934), .A2(n399), .B1(n7017), .B2(n383), .ZN(n2106) );
  AOI222_X1 U3065 ( .A1(\regfile/reg_out[16][22] ), .A2(n1936), .B1(
        \regfile/reg_out[9][22] ), .B2(n1937), .C1(\regfile/reg_out[17][22] ), 
        .C2(n1938), .ZN(n2095) );
  INV_X1 U3066 ( .A(n89), .ZN(n5574) );
  NAND4_X1 U3067 ( .A1(n2107), .A2(n2108), .A3(n2109), .A4(n2110), .ZN(n89) );
  NOR4_X1 U3068 ( .A1(n2111), .A2(n2112), .A3(n2113), .A4(n2114), .ZN(n2110)
         );
  NAND3_X1 U3069 ( .A1(n5918), .A2(n5917), .A3(n5919), .ZN(n2114) );
  OAI211_X1 U3070 ( .C1(n5779), .C2(n1333), .A(n5915), .B(n5916), .ZN(n2113)
         );
  OAI222_X1 U3071 ( .A1(n5777), .A2(n1305), .B1(n7025), .B2(n1161), .C1(n5778), 
        .C2(n1189), .ZN(n2112) );
  OAI221_X1 U3072 ( .B1(n7492), .B2(n1361), .C1(n5772), .C2(n1217), .A(n2115), 
        .ZN(n2111) );
  AOI22_X1 U3073 ( .A1(\regfile/reg_out[2][23] ), .A2(n1926), .B1(
        \regfile/reg_out[3][23] ), .B2(n1927), .ZN(n2115) );
  AOI211_X1 U3074 ( .C1(\regfile/reg_out[30][23] ), .C2(n6892), .A(n2116), .B(
        n2117), .ZN(n2109) );
  OAI22_X1 U3075 ( .A1(n7026), .A2(n1247), .B1(n5760), .B2(n1119), .ZN(n2117)
         );
  OAI222_X1 U3078 ( .A1(n5755), .A2(n1133), .B1(n6906), .B2(n1277), .C1(n5759), 
        .C2(n1263), .ZN(n2116) );
  AOI221_X1 U3082 ( .B1(\regfile/reg_out[1][23] ), .B2(n1931), .C1(
        \regfile/reg_out[12][23] ), .C2(n1932), .A(n2118), .ZN(n2108) );
  OAI22_X1 U3083 ( .A1(n1934), .A2(n1203), .B1(n7017), .B2(n1319), .ZN(n2118)
         );
  AOI222_X1 U3085 ( .A1(\regfile/reg_out[16][23] ), .A2(n1936), .B1(
        \regfile/reg_out[9][23] ), .B2(n1937), .C1(\regfile/reg_out[17][23] ), 
        .C2(n1938), .ZN(n2107) );
  INV_X1 U3086 ( .A(n85), .ZN(n5571) );
  NAND4_X1 U3087 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(n85) );
  NOR4_X1 U3088 ( .A1(n2123), .A2(n2124), .A3(n2125), .A4(n2126), .ZN(n2122)
         );
  NAND3_X1 U3089 ( .A1(n5909), .A2(n5908), .A3(n5910), .ZN(n2126) );
  OAI211_X1 U3090 ( .C1(n5779), .C2(n337), .A(n5906), .B(n5907), .ZN(n2125) );
  OAI222_X1 U3091 ( .A1(n5777), .A2(n341), .B1(n7025), .B2(n340), .C1(n5778), 
        .C2(n336), .ZN(n2124) );
  OAI221_X1 U3092 ( .B1(n7491), .B2(n354), .C1(n5772), .C2(n353), .A(n2127), 
        .ZN(n2123) );
  AOI22_X1 U3093 ( .A1(\regfile/reg_out[2][24] ), .A2(n1926), .B1(
        \regfile/reg_out[3][24] ), .B2(n1927), .ZN(n2127) );
  AOI211_X1 U3094 ( .C1(\regfile/reg_out[30][24] ), .C2(n6892), .A(n2128), .B(
        n2129), .ZN(n2121) );
  OAI22_X1 U3095 ( .A1(n7026), .A2(n351), .B1(n5760), .B2(n347), .ZN(n2129) );
  OAI222_X1 U3098 ( .A1(n5755), .A2(n345), .B1(n6906), .B2(n346), .C1(n5759), 
        .C2(n348), .ZN(n2128) );
  AOI221_X1 U3102 ( .B1(\regfile/reg_out[1][24] ), .B2(n1931), .C1(
        \regfile/reg_out[12][24] ), .C2(n1932), .A(n2130), .ZN(n2120) );
  OAI22_X1 U3103 ( .A1(n1934), .A2(n355), .B1(n7017), .B2(n339), .ZN(n2130) );
  AOI222_X1 U3105 ( .A1(\regfile/reg_out[16][24] ), .A2(n1936), .B1(
        \regfile/reg_out[9][24] ), .B2(n1937), .C1(\regfile/reg_out[17][24] ), 
        .C2(n1938), .ZN(n2119) );
  INV_X1 U3106 ( .A(n81), .ZN(n5568) );
  NAND4_X1 U3107 ( .A1(n2131), .A2(n2132), .A3(n2133), .A4(n2134), .ZN(n81) );
  NOR4_X1 U3108 ( .A1(n2135), .A2(n2136), .A3(n2137), .A4(n2138), .ZN(n2134)
         );
  NAND3_X1 U3109 ( .A1(n5899), .A2(n5898), .A3(n5900), .ZN(n2138) );
  OAI211_X1 U3110 ( .C1(n5779), .C2(n241), .A(n5896), .B(n5897), .ZN(n2137) );
  OAI222_X1 U3111 ( .A1(n5777), .A2(n253), .B1(n7025), .B2(n250), .C1(n5778), 
        .C2(n238), .ZN(n2136) );
  OAI221_X1 U3112 ( .B1(n7493), .B2(n312), .C1(n5772), .C2(n309), .A(n2139), 
        .ZN(n2135) );
  AOI22_X1 U3113 ( .A1(\regfile/reg_out[2][25] ), .A2(n1926), .B1(
        \regfile/reg_out[3][25] ), .B2(n1927), .ZN(n2139) );
  AOI211_X1 U3114 ( .C1(\regfile/reg_out[30][25] ), .C2(n1928), .A(n2140), .B(
        n2141), .ZN(n2133) );
  OAI22_X1 U3115 ( .A1(n7026), .A2(n299), .B1(n5760), .B2(n283), .ZN(n2141) );
  OAI222_X1 U3118 ( .A1(n5755), .A2(n273), .B1(n6906), .B2(n276), .C1(n5759), 
        .C2(n286), .ZN(n2140) );
  AOI221_X1 U3122 ( .B1(\regfile/reg_out[1][25] ), .B2(n1931), .C1(
        \regfile/reg_out[12][25] ), .C2(n1932), .A(n2142), .ZN(n2132) );
  OAI22_X1 U3123 ( .A1(n1934), .A2(n315), .B1(n7017), .B2(n247), .ZN(n2142) );
  AOI222_X1 U3125 ( .A1(\regfile/reg_out[16][25] ), .A2(n1936), .B1(
        \regfile/reg_out[9][25] ), .B2(n1937), .C1(\regfile/reg_out[17][25] ), 
        .C2(n1938), .ZN(n2131) );
  INV_X1 U3126 ( .A(n77), .ZN(n5565) );
  NAND4_X1 U3127 ( .A1(n2143), .A2(n2144), .A3(n2145), .A4(n2146), .ZN(n77) );
  NOR4_X1 U3128 ( .A1(n2147), .A2(n2148), .A3(n2149), .A4(n2150), .ZN(n2146)
         );
  NAND3_X1 U3129 ( .A1(n5888), .A2(n5887), .A3(n5889), .ZN(n2150) );
  OAI211_X1 U3130 ( .C1(n5779), .C2(n1332), .A(n5885), .B(n5886), .ZN(n2149)
         );
  OAI222_X1 U3131 ( .A1(n5777), .A2(n1304), .B1(n7025), .B2(n1160), .C1(n5778), 
        .C2(n1188), .ZN(n2148) );
  OAI221_X1 U3132 ( .B1(n7492), .B2(n1360), .C1(n5772), .C2(n1216), .A(n2151), 
        .ZN(n2147) );
  AOI22_X1 U3133 ( .A1(\regfile/reg_out[2][26] ), .A2(n1926), .B1(
        \regfile/reg_out[3][26] ), .B2(n1927), .ZN(n2151) );
  AOI211_X1 U3134 ( .C1(\regfile/reg_out[30][26] ), .C2(n1928), .A(n2152), .B(
        n2153), .ZN(n2145) );
  OAI22_X1 U3135 ( .A1(n7026), .A2(n1246), .B1(n5760), .B2(n1118), .ZN(n2153)
         );
  OAI222_X1 U3138 ( .A1(n5755), .A2(n1132), .B1(n6906), .B2(n1276), .C1(n5759), 
        .C2(n1262), .ZN(n2152) );
  AOI221_X1 U3142 ( .B1(\regfile/reg_out[1][26] ), .B2(n1931), .C1(
        \regfile/reg_out[12][26] ), .C2(n1932), .A(n2154), .ZN(n2144) );
  OAI22_X1 U3143 ( .A1(n1934), .A2(n1202), .B1(n7017), .B2(n1318), .ZN(n2154)
         );
  AOI222_X1 U3145 ( .A1(\regfile/reg_out[16][26] ), .A2(n1936), .B1(
        \regfile/reg_out[9][26] ), .B2(n1937), .C1(\regfile/reg_out[17][26] ), 
        .C2(n1938), .ZN(n2143) );
  INV_X1 U3146 ( .A(n73), .ZN(n5562) );
  NAND4_X1 U3147 ( .A1(n2155), .A2(n2156), .A3(n2157), .A4(n2158), .ZN(n73) );
  NOR4_X1 U3148 ( .A1(n2159), .A2(n2160), .A3(n2161), .A4(n2162), .ZN(n2158)
         );
  NAND3_X1 U3149 ( .A1(n5878), .A2(n5877), .A3(n5879), .ZN(n2162) );
  OAI211_X1 U3150 ( .C1(n5779), .C2(n1331), .A(n5875), .B(n5876), .ZN(n2161)
         );
  OAI222_X1 U3151 ( .A1(n5777), .A2(n1303), .B1(n7024), .B2(n1159), .C1(n5778), 
        .C2(n1187), .ZN(n2160) );
  OAI221_X1 U3152 ( .B1(n7492), .B2(n1359), .C1(n5772), .C2(n1215), .A(n2163), 
        .ZN(n2159) );
  AOI22_X1 U3153 ( .A1(\regfile/reg_out[2][27] ), .A2(n1926), .B1(
        \regfile/reg_out[3][27] ), .B2(n1927), .ZN(n2163) );
  AOI211_X1 U3154 ( .C1(\regfile/reg_out[30][27] ), .C2(n6892), .A(n2164), .B(
        n2165), .ZN(n2157) );
  OAI22_X1 U3155 ( .A1(n7026), .A2(n1245), .B1(n5760), .B2(n1117), .ZN(n2165)
         );
  OAI222_X1 U3158 ( .A1(n5755), .A2(n1131), .B1(n6906), .B2(n1275), .C1(n5759), 
        .C2(n1261), .ZN(n2164) );
  AOI221_X1 U3162 ( .B1(\regfile/reg_out[1][27] ), .B2(n1931), .C1(
        \regfile/reg_out[12][27] ), .C2(n1932), .A(n2166), .ZN(n2156) );
  OAI22_X1 U3163 ( .A1(n1934), .A2(n1201), .B1(n7017), .B2(n1317), .ZN(n2166)
         );
  AOI222_X1 U3165 ( .A1(\regfile/reg_out[16][27] ), .A2(n1936), .B1(
        \regfile/reg_out[9][27] ), .B2(n1937), .C1(\regfile/reg_out[17][27] ), 
        .C2(n1938), .ZN(n2155) );
  INV_X1 U3166 ( .A(n69), .ZN(n5559) );
  NAND4_X1 U3167 ( .A1(n2167), .A2(n2168), .A3(n2169), .A4(n2170), .ZN(n69) );
  NOR4_X1 U3168 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(n2170)
         );
  NAND3_X1 U3169 ( .A1(n5873), .A2(n5872), .A3(n5874), .ZN(n2174) );
  OAI211_X1 U3170 ( .C1(n5779), .C2(n1330), .A(n5870), .B(n5871), .ZN(n2173)
         );
  OAI222_X1 U3171 ( .A1(n5777), .A2(n1302), .B1(n7024), .B2(n1158), .C1(n5778), 
        .C2(n1186), .ZN(n2172) );
  OAI221_X1 U3172 ( .B1(n7493), .B2(n1358), .C1(n5772), .C2(n1214), .A(n2175), 
        .ZN(n2171) );
  AOI22_X1 U3173 ( .A1(\regfile/reg_out[2][28] ), .A2(n1926), .B1(
        \regfile/reg_out[3][28] ), .B2(n1927), .ZN(n2175) );
  AOI211_X1 U3174 ( .C1(\regfile/reg_out[30][28] ), .C2(n1928), .A(n2176), .B(
        n2177), .ZN(n2169) );
  OAI22_X1 U3175 ( .A1(n7026), .A2(n1244), .B1(n5760), .B2(n1116), .ZN(n2177)
         );
  OAI222_X1 U3178 ( .A1(n5755), .A2(n1130), .B1(n6906), .B2(n1274), .C1(n5759), 
        .C2(n1260), .ZN(n2176) );
  AOI221_X1 U3182 ( .B1(\regfile/reg_out[1][28] ), .B2(n1931), .C1(
        \regfile/reg_out[12][28] ), .C2(n1932), .A(n2178), .ZN(n2168) );
  OAI22_X1 U3183 ( .A1(n1934), .A2(n1200), .B1(n7017), .B2(n1316), .ZN(n2178)
         );
  AOI222_X1 U3185 ( .A1(\regfile/reg_out[16][28] ), .A2(n1936), .B1(
        \regfile/reg_out[9][28] ), .B2(n1937), .C1(\regfile/reg_out[17][28] ), 
        .C2(n1938), .ZN(n2167) );
  INV_X1 U3186 ( .A(n65), .ZN(n5556) );
  NAND4_X1 U3187 ( .A1(n2179), .A2(n2180), .A3(n2181), .A4(n2182), .ZN(n65) );
  NOR4_X1 U3188 ( .A1(n2183), .A2(n2184), .A3(n2185), .A4(n2186), .ZN(n2182)
         );
  NAND3_X1 U3189 ( .A1(n5868), .A2(n5867), .A3(n5869), .ZN(n2186) );
  OAI211_X1 U3190 ( .C1(n5779), .C2(n1329), .A(n5865), .B(n5866), .ZN(n2185)
         );
  OAI222_X1 U3191 ( .A1(n5777), .A2(n1301), .B1(n7025), .B2(n1157), .C1(n5778), 
        .C2(n1185), .ZN(n2184) );
  OAI221_X1 U3192 ( .B1(n7493), .B2(n1357), .C1(n5772), .C2(n1213), .A(n2187), 
        .ZN(n2183) );
  AOI22_X1 U3193 ( .A1(\regfile/reg_out[2][29] ), .A2(n1926), .B1(
        \regfile/reg_out[3][29] ), .B2(n1927), .ZN(n2187) );
  AOI211_X1 U3194 ( .C1(\regfile/reg_out[30][29] ), .C2(n1928), .A(n2188), .B(
        n2189), .ZN(n2181) );
  OAI22_X1 U3195 ( .A1(n7026), .A2(n1243), .B1(n5760), .B2(n1115), .ZN(n2189)
         );
  OAI222_X1 U3198 ( .A1(n5755), .A2(n1129), .B1(n6906), .B2(n1273), .C1(n5759), 
        .C2(n1259), .ZN(n2188) );
  AOI221_X1 U3202 ( .B1(\regfile/reg_out[1][29] ), .B2(n1931), .C1(
        \regfile/reg_out[12][29] ), .C2(n1932), .A(n2190), .ZN(n2180) );
  OAI22_X1 U3203 ( .A1(n1934), .A2(n1199), .B1(n7017), .B2(n1315), .ZN(n2190)
         );
  AOI222_X1 U3205 ( .A1(\regfile/reg_out[16][29] ), .A2(n1936), .B1(
        \regfile/reg_out[9][29] ), .B2(n1937), .C1(\regfile/reg_out[17][29] ), 
        .C2(n1938), .ZN(n2179) );
  INV_X1 U3206 ( .A(n173), .ZN(n5553) );
  NAND4_X1 U3207 ( .A1(n2191), .A2(n2192), .A3(n2193), .A4(n2194), .ZN(n173)
         );
  NOR4_X1 U3208 ( .A1(n2195), .A2(n2196), .A3(n2197), .A4(n2198), .ZN(n2194)
         );
  NAND3_X1 U3209 ( .A1(n5863), .A2(n5862), .A3(n5864), .ZN(n2198) );
  OAI211_X1 U3210 ( .C1(n5779), .C2(n1328), .A(n5860), .B(n5861), .ZN(n2197)
         );
  OAI222_X1 U3211 ( .A1(n5777), .A2(n1300), .B1(n7025), .B2(n1156), .C1(n5778), 
        .C2(n1184), .ZN(n2196) );
  OAI221_X1 U3212 ( .B1(n7493), .B2(n1356), .C1(n5772), .C2(n1212), .A(n2199), 
        .ZN(n2195) );
  AOI22_X1 U3213 ( .A1(\regfile/reg_out[2][2] ), .A2(n1926), .B1(
        \regfile/reg_out[3][2] ), .B2(n1927), .ZN(n2199) );
  AOI211_X1 U3214 ( .C1(\regfile/reg_out[30][2] ), .C2(n1928), .A(n2200), .B(
        n2201), .ZN(n2193) );
  OAI22_X1 U3215 ( .A1(n7026), .A2(n1242), .B1(n5760), .B2(n1114), .ZN(n2201)
         );
  OAI222_X1 U3218 ( .A1(n5755), .A2(n1128), .B1(n6906), .B2(n1272), .C1(n5759), 
        .C2(n1258), .ZN(n2200) );
  AOI221_X1 U3222 ( .B1(\regfile/reg_out[1][2] ), .B2(n1931), .C1(
        \regfile/reg_out[12][2] ), .C2(n1932), .A(n2202), .ZN(n2192) );
  OAI22_X1 U3223 ( .A1(n1934), .A2(n1198), .B1(n7017), .B2(n1314), .ZN(n2202)
         );
  AOI222_X1 U3225 ( .A1(\regfile/reg_out[16][2] ), .A2(n1936), .B1(
        \regfile/reg_out[9][2] ), .B2(n1937), .C1(\regfile/reg_out[17][2] ), 
        .C2(n1938), .ZN(n2191) );
  INV_X1 U3226 ( .A(n61), .ZN(n5550) );
  NAND4_X1 U3227 ( .A1(n2203), .A2(n2204), .A3(n2205), .A4(n2206), .ZN(n61) );
  NOR4_X1 U3228 ( .A1(n2207), .A2(n2208), .A3(n2209), .A4(n2210), .ZN(n2206)
         );
  NAND3_X1 U3229 ( .A1(n5852), .A2(n5851), .A3(n5853), .ZN(n2210) );
  OAI211_X1 U3230 ( .C1(n5779), .C2(n1327), .A(n5849), .B(n5850), .ZN(n2209)
         );
  OAI222_X1 U3231 ( .A1(n5777), .A2(n1299), .B1(n7024), .B2(n1155), .C1(n5778), 
        .C2(n1183), .ZN(n2208) );
  OAI221_X1 U3232 ( .B1(n7493), .B2(n1355), .C1(n5772), .C2(n1211), .A(n2211), 
        .ZN(n2207) );
  AOI22_X1 U3233 ( .A1(\regfile/reg_out[2][30] ), .A2(n1926), .B1(
        \regfile/reg_out[3][30] ), .B2(n1927), .ZN(n2211) );
  AOI211_X1 U3234 ( .C1(\regfile/reg_out[30][30] ), .C2(n6892), .A(n2212), .B(
        n2213), .ZN(n2205) );
  OAI22_X1 U3235 ( .A1(n7026), .A2(n1241), .B1(n5760), .B2(n1113), .ZN(n2213)
         );
  OAI222_X1 U3238 ( .A1(n5755), .A2(n1127), .B1(n6906), .B2(n1271), .C1(n5759), 
        .C2(n1257), .ZN(n2212) );
  AOI221_X1 U3242 ( .B1(\regfile/reg_out[1][30] ), .B2(n1931), .C1(
        \regfile/reg_out[12][30] ), .C2(n1932), .A(n2214), .ZN(n2204) );
  OAI22_X1 U3243 ( .A1(n1934), .A2(n1197), .B1(n7017), .B2(n1313), .ZN(n2214)
         );
  AOI222_X1 U3245 ( .A1(\regfile/reg_out[16][30] ), .A2(n1936), .B1(
        \regfile/reg_out[9][30] ), .B2(n1937), .C1(\regfile/reg_out[17][30] ), 
        .C2(n1938), .ZN(n2203) );
  INV_X1 U3246 ( .A(n56), .ZN(n5547) );
  NAND4_X1 U3247 ( .A1(n2215), .A2(n2216), .A3(n2217), .A4(n2218), .ZN(n56) );
  NOR4_X1 U3248 ( .A1(n2219), .A2(n2220), .A3(n2221), .A4(n2222), .ZN(n2218)
         );
  NAND3_X1 U3249 ( .A1(n5843), .A2(n5842), .A3(n5844), .ZN(n2222) );
  OAI211_X1 U3250 ( .C1(n5779), .C2(n1326), .A(n5840), .B(n5841), .ZN(n2221)
         );
  OAI222_X1 U3251 ( .A1(n5777), .A2(n1298), .B1(n7024), .B2(n1154), .C1(n5778), 
        .C2(n1182), .ZN(n2220) );
  OAI221_X1 U3252 ( .B1(n7493), .B2(n1354), .C1(n5772), .C2(n1210), .A(n2223), 
        .ZN(n2219) );
  AOI22_X1 U3253 ( .A1(\regfile/reg_out[2][31] ), .A2(n1926), .B1(
        \regfile/reg_out[3][31] ), .B2(n1927), .ZN(n2223) );
  AOI211_X1 U3254 ( .C1(\regfile/reg_out[30][31] ), .C2(n1928), .A(n2224), .B(
        n2225), .ZN(n2217) );
  OAI22_X1 U3255 ( .A1(n7026), .A2(n1240), .B1(n5760), .B2(n1112), .ZN(n2225)
         );
  OAI222_X1 U3258 ( .A1(n5755), .A2(n1126), .B1(n6906), .B2(n1270), .C1(n5759), 
        .C2(n1256), .ZN(n2224) );
  AOI221_X1 U3262 ( .B1(\regfile/reg_out[1][31] ), .B2(n1931), .C1(
        \regfile/reg_out[12][31] ), .C2(n1932), .A(n2226), .ZN(n2216) );
  OAI22_X1 U3263 ( .A1(n1934), .A2(n1196), .B1(n7017), .B2(n1312), .ZN(n2226)
         );
  AOI222_X1 U3265 ( .A1(\regfile/reg_out[16][31] ), .A2(n1936), .B1(
        \regfile/reg_out[9][31] ), .B2(n1937), .C1(\regfile/reg_out[17][31] ), 
        .C2(n1938), .ZN(n2215) );
  INV_X1 U3266 ( .A(n169), .ZN(n5544) );
  NAND4_X1 U3267 ( .A1(n2227), .A2(n2228), .A3(n2229), .A4(n2230), .ZN(n169)
         );
  NOR4_X1 U3268 ( .A1(n2231), .A2(n2232), .A3(n2233), .A4(n2234), .ZN(n2230)
         );
  NAND3_X1 U3269 ( .A1(n5838), .A2(n5837), .A3(n5839), .ZN(n2234) );
  OAI211_X1 U3270 ( .C1(n5779), .C2(n1325), .A(n5835), .B(n5836), .ZN(n2233)
         );
  OAI222_X1 U3271 ( .A1(n5777), .A2(n1297), .B1(n7025), .B2(n1153), .C1(n5778), 
        .C2(n1181), .ZN(n2232) );
  OAI221_X1 U3272 ( .B1(n7492), .B2(n1353), .C1(n5772), .C2(n1209), .A(n2235), 
        .ZN(n2231) );
  AOI22_X1 U3273 ( .A1(\regfile/reg_out[2][3] ), .A2(n1926), .B1(
        \regfile/reg_out[3][3] ), .B2(n1927), .ZN(n2235) );
  AOI211_X1 U3274 ( .C1(\regfile/reg_out[30][3] ), .C2(n6892), .A(n2236), .B(
        n2237), .ZN(n2229) );
  OAI22_X1 U3275 ( .A1(n7026), .A2(n1239), .B1(n5760), .B2(n1111), .ZN(n2237)
         );
  OAI222_X1 U3278 ( .A1(n5755), .A2(n1125), .B1(n6906), .B2(n1269), .C1(n5759), 
        .C2(n1255), .ZN(n2236) );
  AOI221_X1 U3282 ( .B1(\regfile/reg_out[1][3] ), .B2(n1931), .C1(
        \regfile/reg_out[12][3] ), .C2(n1932), .A(n2238), .ZN(n2228) );
  OAI22_X1 U3283 ( .A1(n1934), .A2(n1195), .B1(n7017), .B2(n1311), .ZN(n2238)
         );
  AOI222_X1 U3285 ( .A1(\regfile/reg_out[16][3] ), .A2(n1936), .B1(
        \regfile/reg_out[9][3] ), .B2(n1937), .C1(\regfile/reg_out[17][3] ), 
        .C2(n1938), .ZN(n2227) );
  INV_X1 U3286 ( .A(n165), .ZN(n5541) );
  NAND4_X1 U3287 ( .A1(n2239), .A2(n2240), .A3(n2241), .A4(n2242), .ZN(n165)
         );
  NOR4_X1 U3288 ( .A1(n2243), .A2(n2244), .A3(n2245), .A4(n2246), .ZN(n2242)
         );
  NAND3_X1 U3289 ( .A1(n5828), .A2(n5827), .A3(n5829), .ZN(n2246) );
  OAI211_X1 U3290 ( .C1(n5779), .C2(n1324), .A(n5825), .B(n5826), .ZN(n2245)
         );
  OAI222_X1 U3291 ( .A1(n5777), .A2(n1296), .B1(n7025), .B2(n1152), .C1(n5778), 
        .C2(n1180), .ZN(n2244) );
  OAI221_X1 U3292 ( .B1(n7491), .B2(n1352), .C1(n5772), .C2(n1208), .A(n2247), 
        .ZN(n2243) );
  AOI22_X1 U3293 ( .A1(\regfile/reg_out[2][4] ), .A2(n1926), .B1(
        \regfile/reg_out[3][4] ), .B2(n1927), .ZN(n2247) );
  AOI211_X1 U3294 ( .C1(\regfile/reg_out[30][4] ), .C2(n6892), .A(n2248), .B(
        n2249), .ZN(n2241) );
  OAI22_X1 U3295 ( .A1(n7026), .A2(n1238), .B1(n5760), .B2(n1110), .ZN(n2249)
         );
  OAI222_X1 U3298 ( .A1(n5755), .A2(n1124), .B1(n6906), .B2(n1268), .C1(n5759), 
        .C2(n1254), .ZN(n2248) );
  AOI221_X1 U3302 ( .B1(\regfile/reg_out[1][4] ), .B2(n1931), .C1(
        \regfile/reg_out[12][4] ), .C2(n1932), .A(n2250), .ZN(n2240) );
  OAI22_X1 U3303 ( .A1(n1934), .A2(n1194), .B1(n7017), .B2(n1310), .ZN(n2250)
         );
  AOI222_X1 U3305 ( .A1(\regfile/reg_out[16][4] ), .A2(n1936), .B1(
        \regfile/reg_out[9][4] ), .B2(n1937), .C1(\regfile/reg_out[17][4] ), 
        .C2(n1938), .ZN(n2239) );
  INV_X1 U3306 ( .A(n161), .ZN(n5538) );
  NAND4_X1 U3307 ( .A1(n2251), .A2(n2252), .A3(n2253), .A4(n2254), .ZN(n161)
         );
  NOR4_X1 U3308 ( .A1(n2255), .A2(n2256), .A3(n2257), .A4(n2258), .ZN(n2254)
         );
  NAND3_X1 U3309 ( .A1(n5818), .A2(n5817), .A3(n5819), .ZN(n2258) );
  OAI211_X1 U3310 ( .C1(n5779), .C2(n891), .A(n5815), .B(n5816), .ZN(n2257) );
  OAI222_X1 U3311 ( .A1(n5777), .A2(n895), .B1(n7025), .B2(n894), .C1(n5778), 
        .C2(n890), .ZN(n2256) );
  OAI221_X1 U3312 ( .B1(n7492), .B2(n908), .C1(n5772), .C2(n907), .A(n2259), 
        .ZN(n2255) );
  AOI22_X1 U3313 ( .A1(\regfile/reg_out[2][5] ), .A2(n1926), .B1(
        \regfile/reg_out[3][5] ), .B2(n1927), .ZN(n2259) );
  AOI211_X1 U3314 ( .C1(\regfile/reg_out[30][5] ), .C2(n6892), .A(n2260), .B(
        n2261), .ZN(n2253) );
  OAI22_X1 U3315 ( .A1(n7026), .A2(n905), .B1(n5760), .B2(n901), .ZN(n2261) );
  OAI222_X1 U3318 ( .A1(n5755), .A2(n899), .B1(n6906), .B2(n900), .C1(n5759), 
        .C2(n902), .ZN(n2260) );
  AOI221_X1 U3322 ( .B1(\regfile/reg_out[1][5] ), .B2(n1931), .C1(
        \regfile/reg_out[12][5] ), .C2(n1932), .A(n2262), .ZN(n2252) );
  OAI22_X1 U3323 ( .A1(n1934), .A2(n909), .B1(n7017), .B2(n893), .ZN(n2262) );
  AOI222_X1 U3325 ( .A1(\regfile/reg_out[16][5] ), .A2(n1936), .B1(
        \regfile/reg_out[9][5] ), .B2(n1937), .C1(\regfile/reg_out[17][5] ), 
        .C2(n1938), .ZN(n2251) );
  INV_X1 U3326 ( .A(n157), .ZN(n5535) );
  NAND4_X1 U3327 ( .A1(n2263), .A2(n2264), .A3(n2265), .A4(n2266), .ZN(n157)
         );
  NOR4_X1 U3328 ( .A1(n2267), .A2(n2268), .A3(n2269), .A4(n2270), .ZN(n2266)
         );
  NAND3_X1 U3329 ( .A1(n5808), .A2(n5807), .A3(n5809), .ZN(n2270) );
  OAI211_X1 U3330 ( .C1(n5779), .C2(n935), .A(n5805), .B(n5806), .ZN(n2269) );
  OAI222_X1 U3331 ( .A1(n5777), .A2(n939), .B1(n7025), .B2(n938), .C1(n5778), 
        .C2(n934), .ZN(n2268) );
  OAI221_X1 U3332 ( .B1(n7493), .B2(n952), .C1(n5772), .C2(n951), .A(n2271), 
        .ZN(n2267) );
  AOI22_X1 U3333 ( .A1(\regfile/reg_out[2][6] ), .A2(n1926), .B1(
        \regfile/reg_out[3][6] ), .B2(n1927), .ZN(n2271) );
  AOI211_X1 U3334 ( .C1(\regfile/reg_out[30][6] ), .C2(n6892), .A(n2272), .B(
        n2273), .ZN(n2265) );
  OAI22_X1 U3335 ( .A1(n7026), .A2(n949), .B1(n5760), .B2(n945), .ZN(n2273) );
  OAI222_X1 U3338 ( .A1(n5755), .A2(n943), .B1(n6906), .B2(n944), .C1(n5759), 
        .C2(n946), .ZN(n2272) );
  AOI221_X1 U3342 ( .B1(\regfile/reg_out[1][6] ), .B2(n1931), .C1(
        \regfile/reg_out[12][6] ), .C2(n1932), .A(n2274), .ZN(n2264) );
  OAI22_X1 U3343 ( .A1(n1934), .A2(n953), .B1(n7017), .B2(n937), .ZN(n2274) );
  AOI222_X1 U3345 ( .A1(\regfile/reg_out[16][6] ), .A2(n1936), .B1(
        \regfile/reg_out[9][6] ), .B2(n1937), .C1(\regfile/reg_out[17][6] ), 
        .C2(n1938), .ZN(n2263) );
  INV_X1 U3346 ( .A(n153), .ZN(n5532) );
  NAND4_X1 U3347 ( .A1(n2275), .A2(n2276), .A3(n2277), .A4(n2278), .ZN(n153)
         );
  NOR4_X1 U3348 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2278)
         );
  NAND3_X1 U3349 ( .A1(n5796), .A2(n5795), .A3(n5797), .ZN(n2282) );
  OAI211_X1 U3350 ( .C1(n5779), .C2(n974), .A(n5793), .B(n5794), .ZN(n2281) );
  OAI222_X1 U3351 ( .A1(n5777), .A2(n978), .B1(n7025), .B2(n977), .C1(n5778), 
        .C2(n973), .ZN(n2280) );
  OAI221_X1 U3352 ( .B1(n7493), .B2(n991), .C1(n5772), .C2(n990), .A(n2283), 
        .ZN(n2279) );
  AOI22_X1 U3353 ( .A1(\regfile/reg_out[2][7] ), .A2(n1926), .B1(
        \regfile/reg_out[3][7] ), .B2(n1927), .ZN(n2283) );
  AOI211_X1 U3354 ( .C1(\regfile/reg_out[30][7] ), .C2(n1928), .A(n2284), .B(
        n2285), .ZN(n2277) );
  OAI22_X1 U3355 ( .A1(n7026), .A2(n988), .B1(n5760), .B2(n984), .ZN(n2285) );
  OAI222_X1 U3358 ( .A1(n5755), .A2(n982), .B1(n6906), .B2(n983), .C1(n5759), 
        .C2(n985), .ZN(n2284) );
  AOI221_X1 U3362 ( .B1(\regfile/reg_out[1][7] ), .B2(n1931), .C1(
        \regfile/reg_out[12][7] ), .C2(n1932), .A(n2286), .ZN(n2276) );
  OAI22_X1 U3363 ( .A1(n1934), .A2(n992), .B1(n7017), .B2(n976), .ZN(n2286) );
  AOI222_X1 U3365 ( .A1(\regfile/reg_out[16][7] ), .A2(n1936), .B1(
        \regfile/reg_out[9][7] ), .B2(n1937), .C1(\regfile/reg_out[17][7] ), 
        .C2(n1938), .ZN(n2275) );
  INV_X1 U3366 ( .A(n149), .ZN(n5529) );
  NAND4_X1 U3367 ( .A1(n2287), .A2(n2288), .A3(n2289), .A4(n2290), .ZN(n149)
         );
  NOR4_X1 U3368 ( .A1(n2291), .A2(n2292), .A3(n2293), .A4(n2294), .ZN(n2290)
         );
  NAND3_X1 U3369 ( .A1(n5783), .A2(n5782), .A3(n5784), .ZN(n2294) );
  OAI211_X1 U3370 ( .C1(n5779), .C2(n1323), .A(n5780), .B(n5781), .ZN(n2293)
         );
  OAI222_X1 U3371 ( .A1(n5777), .A2(n1295), .B1(n7025), .B2(n1151), .C1(n5778), 
        .C2(n1179), .ZN(n2292) );
  OAI221_X1 U3372 ( .B1(n7493), .B2(n1351), .C1(n5772), .C2(n1207), .A(n2295), 
        .ZN(n2291) );
  AOI22_X1 U3373 ( .A1(\regfile/reg_out[2][8] ), .A2(n1926), .B1(
        \regfile/reg_out[3][8] ), .B2(n1927), .ZN(n2295) );
  AOI211_X1 U3374 ( .C1(\regfile/reg_out[30][8] ), .C2(n1928), .A(n2296), .B(
        n2297), .ZN(n2289) );
  OAI22_X1 U3375 ( .A1(n7026), .A2(n1237), .B1(n5760), .B2(n1109), .ZN(n2297)
         );
  OAI222_X1 U3378 ( .A1(n5755), .A2(n1123), .B1(n6906), .B2(n1267), .C1(n5759), 
        .C2(n1253), .ZN(n2296) );
  AOI221_X1 U3382 ( .B1(\regfile/reg_out[1][8] ), .B2(n1931), .C1(
        \regfile/reg_out[12][8] ), .C2(n1932), .A(n2298), .ZN(n2288) );
  OAI22_X1 U3383 ( .A1(n1934), .A2(n1193), .B1(n7017), .B2(n1309), .ZN(n2298)
         );
  AOI222_X1 U3385 ( .A1(\regfile/reg_out[16][8] ), .A2(n1936), .B1(
        \regfile/reg_out[9][8] ), .B2(n1937), .C1(\regfile/reg_out[17][8] ), 
        .C2(n1938), .ZN(n2287) );
  INV_X1 U3386 ( .A(n145), .ZN(n5524) );
  NAND4_X1 U3387 ( .A1(n2299), .A2(n2300), .A3(n2301), .A4(n2302), .ZN(n145)
         );
  NOR4_X1 U3388 ( .A1(n2303), .A2(n2304), .A3(n2305), .A4(n2306), .ZN(n2302)
         );
  NAND3_X1 U3389 ( .A1(n5766), .A2(n5761), .A3(n5773), .ZN(n2306) );
  OAI211_X1 U3390 ( .C1(n5779), .C2(n1013), .A(n5751), .B(n5756), .ZN(n2305)
         );
  OAI222_X1 U3391 ( .A1(n5777), .A2(n1017), .B1(n7025), .B2(n1016), .C1(n5778), 
        .C2(n1012), .ZN(n2304) );
  OAI221_X1 U3392 ( .B1(n7493), .B2(n1030), .C1(n5772), .C2(n1029), .A(n2307), 
        .ZN(n2303) );
  AOI22_X1 U3393 ( .A1(\regfile/reg_out[2][9] ), .A2(n1926), .B1(
        \regfile/reg_out[3][9] ), .B2(n1927), .ZN(n2307) );
  AOI211_X1 U3396 ( .C1(\regfile/reg_out[30][9] ), .C2(n1928), .A(n2308), .B(
        n2309), .ZN(n2301) );
  OAI22_X1 U3397 ( .A1(n7026), .A2(n1027), .B1(n5760), .B2(n1023), .ZN(n2309)
         );
  OAI222_X1 U3400 ( .A1(n5755), .A2(n1021), .B1(n6906), .B2(n1022), .C1(n5759), 
        .C2(n1024), .ZN(n2308) );
  INV_X1 U3404 ( .A(n5765), .ZN(n1928) );
  AOI221_X1 U3405 ( .B1(\regfile/reg_out[1][9] ), .B2(n1931), .C1(
        \regfile/reg_out[12][9] ), .C2(n1932), .A(n2310), .ZN(n2300) );
  OAI22_X1 U3406 ( .A1(n1934), .A2(n1031), .B1(n7017), .B2(n1015), .ZN(n2310)
         );
  NAND3_X1 U3408 ( .A1(n6025), .A2(rs2_addr[3]), .A3(n6037), .ZN(n1935) );
  INV_X1 U3410 ( .A(rs2_addr[0]), .ZN(n2311) );
  INV_X1 U3412 ( .A(rs2_addr[4]), .ZN(n2312) );
  AOI222_X1 U3414 ( .A1(\regfile/reg_out[16][9] ), .A2(n1936), .B1(
        \regfile/reg_out[9][9] ), .B2(n1937), .C1(\regfile/reg_out[17][9] ), 
        .C2(n1938), .ZN(n2299) );
  INV_X1 U3418 ( .A(n1667), .ZN(n5514) );
  NAND4_X1 U3419 ( .A1(n2313), .A2(n2314), .A3(n2315), .A4(n2316), .ZN(n1667)
         );
  NOR4_X1 U3420 ( .A1(n2317), .A2(n2318), .A3(n2319), .A4(n2320), .ZN(n2316)
         );
  NAND3_X1 U3421 ( .A1(n5711), .A2(n5710), .A3(n5712), .ZN(n2320) );
  OAI211_X1 U3422 ( .C1(n5654), .C2(n1336), .A(n5708), .B(n5709), .ZN(n2319)
         );
  OAI222_X1 U3424 ( .A1(n5652), .A2(n1308), .B1(n7518), .B2(n1164), .C1(n7482), 
        .C2(n1192), .ZN(n2318) );
  OAI221_X1 U3428 ( .B1(n5646), .B2(n1364), .C1(n5647), .C2(n1220), .A(n2321), 
        .ZN(n2317) );
  AOI22_X1 U3429 ( .A1(\regfile/reg_out[2][0] ), .A2(n7641), .B1(
        \regfile/reg_out[3][0] ), .B2(n2323), .ZN(n2321) );
  AOI211_X1 U3432 ( .C1(\regfile/reg_out[16][0] ), .C2(n2324), .A(n2325), .B(
        n2326), .ZN(n2315) );
  OAI22_X1 U3433 ( .A1(n5624), .A2(n1294), .B1(n1350), .B2(n2327), .ZN(n2326)
         );
  OAI221_X1 U3436 ( .B1(n1410), .B2(n2328), .C1(n1206), .C2(n2329), .A(n2330), 
        .ZN(n2325) );
  AOI22_X1 U3437 ( .A1(n2331), .A2(\regfile/reg_out[12][0] ), .B1(n2332), .B2(
        \regfile/reg_out[13][0] ), .ZN(n2330) );
  AOI222_X1 U3440 ( .A1(\regfile/reg_out[27][0] ), .A2(n2333), .B1(
        \regfile/reg_out[23][0] ), .B2(n2334), .C1(\regfile/reg_out[22][0] ), 
        .C2(n2335), .ZN(n2314) );
  AOI222_X1 U3441 ( .A1(\regfile/reg_out[30][0] ), .A2(n2336), .B1(
        \regfile/reg_out[26][0] ), .B2(n2337), .C1(\regfile/reg_out[31][0] ), 
        .C2(n2338), .ZN(n2313) );
  INV_X1 U3442 ( .A(n335), .ZN(n5513) );
  NAND4_X1 U3443 ( .A1(n2339), .A2(n2340), .A3(n2341), .A4(n2342), .ZN(n335)
         );
  NAND3_X1 U3445 ( .A1(n5703), .A2(n5702), .A3(n5704), .ZN(n2346) );
  OAI211_X1 U3446 ( .C1(n5654), .C2(n337), .A(n5700), .B(n5701), .ZN(n2345) );
  OAI222_X1 U3448 ( .A1(n5652), .A2(n341), .B1(n7519), .B2(n340), .C1(n7484), 
        .C2(n336), .ZN(n2344) );
  OAI221_X1 U3452 ( .B1(n5646), .B2(n354), .C1(n5647), .C2(n353), .A(n2347), 
        .ZN(n2343) );
  AOI22_X1 U3453 ( .A1(\regfile/reg_out[2][24] ), .A2(n7641), .B1(
        \regfile/reg_out[3][24] ), .B2(n2323), .ZN(n2347) );
  AOI211_X1 U3456 ( .C1(\regfile/reg_out[16][24] ), .C2(n2324), .A(n2348), .B(
        n2349), .ZN(n2341) );
  OAI22_X1 U3457 ( .A1(n5624), .A2(n343), .B1(n356), .B2(n2327), .ZN(n2349) );
  OAI221_X1 U3460 ( .B1(n344), .B2(n2328), .C1(n355), .C2(n2329), .A(n2350), 
        .ZN(n2348) );
  AOI22_X1 U3461 ( .A1(n2331), .A2(\regfile/reg_out[12][24] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][24] ), .ZN(n2350) );
  AOI222_X1 U3464 ( .A1(\regfile/reg_out[27][24] ), .A2(n2333), .B1(
        \regfile/reg_out[23][24] ), .B2(n2334), .C1(\regfile/reg_out[22][24] ), 
        .C2(n2335), .ZN(n2340) );
  AOI222_X1 U3465 ( .A1(\regfile/reg_out[30][24] ), .A2(n2336), .B1(
        \regfile/reg_out[26][24] ), .B2(n2337), .C1(\regfile/reg_out[31][24] ), 
        .C2(n2338), .ZN(n2339) );
  INV_X1 U3466 ( .A(n236), .ZN(n5512) );
  NAND4_X1 U3467 ( .A1(n2351), .A2(n2352), .A3(n2353), .A4(n2354), .ZN(n236)
         );
  NAND3_X1 U3469 ( .A1(n5695), .A2(n5694), .A3(n5696), .ZN(n2358) );
  OAI211_X1 U3470 ( .C1(n5654), .C2(n241), .A(n5692), .B(n5693), .ZN(n2357) );
  OAI222_X1 U3472 ( .A1(n5652), .A2(n253), .B1(n7519), .B2(n250), .C1(n7483), 
        .C2(n238), .ZN(n2356) );
  OAI221_X1 U3476 ( .B1(n5646), .B2(n312), .C1(n5647), .C2(n309), .A(n2359), 
        .ZN(n2355) );
  AOI22_X1 U3477 ( .A1(\regfile/reg_out[2][25] ), .A2(n7642), .B1(
        \regfile/reg_out[3][25] ), .B2(n2323), .ZN(n2359) );
  AOI211_X1 U3480 ( .C1(\regfile/reg_out[16][25] ), .C2(n2324), .A(n2360), .B(
        n2361), .ZN(n2353) );
  OAI22_X1 U3481 ( .A1(n5624), .A2(n259), .B1(n318), .B2(n2327), .ZN(n2361) );
  OAI221_X1 U3484 ( .B1(n266), .B2(n2328), .C1(n315), .C2(n2329), .A(n2362), 
        .ZN(n2360) );
  AOI22_X1 U3485 ( .A1(n2331), .A2(\regfile/reg_out[12][25] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][25] ), .ZN(n2362) );
  AOI222_X1 U3488 ( .A1(\regfile/reg_out[27][25] ), .A2(n2333), .B1(
        \regfile/reg_out[23][25] ), .B2(n2334), .C1(\regfile/reg_out[22][25] ), 
        .C2(n2335), .ZN(n2352) );
  AOI222_X1 U3489 ( .A1(\regfile/reg_out[30][25] ), .A2(n2336), .B1(
        \regfile/reg_out[26][25] ), .B2(n2337), .C1(\regfile/reg_out[31][25] ), 
        .C2(n2338), .ZN(n2351) );
  INV_X1 U3490 ( .A(n1614), .ZN(n5511) );
  NAND4_X1 U3491 ( .A1(n2363), .A2(n2364), .A3(n2365), .A4(n2366), .ZN(n1614)
         );
  NOR4_X1 U3492 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(n2366)
         );
  NAND3_X1 U3493 ( .A1(n5687), .A2(n5686), .A3(n5688), .ZN(n2370) );
  OAI211_X1 U3494 ( .C1(n5654), .C2(n1332), .A(n5684), .B(n5685), .ZN(n2369)
         );
  OAI222_X1 U3496 ( .A1(n5652), .A2(n1304), .B1(n7518), .B2(n1160), .C1(n7484), 
        .C2(n1188), .ZN(n2368) );
  OAI221_X1 U3500 ( .B1(n5646), .B2(n1360), .C1(n5647), .C2(n1216), .A(n2371), 
        .ZN(n2367) );
  AOI22_X1 U3501 ( .A1(\regfile/reg_out[2][26] ), .A2(n7642), .B1(
        \regfile/reg_out[3][26] ), .B2(n2323), .ZN(n2371) );
  AOI211_X1 U3504 ( .C1(\regfile/reg_out[16][26] ), .C2(n2324), .A(n2372), .B(
        n2373), .ZN(n2365) );
  OAI22_X1 U3505 ( .A1(n5624), .A2(n1290), .B1(n1346), .B2(n2327), .ZN(n2373)
         );
  OAI221_X1 U3508 ( .B1(n1402), .B2(n2328), .C1(n1202), .C2(n2329), .A(n2374), 
        .ZN(n2372) );
  AOI22_X1 U3509 ( .A1(n2331), .A2(\regfile/reg_out[12][26] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][26] ), .ZN(n2374) );
  AOI222_X1 U3512 ( .A1(\regfile/reg_out[27][26] ), .A2(n2333), .B1(
        \regfile/reg_out[23][26] ), .B2(n2334), .C1(\regfile/reg_out[22][26] ), 
        .C2(n2335), .ZN(n2364) );
  AOI222_X1 U3513 ( .A1(\regfile/reg_out[30][26] ), .A2(n2336), .B1(
        \regfile/reg_out[26][26] ), .B2(n2337), .C1(\regfile/reg_out[31][26] ), 
        .C2(n2338), .ZN(n2363) );
  INV_X1 U3514 ( .A(n1616), .ZN(n5510) );
  NAND4_X1 U3515 ( .A1(n2375), .A2(n2376), .A3(n2377), .A4(n2378), .ZN(n1616)
         );
  NOR4_X1 U3516 ( .A1(n2379), .A2(n2380), .A3(n2381), .A4(n2382), .ZN(n2378)
         );
  NAND3_X1 U3517 ( .A1(n5679), .A2(n5678), .A3(n5680), .ZN(n2382) );
  OAI211_X1 U3518 ( .C1(n5654), .C2(n1331), .A(n5676), .B(n5677), .ZN(n2381)
         );
  OAI222_X1 U3520 ( .A1(n5652), .A2(n1303), .B1(n7518), .B2(n1159), .C1(n7484), 
        .C2(n1187), .ZN(n2380) );
  OAI221_X1 U3524 ( .B1(n5646), .B2(n1359), .C1(n5647), .C2(n1215), .A(n2383), 
        .ZN(n2379) );
  AOI22_X1 U3525 ( .A1(\regfile/reg_out[2][27] ), .A2(n7641), .B1(
        \regfile/reg_out[3][27] ), .B2(n2323), .ZN(n2383) );
  AOI211_X1 U3528 ( .C1(\regfile/reg_out[16][27] ), .C2(n2324), .A(n2384), .B(
        n2385), .ZN(n2377) );
  OAI22_X1 U3529 ( .A1(n5624), .A2(n1289), .B1(n1345), .B2(n2327), .ZN(n2385)
         );
  OAI221_X1 U3532 ( .B1(n1401), .B2(n2328), .C1(n1201), .C2(n2329), .A(n2386), 
        .ZN(n2384) );
  AOI22_X1 U3533 ( .A1(n2331), .A2(\regfile/reg_out[12][27] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][27] ), .ZN(n2386) );
  AOI222_X1 U3536 ( .A1(\regfile/reg_out[27][27] ), .A2(n2333), .B1(
        \regfile/reg_out[23][27] ), .B2(n2334), .C1(\regfile/reg_out[22][27] ), 
        .C2(n2335), .ZN(n2376) );
  AOI222_X1 U3537 ( .A1(\regfile/reg_out[30][27] ), .A2(n2336), .B1(
        \regfile/reg_out[26][27] ), .B2(n2337), .C1(\regfile/reg_out[31][27] ), 
        .C2(n2338), .ZN(n2375) );
  INV_X1 U3538 ( .A(n1618), .ZN(n5509) );
  NAND4_X1 U3539 ( .A1(n2387), .A2(n2388), .A3(n2389), .A4(n2390), .ZN(n1618)
         );
  NOR4_X1 U3540 ( .A1(n2391), .A2(n2392), .A3(n2393), .A4(n2394), .ZN(n2390)
         );
  NAND3_X1 U3541 ( .A1(n5671), .A2(n5670), .A3(n5672), .ZN(n2394) );
  OAI211_X1 U3542 ( .C1(n5654), .C2(n1330), .A(n5668), .B(n5669), .ZN(n2393)
         );
  OAI222_X1 U3544 ( .A1(n5652), .A2(n1302), .B1(n7519), .B2(n1158), .C1(n7484), 
        .C2(n1186), .ZN(n2392) );
  OAI221_X1 U3548 ( .B1(n5646), .B2(n1358), .C1(n5647), .C2(n1214), .A(n2395), 
        .ZN(n2391) );
  AOI22_X1 U3549 ( .A1(\regfile/reg_out[2][28] ), .A2(n7642), .B1(
        \regfile/reg_out[3][28] ), .B2(n2323), .ZN(n2395) );
  AOI211_X1 U3552 ( .C1(\regfile/reg_out[16][28] ), .C2(n2324), .A(n2396), .B(
        n2397), .ZN(n2389) );
  OAI22_X1 U3553 ( .A1(n5624), .A2(n1288), .B1(n1344), .B2(n2327), .ZN(n2397)
         );
  OAI221_X1 U3556 ( .B1(n1400), .B2(n2328), .C1(n1200), .C2(n2329), .A(n2398), 
        .ZN(n2396) );
  AOI22_X1 U3557 ( .A1(n2331), .A2(\regfile/reg_out[12][28] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][28] ), .ZN(n2398) );
  AOI222_X1 U3560 ( .A1(\regfile/reg_out[27][28] ), .A2(n2333), .B1(
        \regfile/reg_out[23][28] ), .B2(n2334), .C1(\regfile/reg_out[22][28] ), 
        .C2(n2335), .ZN(n2388) );
  AOI222_X1 U3561 ( .A1(\regfile/reg_out[30][28] ), .A2(n2336), .B1(
        \regfile/reg_out[26][28] ), .B2(n2337), .C1(\regfile/reg_out[31][28] ), 
        .C2(n2338), .ZN(n2387) );
  INV_X1 U3562 ( .A(n1620), .ZN(n5508) );
  NAND4_X1 U3563 ( .A1(n2399), .A2(n2400), .A3(n2401), .A4(n2402), .ZN(n1620)
         );
  NOR4_X1 U3564 ( .A1(n2403), .A2(n2404), .A3(n2405), .A4(n2406), .ZN(n2402)
         );
  NAND3_X1 U3565 ( .A1(n5663), .A2(n5662), .A3(n5664), .ZN(n2406) );
  OAI211_X1 U3566 ( .C1(n5654), .C2(n1329), .A(n5660), .B(n5661), .ZN(n2405)
         );
  OAI222_X1 U3568 ( .A1(n5652), .A2(n1301), .B1(n7519), .B2(n1157), .C1(n7484), 
        .C2(n1185), .ZN(n2404) );
  OAI221_X1 U3572 ( .B1(n5646), .B2(n1357), .C1(n5647), .C2(n1213), .A(n2407), 
        .ZN(n2403) );
  AOI22_X1 U3573 ( .A1(\regfile/reg_out[2][29] ), .A2(n7641), .B1(
        \regfile/reg_out[3][29] ), .B2(n2323), .ZN(n2407) );
  AOI211_X1 U3576 ( .C1(\regfile/reg_out[16][29] ), .C2(n2324), .A(n2408), .B(
        n2409), .ZN(n2401) );
  OAI22_X1 U3577 ( .A1(n5624), .A2(n1287), .B1(n1343), .B2(n2327), .ZN(n2409)
         );
  OAI221_X1 U3580 ( .B1(n1399), .B2(n2328), .C1(n1199), .C2(n2329), .A(n2410), 
        .ZN(n2408) );
  AOI22_X1 U3581 ( .A1(n2331), .A2(\regfile/reg_out[12][29] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][29] ), .ZN(n2410) );
  AOI222_X1 U3584 ( .A1(\regfile/reg_out[27][29] ), .A2(n2333), .B1(
        \regfile/reg_out[23][29] ), .B2(n2334), .C1(\regfile/reg_out[22][29] ), 
        .C2(n2335), .ZN(n2400) );
  AOI222_X1 U3585 ( .A1(\regfile/reg_out[30][29] ), .A2(n2336), .B1(
        \regfile/reg_out[26][29] ), .B2(n2337), .C1(\regfile/reg_out[31][29] ), 
        .C2(n2338), .ZN(n2399) );
  INV_X1 U3586 ( .A(n1622), .ZN(n5507) );
  NAND4_X1 U3587 ( .A1(n2414), .A2(n2412), .A3(n2413), .A4(n2411), .ZN(n1622)
         );
  NAND3_X1 U3589 ( .A1(n5641), .A2(n5636), .A3(n5648), .ZN(n2418) );
  OAI211_X1 U3590 ( .C1(n5654), .C2(n1327), .A(n5626), .B(n5631), .ZN(n2417)
         );
  OAI222_X1 U3592 ( .A1(n5652), .A2(n1299), .B1(n7517), .B2(n1155), .C1(n7483), 
        .C2(n1183), .ZN(n2416) );
  OAI221_X1 U3596 ( .B1(n5646), .B2(n1355), .C1(n5647), .C2(n1211), .A(n2419), 
        .ZN(n2415) );
  AOI22_X1 U3597 ( .A1(\regfile/reg_out[2][30] ), .A2(n7641), .B1(
        \regfile/reg_out[3][30] ), .B2(n2323), .ZN(n2419) );
  AOI211_X1 U3600 ( .C1(\regfile/reg_out[16][30] ), .C2(n2324), .A(n2420), .B(
        n2421), .ZN(n2413) );
  OAI22_X1 U3601 ( .A1(n5624), .A2(n1285), .B1(n1341), .B2(n2327), .ZN(n2421)
         );
  OAI221_X1 U3604 ( .B1(n1391), .B2(n2328), .C1(n1197), .C2(n2329), .A(n2422), 
        .ZN(n2420) );
  AOI22_X1 U3605 ( .A1(n2331), .A2(\regfile/reg_out[12][30] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][30] ), .ZN(n2422) );
  AOI222_X1 U3608 ( .A1(\regfile/reg_out[27][30] ), .A2(n2333), .B1(
        \regfile/reg_out[23][30] ), .B2(n2334), .C1(\regfile/reg_out[22][30] ), 
        .C2(n2335), .ZN(n2412) );
  AOI222_X1 U3609 ( .A1(\regfile/reg_out[30][30] ), .A2(n2336), .B1(
        \regfile/reg_out[26][30] ), .B2(n2337), .C1(\regfile/reg_out[31][30] ), 
        .C2(n2338), .ZN(n2411) );
  INV_X1 U3610 ( .A(n1086), .ZN(n5506) );
  NAND4_X1 U3611 ( .A1(n2426), .A2(n2424), .A3(n2425), .A4(n2423), .ZN(n1086)
         );
  NAND3_X1 U3613 ( .A1(n6427), .A2(n6423), .A3(n6432), .ZN(n2430) );
  OAI211_X1 U3614 ( .C1(n5654), .C2(n1326), .A(n6412), .B(n6419), .ZN(n2429)
         );
  OAI222_X1 U3616 ( .A1(n5652), .A2(n1298), .B1(n7517), .B2(n1154), .C1(n7483), 
        .C2(n1182), .ZN(n2428) );
  AOI22_X1 U3621 ( .A1(\regfile/reg_out[2][31] ), .A2(n7642), .B1(
        \regfile/reg_out[3][31] ), .B2(n2323), .ZN(n2431) );
  OAI22_X1 U3625 ( .A1(n5624), .A2(n1284), .B1(n1340), .B2(n2327), .ZN(n2433)
         );
  OAI221_X1 U3628 ( .B1(n1389), .B2(n2328), .C1(n1196), .C2(n2329), .A(n2434), 
        .ZN(n2432) );
  AOI22_X1 U3629 ( .A1(n2331), .A2(\regfile/reg_out[12][31] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][31] ), .ZN(n2434) );
  AOI222_X1 U3632 ( .A1(\regfile/reg_out[27][31] ), .A2(n2333), .B1(
        \regfile/reg_out[23][31] ), .B2(n2334), .C1(\regfile/reg_out[22][31] ), 
        .C2(n2335), .ZN(n2424) );
  AOI222_X1 U3633 ( .A1(\regfile/reg_out[30][31] ), .A2(n2336), .B1(
        \regfile/reg_out[26][31] ), .B2(n2337), .C1(\regfile/reg_out[31][31] ), 
        .C2(n2338), .ZN(n2423) );
  INV_X1 U3634 ( .A(\x_mem_command[MB] ), .ZN(n5505) );
  NAND2_X1 U3635 ( .A1(n1546), .A2(n1519), .ZN(\x_mem_command[MB] ) );
  AOI21_X1 U3637 ( .B1(\Scc_coproc/cause[4] ), .B2(serve_exception), .A(n1596), 
        .ZN(n4510) );
  NAND2_X1 U3638 ( .A1(n2435), .A2(n2436), .ZN(n1596) );
  NAND3_X1 U3639 ( .A1(\Scc_coproc/x_exc_word[4] ), .A2(n1585), .A3(n883), 
        .ZN(n2436) );
  AOI21_X1 U3640 ( .B1(\Scc_coproc/cause[5] ), .B2(serve_exception), .A(n1038), 
        .ZN(n4509) );
  NAND2_X1 U3641 ( .A1(n2435), .A2(n2437), .ZN(n1038) );
  NAND3_X1 U3642 ( .A1(n7130), .A2(n1585), .A3(n883), .ZN(n2437) );
  NOR2_X1 U3643 ( .A1(n1610), .A2(n7163), .ZN(n883) );
  INV_X1 U3644 ( .A(\Scc_coproc/interrupt_active ), .ZN(n1610) );
  INV_X1 U3645 ( .A(n5740), .ZN(n1585) );
  NAND3_X1 U3646 ( .A1(n1591), .A2(n1590), .A3(n1587), .ZN(n2435) );
  NOR4_X1 U3647 ( .A1(\Scc_coproc/interrupt[3] ), .A2(n5740), .A3(n1579), .A4(
        n2438), .ZN(n1587) );
  NAND2_X1 U3648 ( .A1(n6492), .A2(n1581), .ZN(n2438) );
  NOR4_X1 U3649 ( .A1(\Scc_coproc/interrupt[4] ), .A2(
        \Scc_coproc/interrupt[5] ), .A3(\Scc_coproc/interrupt[6] ), .A4(
        \Scc_coproc/interrupt[7] ), .ZN(n1581) );
  INV_X1 U3650 ( .A(\Scc_coproc/N551 ), .ZN(n1579) );
  INV_X1 U3652 ( .A(\x_mem_command[MH] ), .ZN(n4508) );
  NAND2_X1 U3653 ( .A1(n1546), .A2(n1526), .ZN(\x_mem_command[MH] ) );
  INV_X1 U3655 ( .A(\x_mem_command[MR] ), .ZN(n4507) );
  NAND2_X1 U3656 ( .A1(n1546), .A2(n1530), .ZN(\x_mem_command[MR] ) );
  AOI22_X1 U3660 ( .A1(\Mpath/the_alu/diff[1] ), .A2(n1698), .B1(
        \Mpath/the_alu/sum[1] ), .B2(n7634), .ZN(n2440) );
  INV_X1 U3662 ( .A(\Mpath/the_alu/N82 ), .ZN(n2443) );
  OAI221_X1 U3663 ( .B1(\Mpath/the_alu/N81 ), .B2(n1693), .C1(n1841), .C2(
        n2444), .A(n1694), .ZN(n2442) );
  OAI22_X1 U3665 ( .A1(n7186), .A2(n2444), .B1(\Mpath/the_alu/N81 ), .B2(n1841), .ZN(n2441) );
  INV_X1 U3667 ( .A(\Mpath/the_alu/N486 ), .ZN(n2445) );
  INV_X1 U3668 ( .A(\Mpath/the_alu/N81 ), .ZN(n2444) );
  NAND2_X1 U3677 ( .A1(n2449), .A2(n2450), .ZN(daddr_out[0]) );
  AND2_X1 U3681 ( .A1(\Mpath/the_alu/N503 ), .A2(\Mpath/the_alu/N498 ), .ZN(
        n2454) );
  INV_X1 U3683 ( .A(n2452), .ZN(n2456) );
  AOI22_X1 U3684 ( .A1(\Mpath/the_alu/sum[0] ), .A2(n7634), .B1(n6504), .B2(
        n6499), .ZN(n2449) );
  INV_X1 U3689 ( .A(\Mpath/the_alu/N468 ), .ZN(n2457) );
  INV_X1 U3690 ( .A(\Mcontrol/st_logic/N42 ), .ZN(byp_controlB[0]) );
  INV_X1 U3701 ( .A(n1078), .ZN(n2464) );
  NAND4_X1 U3702 ( .A1(n2465), .A2(n2466), .A3(n2467), .A4(n2468), .ZN(n1078)
         );
  NOR4_X1 U3703 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(n2468)
         );
  NAND3_X1 U3704 ( .A1(n6084), .A2(n6083), .A3(n6085), .ZN(n2472) );
  OAI211_X1 U3705 ( .C1(n5654), .C2(n1334), .A(n6081), .B(n6082), .ZN(n2471)
         );
  OAI222_X1 U3707 ( .A1(n5652), .A2(n1306), .B1(n7519), .B2(n1162), .C1(n7484), 
        .C2(n1190), .ZN(n2470) );
  OAI221_X1 U3711 ( .B1(n5646), .B2(n1362), .C1(n5647), .C2(n1218), .A(n2473), 
        .ZN(n2469) );
  AOI22_X1 U3712 ( .A1(\regfile/reg_out[2][1] ), .A2(n7642), .B1(
        \regfile/reg_out[3][1] ), .B2(n2323), .ZN(n2473) );
  AOI211_X1 U3715 ( .C1(\regfile/reg_out[16][1] ), .C2(n2324), .A(n2474), .B(
        n2475), .ZN(n2467) );
  OAI22_X1 U3716 ( .A1(n5624), .A2(n1292), .B1(n1348), .B2(n2327), .ZN(n2475)
         );
  OAI221_X1 U3719 ( .B1(n1405), .B2(n2328), .C1(n1204), .C2(n2329), .A(n2476), 
        .ZN(n2474) );
  AOI22_X1 U3720 ( .A1(n2331), .A2(\regfile/reg_out[12][1] ), .B1(n2332), .B2(
        \regfile/reg_out[13][1] ), .ZN(n2476) );
  AOI222_X1 U3723 ( .A1(\regfile/reg_out[27][1] ), .A2(n2333), .B1(
        \regfile/reg_out[23][1] ), .B2(n2334), .C1(\regfile/reg_out[22][1] ), 
        .C2(n2335), .ZN(n2466) );
  AOI222_X1 U3724 ( .A1(\regfile/reg_out[30][1] ), .A2(n2336), .B1(
        \regfile/reg_out[26][1] ), .B2(n2337), .C1(\regfile/reg_out[31][1] ), 
        .C2(n2338), .ZN(n2465) );
  NAND2_X1 U3725 ( .A1(n6478), .A2(n2477), .ZN(\Scc_coproc/x_exc_word[5] ) );
  NAND2_X1 U3726 ( .A1(n1054), .A2(n6479), .ZN(\Scc_coproc/x_exc_word[4] ) );
  OAI21_X1 U3728 ( .B1(\Scc_coproc/N575 ), .B2(n1057), .A(n2477), .ZN(
        \Scc_coproc/x_exc_word[3] ) );
  OAI21_X1 U3730 ( .B1(\Scc_coproc/N575 ), .B2(n1058), .A(n2478), .ZN(
        \Scc_coproc/x_exc_word[2] ) );
  OAI21_X1 U3731 ( .B1(\exc[DMEM_MISALIGN] ), .B2(n2479), .A(\Scc_coproc/N575 ), .ZN(n2478) );
  OAI211_X1 U3733 ( .C1(\Scc_coproc/N575 ), .C2(n1052), .A(n2480), .B(n2477), 
        .ZN(\Scc_coproc/x_exc_word[1] ) );
  OR3_X1 U3734 ( .A1(n6479), .A2(\exc[DMEM_MISALIGN] ), .A3(n2479), .ZN(n2480)
         );
  INV_X1 U3735 ( .A(\exc[ALU_OFLOW1] ), .ZN(n2479) );
  OAI221_X1 U3737 ( .B1(n6479), .B2(n1684), .C1(\Scc_coproc/N575 ), .C2(n1551), 
        .A(n2477), .ZN(\Scc_coproc/x_exc_word[0] ) );
  INV_X1 U3741 ( .A(\Scc_coproc/N575 ), .ZN(n6479) );
  INV_X1 U3742 ( .A(n1590), .ZN(\Scc_coproc/interrupt[9] ) );
  NAND2_X1 U3743 ( .A1(INTERRUPT_VECTOR[7]), .A2(n2481), .ZN(n1590) );
  INV_X1 U3744 ( .A(n5721), .ZN(n2481) );
  INV_X1 U3745 ( .A(n1591), .ZN(\Scc_coproc/interrupt[8] ) );
  NAND2_X1 U3746 ( .A1(INTERRUPT_VECTOR[6]), .A2(n2482), .ZN(n1591) );
  INV_X1 U3747 ( .A(n5723), .ZN(n2482) );
  NOR2_X1 U3748 ( .A1(n2483), .A2(n5725), .ZN(\Scc_coproc/interrupt[7] ) );
  INV_X1 U3749 ( .A(INTERRUPT_VECTOR[5]), .ZN(n2483) );
  NOR2_X1 U3750 ( .A1(n2484), .A2(n5727), .ZN(\Scc_coproc/interrupt[6] ) );
  INV_X1 U3751 ( .A(INTERRUPT_VECTOR[4]), .ZN(n2484) );
  NOR2_X1 U3752 ( .A1(n2485), .A2(n5729), .ZN(\Scc_coproc/interrupt[5] ) );
  INV_X1 U3753 ( .A(INTERRUPT_VECTOR[3]), .ZN(n2485) );
  INV_X1 U3754 ( .A(n5742), .ZN(\Scc_coproc/interrupt[4] ) );
  NAND2_X1 U3755 ( .A1(INTERRUPT_VECTOR[2]), .A2(n2486), .ZN(n5742) );
  INV_X1 U3756 ( .A(n5731), .ZN(n2486) );
  NOR2_X1 U3757 ( .A1(n2487), .A2(n5733), .ZN(\Scc_coproc/interrupt[3] ) );
  INV_X1 U3758 ( .A(INTERRUPT_VECTOR[1]), .ZN(n2487) );
  NOR2_X1 U3760 ( .A1(\Scc_coproc/N587 ), .A2(n1580), .ZN(
        \Scc_coproc/interrupt_active ) );
  INV_X1 U3761 ( .A(n6492), .ZN(n1580) );
  INV_X1 U3762 ( .A(\Mpath/the_alu/N491 ), .ZN(\Mpath/the_alu/N492 ) );
  INV_X1 U3764 ( .A(\Mcontrol/bp_logicA/exec_main ), .ZN(n2488) );
  NAND2_X1 U3765 ( .A1(\Mcontrol/bp_logicB/memory_main ), .A2(n2489), .ZN(
        \Mcontrol/st_logic/N42 ) );
  INV_X1 U3766 ( .A(\Mcontrol/bp_logicB/exec_main ), .ZN(n2489) );
  INV_X1 U3769 ( .A(n6044), .ZN(n6041) );
  NAND2_X1 U3770 ( .A1(\Mcontrol/d_sampled_finstr [20]), .A2(n7207), .ZN(n6044) );
  OAI21_X1 U3771 ( .B1(n7534), .B2(n7571), .A(n6971), .ZN(n2490) );
  NAND2_X1 U3776 ( .A1(\Mcontrol/d_sampled_finstr [19]), .A2(n7207), .ZN(n6046) );
  AOI21_X1 U3778 ( .B1(n7451), .B2(n1423), .A(n2495), .ZN(n2493) );
  AOI21_X1 U3779 ( .B1(n6060), .B2(n2496), .A(n2497), .ZN(n2495) );
  INV_X1 U3780 ( .A(n6069), .ZN(n2496) );
  INV_X1 U3781 ( .A(n7547), .ZN(n6060) );
  INV_X1 U3782 ( .A(n6039), .ZN(n1423) );
  NAND2_X1 U3783 ( .A1(\Mcontrol/d_sampled_finstr [18]), .A2(n7207), .ZN(n6039) );
  OAI21_X1 U3784 ( .B1(n5743), .B2(n2498), .A(n1673), .ZN(
        \Mcontrol/d_jump_type[1] ) );
  AOI21_X1 U3785 ( .B1(n2492), .B2(n6038), .A(net56977), .ZN(n2498) );
  INV_X1 U3788 ( .A(n6049), .ZN(n6038) );
  NAND2_X1 U3789 ( .A1(\Mcontrol/d_sampled_finstr [17]), .A2(n7207), .ZN(n6049) );
  NAND2_X1 U3790 ( .A1(n7571), .A2(n7576), .ZN(n2492) );
  OAI21_X1 U3798 ( .B1(n6042), .B2(n7534), .A(n2502), .ZN(n2501) );
  INV_X1 U3802 ( .A(\Mcontrol/Operation_decoding32/N1928 ), .ZN(n1846) );
  INV_X1 U3804 ( .A(n6042), .ZN(n1417) );
  NAND2_X1 U3805 ( .A1(\Mcontrol/d_sampled_finstr [16]), .A2(n7207), .ZN(n6042) );
  INV_X1 U3812 ( .A(\Mcontrol/Operation_decoding32/N1975 ), .ZN(
        \Mcontrol/Operation_decoding32/N1976 ) );
  INV_X1 U3813 ( .A(\Mcontrol/Operation_decoding32/N1969 ), .ZN(
        \Mcontrol/Operation_decoding32/N1970 ) );
  INV_X1 U3814 ( .A(n7391), .ZN(\Mcontrol/Operation_decoding32/N1964 ) );
  INV_X1 U3815 ( .A(n7218), .ZN(\Mcontrol/Operation_decoding32/N1958 ) );
  INV_X1 U3816 ( .A(n7064), .ZN(\Mcontrol/Operation_decoding32/N1952 ) );
  OAI211_X1 U3818 ( .C1(n2504), .C2(n1557), .A(n2505), .B(n2506), .ZN(n7882)
         );
  AOI22_X1 U3820 ( .A1(epc[9]), .A2(n1562), .B1(n1563), .B2(break_code[9]), 
        .ZN(n2505) );
  OAI22_X1 U3821 ( .A1(n2507), .A2(n2508), .B1(n5904), .B2(n2509), .ZN(
        break_code[9]) );
  NAND2_X1 U3822 ( .A1(\Mcontrol/d_sampled_finstr [9]), .A2(n7207), .ZN(n5904)
         );
  INV_X1 U3823 ( .A(n6104), .ZN(n2508) );
  INV_X1 U3824 ( .A(branch_rega[9]), .ZN(n2504) );
  INV_X1 U3826 ( .A(n1011), .ZN(n2510) );
  NAND4_X1 U3827 ( .A1(n2511), .A2(n2512), .A3(n2513), .A4(n2514), .ZN(n1011)
         );
  NAND3_X1 U3829 ( .A1(n6111), .A2(n6110), .A3(n6112), .ZN(n2518) );
  OAI211_X1 U3830 ( .C1(n5654), .C2(n1013), .A(n6108), .B(n6109), .ZN(n2517)
         );
  OAI222_X1 U3832 ( .A1(n5652), .A2(n1017), .B1(n7518), .B2(n1016), .C1(n7484), 
        .C2(n1012), .ZN(n2516) );
  OAI221_X1 U3836 ( .B1(n5646), .B2(n1030), .C1(n5647), .C2(n1029), .A(n2519), 
        .ZN(n2515) );
  AOI22_X1 U3837 ( .A1(\regfile/reg_out[2][9] ), .A2(n7641), .B1(
        \regfile/reg_out[3][9] ), .B2(n2323), .ZN(n2519) );
  AOI211_X1 U3840 ( .C1(\regfile/reg_out[16][9] ), .C2(n2324), .A(n2520), .B(
        n2521), .ZN(n2513) );
  OAI22_X1 U3841 ( .A1(n5624), .A2(n1019), .B1(n1032), .B2(n2327), .ZN(n2521)
         );
  OAI221_X1 U3844 ( .B1(n1020), .B2(n2328), .C1(n1031), .C2(n2329), .A(n2522), 
        .ZN(n2520) );
  AOI22_X1 U3845 ( .A1(n2331), .A2(\regfile/reg_out[12][9] ), .B1(n2332), .B2(
        \regfile/reg_out[13][9] ), .ZN(n2522) );
  AOI222_X1 U3848 ( .A1(\regfile/reg_out[27][9] ), .A2(n2333), .B1(
        \regfile/reg_out[23][9] ), .B2(n2334), .C1(\regfile/reg_out[22][9] ), 
        .C2(n2335), .ZN(n2512) );
  AOI222_X1 U3849 ( .A1(\regfile/reg_out[30][9] ), .A2(n2336), .B1(
        \regfile/reg_out[26][9] ), .B2(n2337), .C1(\regfile/reg_out[31][9] ), 
        .C2(n2338), .ZN(n2511) );
  AOI22_X1 U3852 ( .A1(epc[8]), .A2(n1562), .B1(n1563), .B2(break_code[8]), 
        .ZN(n2524) );
  NAND2_X1 U3854 ( .A1(\Mcontrol/d_sampled_finstr [8]), .A2(n7207), .ZN(n5914)
         );
  INV_X1 U3855 ( .A(n6119), .ZN(n2526) );
  INV_X1 U3856 ( .A(branch_rega[8]), .ZN(n2523) );
  INV_X1 U3858 ( .A(n1092), .ZN(n2527) );
  NAND4_X1 U3859 ( .A1(n2528), .A2(n2529), .A3(n2530), .A4(n2531), .ZN(n1092)
         );
  NAND3_X1 U3861 ( .A1(n6124), .A2(n6123), .A3(n6125), .ZN(n2535) );
  OAI211_X1 U3862 ( .C1(n5654), .C2(n1323), .A(n6121), .B(n6122), .ZN(n2534)
         );
  OAI222_X1 U3864 ( .A1(n5652), .A2(n1295), .B1(n7518), .B2(n1151), .C1(n7484), 
        .C2(n1179), .ZN(n2533) );
  OAI221_X1 U3868 ( .B1(n5646), .B2(n1351), .C1(n5647), .C2(n1207), .A(n2536), 
        .ZN(n2532) );
  AOI22_X1 U3869 ( .A1(\regfile/reg_out[2][8] ), .A2(n7642), .B1(
        \regfile/reg_out[3][8] ), .B2(n2323), .ZN(n2536) );
  AOI211_X1 U3872 ( .C1(\regfile/reg_out[16][8] ), .C2(n2324), .A(n2537), .B(
        n2538), .ZN(n2530) );
  OAI22_X1 U3873 ( .A1(n5624), .A2(n1281), .B1(n1337), .B2(n2327), .ZN(n2538)
         );
  OAI221_X1 U3876 ( .B1(n1380), .B2(n2328), .C1(n1193), .C2(n2329), .A(n2539), 
        .ZN(n2537) );
  AOI22_X1 U3877 ( .A1(n2331), .A2(\regfile/reg_out[12][8] ), .B1(n2332), .B2(
        \regfile/reg_out[13][8] ), .ZN(n2539) );
  AOI222_X1 U3880 ( .A1(\regfile/reg_out[27][8] ), .A2(n2333), .B1(
        \regfile/reg_out[23][8] ), .B2(n2334), .C1(\regfile/reg_out[22][8] ), 
        .C2(n2335), .ZN(n2529) );
  AOI222_X1 U3881 ( .A1(\regfile/reg_out[30][8] ), .A2(n2336), .B1(
        \regfile/reg_out[26][8] ), .B2(n2337), .C1(\regfile/reg_out[31][8] ), 
        .C2(n2338), .ZN(n2528) );
  OAI211_X1 U3882 ( .C1(n2540), .C2(n1557), .A(n2541), .B(n2542), .ZN(n7883)
         );
  AOI222_X1 U3883 ( .A1(n6102), .A2(n6540), .B1(
        \Mcontrol/Nextpc_decoding/Bta [7]), .B2(n1560), .C1(jar_in[7]), .C2(
        net57184), .ZN(n2542) );
  AOI22_X1 U3884 ( .A1(epc[7]), .A2(n1562), .B1(n1563), .B2(break_code[7]), 
        .ZN(n2541) );
  OAI22_X1 U3885 ( .A1(n2507), .A2(n2543), .B1(n6106), .B2(n2509), .ZN(
        break_code[7]) );
  NAND2_X1 U3886 ( .A1(\Mcontrol/d_sampled_finstr [7]), .A2(n7207), .ZN(n6106)
         );
  INV_X1 U3887 ( .A(n6132), .ZN(n2543) );
  INV_X1 U3888 ( .A(branch_rega[7]), .ZN(n2540) );
  OAI222_X1 U3889 ( .A1(n5623), .A2(n5533), .B1(n7486), .B2(n2544), .C1(n5621), 
        .C2(n5531), .ZN(branch_rega[7]) );
  INV_X1 U3890 ( .A(n972), .ZN(n2544) );
  NAND4_X1 U3891 ( .A1(n2545), .A2(n2546), .A3(n2547), .A4(n2548), .ZN(n972)
         );
  NOR4_X1 U3892 ( .A1(n2549), .A2(n2550), .A3(n2551), .A4(n2552), .ZN(n2548)
         );
  NAND3_X1 U3893 ( .A1(n6136), .A2(n6135), .A3(n6137), .ZN(n2552) );
  OAI211_X1 U3894 ( .C1(n5654), .C2(n974), .A(n6133), .B(n6134), .ZN(n2551) );
  OAI222_X1 U3896 ( .A1(n5652), .A2(n978), .B1(n7519), .B2(n977), .C1(n7484), 
        .C2(n973), .ZN(n2550) );
  OAI221_X1 U3900 ( .B1(n5646), .B2(n991), .C1(n5647), .C2(n990), .A(n2553), 
        .ZN(n2549) );
  AOI22_X1 U3901 ( .A1(\regfile/reg_out[2][7] ), .A2(n7642), .B1(
        \regfile/reg_out[3][7] ), .B2(n2323), .ZN(n2553) );
  AOI211_X1 U3904 ( .C1(\regfile/reg_out[16][7] ), .C2(n2324), .A(n2554), .B(
        n2555), .ZN(n2547) );
  OAI22_X1 U3905 ( .A1(n5624), .A2(n980), .B1(n993), .B2(n2327), .ZN(n2555) );
  OAI221_X1 U3908 ( .B1(n981), .B2(n2328), .C1(n992), .C2(n2329), .A(n2556), 
        .ZN(n2554) );
  AOI22_X1 U3909 ( .A1(n2331), .A2(\regfile/reg_out[12][7] ), .B1(n2332), .B2(
        \regfile/reg_out[13][7] ), .ZN(n2556) );
  AOI222_X1 U3912 ( .A1(\regfile/reg_out[27][7] ), .A2(n2333), .B1(
        \regfile/reg_out[23][7] ), .B2(n2334), .C1(\regfile/reg_out[22][7] ), 
        .C2(n2335), .ZN(n2546) );
  AOI222_X1 U3913 ( .A1(\regfile/reg_out[30][7] ), .A2(n2336), .B1(
        \regfile/reg_out[26][7] ), .B2(n2337), .C1(\regfile/reg_out[31][7] ), 
        .C2(n2338), .ZN(n2545) );
  OAI211_X1 U3914 ( .C1(n2557), .C2(n1557), .A(n2558), .B(n2559), .ZN(n7884)
         );
  AOI222_X1 U3915 ( .A1(n6102), .A2(n6514), .B1(
        \Mcontrol/Nextpc_decoding/Bta [6]), .B2(n1560), .C1(jar_in[6]), .C2(
        net57184), .ZN(n2559) );
  AOI22_X1 U3916 ( .A1(epc[6]), .A2(n1562), .B1(n1563), .B2(break_code[6]), 
        .ZN(n2558) );
  OAI22_X1 U3917 ( .A1(n2507), .A2(n2560), .B1(n6120), .B2(n2509), .ZN(
        break_code[6]) );
  NAND2_X1 U3918 ( .A1(\Mcontrol/d_sampled_finstr [6]), .A2(n7207), .ZN(n6120)
         );
  INV_X1 U3919 ( .A(n6144), .ZN(n2560) );
  INV_X1 U3920 ( .A(branch_rega[6]), .ZN(n2557) );
  INV_X1 U3922 ( .A(n933), .ZN(n2561) );
  NAND4_X1 U3923 ( .A1(n2562), .A2(n2563), .A3(n2564), .A4(n2565), .ZN(n933)
         );
  NOR4_X1 U3924 ( .A1(n2566), .A2(n2567), .A3(n2568), .A4(n2569), .ZN(n2565)
         );
  NAND3_X1 U3925 ( .A1(n6148), .A2(n6147), .A3(n6149), .ZN(n2569) );
  OAI211_X1 U3926 ( .C1(n5654), .C2(n935), .A(n6145), .B(n6146), .ZN(n2568) );
  OAI222_X1 U3928 ( .A1(n5652), .A2(n939), .B1(n7519), .B2(n938), .C1(n7482), 
        .C2(n934), .ZN(n2567) );
  OAI221_X1 U3932 ( .B1(n5646), .B2(n952), .C1(n5647), .C2(n951), .A(n2570), 
        .ZN(n2566) );
  AOI22_X1 U3933 ( .A1(\regfile/reg_out[2][6] ), .A2(n7641), .B1(
        \regfile/reg_out[3][6] ), .B2(n2323), .ZN(n2570) );
  AOI211_X1 U3936 ( .C1(\regfile/reg_out[16][6] ), .C2(n2324), .A(n2571), .B(
        n2572), .ZN(n2564) );
  OAI22_X1 U3937 ( .A1(n5624), .A2(n941), .B1(n954), .B2(n2327), .ZN(n2572) );
  OAI221_X1 U3940 ( .B1(n942), .B2(n2328), .C1(n953), .C2(n2329), .A(n2573), 
        .ZN(n2571) );
  AOI22_X1 U3941 ( .A1(n2331), .A2(\regfile/reg_out[12][6] ), .B1(n2332), .B2(
        \regfile/reg_out[13][6] ), .ZN(n2573) );
  AOI222_X1 U3944 ( .A1(\regfile/reg_out[27][6] ), .A2(n2333), .B1(
        \regfile/reg_out[23][6] ), .B2(n2334), .C1(\regfile/reg_out[22][6] ), 
        .C2(n2335), .ZN(n2563) );
  AOI222_X1 U3945 ( .A1(\regfile/reg_out[30][6] ), .A2(n2336), .B1(
        \regfile/reg_out[26][6] ), .B2(n2337), .C1(\regfile/reg_out[31][6] ), 
        .C2(n2338), .ZN(n2562) );
  AOI22_X1 U3948 ( .A1(epc[5]), .A2(n1562), .B1(n1563), .B2(break_code[5]), 
        .ZN(n2575) );
  INV_X1 U3951 ( .A(n6156), .ZN(n2577) );
  INV_X1 U3952 ( .A(branch_rega[5]), .ZN(n2574) );
  INV_X1 U3954 ( .A(n889), .ZN(n2578) );
  NAND4_X1 U3955 ( .A1(n2579), .A2(n2580), .A3(n2581), .A4(n2582), .ZN(n889)
         );
  NOR4_X1 U3956 ( .A1(n2583), .A2(n2584), .A3(n2585), .A4(n2586), .ZN(n2582)
         );
  NAND3_X1 U3957 ( .A1(n6160), .A2(n6159), .A3(n6161), .ZN(n2586) );
  OAI211_X1 U3958 ( .C1(n5654), .C2(n891), .A(n6157), .B(n6158), .ZN(n2585) );
  OAI222_X1 U3960 ( .A1(n5652), .A2(n895), .B1(n7519), .B2(n894), .C1(n7484), 
        .C2(n890), .ZN(n2584) );
  OAI221_X1 U3964 ( .B1(n5646), .B2(n908), .C1(n5647), .C2(n907), .A(n2587), 
        .ZN(n2583) );
  AOI22_X1 U3965 ( .A1(\regfile/reg_out[2][5] ), .A2(n7641), .B1(
        \regfile/reg_out[3][5] ), .B2(n2323), .ZN(n2587) );
  AOI211_X1 U3968 ( .C1(\regfile/reg_out[16][5] ), .C2(n2324), .A(n2588), .B(
        n2589), .ZN(n2581) );
  OAI22_X1 U3969 ( .A1(n5624), .A2(n897), .B1(n910), .B2(n2327), .ZN(n2589) );
  OAI221_X1 U3972 ( .B1(n898), .B2(n2328), .C1(n909), .C2(n2329), .A(n2590), 
        .ZN(n2588) );
  AOI22_X1 U3973 ( .A1(n2331), .A2(\regfile/reg_out[12][5] ), .B1(n2332), .B2(
        \regfile/reg_out[13][5] ), .ZN(n2590) );
  AOI222_X1 U3976 ( .A1(\regfile/reg_out[27][5] ), .A2(n2333), .B1(
        \regfile/reg_out[23][5] ), .B2(n2334), .C1(\regfile/reg_out[22][5] ), 
        .C2(n2335), .ZN(n2580) );
  AOI222_X1 U3977 ( .A1(\regfile/reg_out[30][5] ), .A2(n2336), .B1(
        \regfile/reg_out[26][5] ), .B2(n2337), .C1(\regfile/reg_out[31][5] ), 
        .C2(n2338), .ZN(n2579) );
  OAI211_X1 U3978 ( .C1(n2591), .C2(n1557), .A(n2592), .B(n2593), .ZN(
        I_ADDR_OUTBUS[4]) );
  AOI222_X1 U3979 ( .A1(n6102), .A2(n6518), .B1(
        \Mcontrol/Nextpc_decoding/Bta [4]), .B2(n7356), .C1(net57184), .C2(
        jar_in[4]), .ZN(n2593) );
  AOI22_X1 U3980 ( .A1(epc[4]), .A2(n1562), .B1(n1563), .B2(break_code[4]), 
        .ZN(n2592) );
  OAI22_X1 U3981 ( .A1(n5516), .A2(n2594), .B1(n2595), .B2(n2596), .ZN(
        break_code[4]) );
  INV_X1 U3982 ( .A(n6169), .ZN(n2596) );
  INV_X1 U3984 ( .A(branch_rega[4]), .ZN(n2591) );
  OAI222_X1 U3985 ( .A1(n5623), .A2(n5542), .B1(n7486), .B2(n2597), .C1(n5621), 
        .C2(n5540), .ZN(branch_rega[4]) );
  INV_X1 U3986 ( .A(n1090), .ZN(n2597) );
  NAND4_X1 U3987 ( .A1(n2598), .A2(n2599), .A3(n2600), .A4(n2601), .ZN(n1090)
         );
  NOR4_X1 U3988 ( .A1(n2602), .A2(n2603), .A3(n2604), .A4(n2605), .ZN(n2601)
         );
  NAND3_X1 U3989 ( .A1(n6177), .A2(n6176), .A3(n6178), .ZN(n2605) );
  OAI211_X1 U3990 ( .C1(n5654), .C2(n1324), .A(n6174), .B(n6175), .ZN(n2604)
         );
  OAI222_X1 U3992 ( .A1(n5652), .A2(n1296), .B1(n7519), .B2(n1152), .C1(n7482), 
        .C2(n1180), .ZN(n2603) );
  OAI221_X1 U3996 ( .B1(n5646), .B2(n1352), .C1(n5647), .C2(n1208), .A(n2606), 
        .ZN(n2602) );
  AOI22_X1 U3997 ( .A1(\regfile/reg_out[2][4] ), .A2(n7641), .B1(
        \regfile/reg_out[3][4] ), .B2(n2323), .ZN(n2606) );
  AOI211_X1 U4000 ( .C1(\regfile/reg_out[16][4] ), .C2(n2324), .A(n2607), .B(
        n2608), .ZN(n2600) );
  OAI22_X1 U4001 ( .A1(n5624), .A2(n1282), .B1(n1338), .B2(n2327), .ZN(n2608)
         );
  OAI221_X1 U4004 ( .B1(n1383), .B2(n2328), .C1(n1194), .C2(n2329), .A(n2609), 
        .ZN(n2607) );
  AOI22_X1 U4005 ( .A1(n2331), .A2(\regfile/reg_out[12][4] ), .B1(n2332), .B2(
        \regfile/reg_out[13][4] ), .ZN(n2609) );
  AOI222_X1 U4008 ( .A1(\regfile/reg_out[27][4] ), .A2(n2333), .B1(
        \regfile/reg_out[23][4] ), .B2(n2334), .C1(\regfile/reg_out[22][4] ), 
        .C2(n2335), .ZN(n2599) );
  AOI222_X1 U4009 ( .A1(\regfile/reg_out[30][4] ), .A2(n2336), .B1(
        \regfile/reg_out[26][4] ), .B2(n2337), .C1(\regfile/reg_out[31][4] ), 
        .C2(n2338), .ZN(n2598) );
  OAI211_X1 U4010 ( .C1(n2610), .C2(n1557), .A(n2611), .B(n2612), .ZN(n7885)
         );
  AOI222_X1 U4011 ( .A1(n6102), .A2(n6520), .B1(
        \Mcontrol/Nextpc_decoding/Bta [3]), .B2(n7356), .C1(jar_in[3]), .C2(
        net57184), .ZN(n2612) );
  AOI22_X1 U4012 ( .A1(epc[3]), .A2(n1562), .B1(n1563), .B2(n7311), .ZN(n2611)
         );
  INV_X1 U4014 ( .A(n6185), .ZN(n2613) );
  INV_X1 U4015 ( .A(branch_rega[3]), .ZN(n2610) );
  INV_X1 U4017 ( .A(n1088), .ZN(n2614) );
  NAND4_X1 U4018 ( .A1(n2615), .A2(n2616), .A3(n2617), .A4(n2618), .ZN(n1088)
         );
  NAND3_X1 U4020 ( .A1(n6191), .A2(n6190), .A3(n6192), .ZN(n2622) );
  OAI211_X1 U4021 ( .C1(n5654), .C2(n1325), .A(n6188), .B(n6189), .ZN(n2621)
         );
  OAI222_X1 U4023 ( .A1(n5652), .A2(n1297), .B1(n7518), .B2(n1153), .C1(n7482), 
        .C2(n1181), .ZN(n2620) );
  OAI221_X1 U4027 ( .B1(n5646), .B2(n1353), .C1(n5647), .C2(n1209), .A(n2623), 
        .ZN(n2619) );
  AOI22_X1 U4028 ( .A1(\regfile/reg_out[2][3] ), .A2(n7641), .B1(
        \regfile/reg_out[3][3] ), .B2(n2323), .ZN(n2623) );
  AOI211_X1 U4031 ( .C1(\regfile/reg_out[16][3] ), .C2(n2324), .A(n2624), .B(
        n2625), .ZN(n2617) );
  OAI22_X1 U4032 ( .A1(n5624), .A2(n1283), .B1(n1339), .B2(n2327), .ZN(n2625)
         );
  OAI221_X1 U4035 ( .B1(n1386), .B2(n2328), .C1(n1195), .C2(n2329), .A(n2626), 
        .ZN(n2624) );
  AOI22_X1 U4036 ( .A1(n2331), .A2(\regfile/reg_out[12][3] ), .B1(n2332), .B2(
        \regfile/reg_out[13][3] ), .ZN(n2626) );
  AOI222_X1 U4039 ( .A1(\regfile/reg_out[27][3] ), .A2(n2333), .B1(
        \regfile/reg_out[23][3] ), .B2(n2334), .C1(\regfile/reg_out[22][3] ), 
        .C2(n2335), .ZN(n2616) );
  AOI222_X1 U4040 ( .A1(\regfile/reg_out[30][3] ), .A2(n2336), .B1(
        \regfile/reg_out[26][3] ), .B2(n2337), .C1(\regfile/reg_out[31][3] ), 
        .C2(n2338), .ZN(n2615) );
  AOI222_X1 U4042 ( .A1(n6102), .A2(n6522), .B1(
        \Mcontrol/Nextpc_decoding/Bta [2]), .B2(n7356), .C1(jar_in[2]), .C2(
        net57184), .ZN(n2629) );
  AOI22_X1 U4043 ( .A1(epc[2]), .A2(n1562), .B1(n1563), .B2(n7353), .ZN(n2628)
         );
  INV_X1 U4045 ( .A(n6199), .ZN(n2630) );
  NAND3_X1 U4046 ( .A1(n5521), .A2(net57954), .A3(n6168), .ZN(n2595) );
  INV_X1 U4050 ( .A(branch_rega[2]), .ZN(n2627) );
  INV_X1 U4052 ( .A(n1083), .ZN(n2632) );
  NAND4_X1 U4053 ( .A1(n2633), .A2(n2634), .A3(n2635), .A4(n2636), .ZN(n1083)
         );
  NOR4_X1 U4054 ( .A1(n2637), .A2(n2638), .A3(n2639), .A4(n2640), .ZN(n2636)
         );
  NAND3_X1 U4055 ( .A1(n6206), .A2(n6205), .A3(n6207), .ZN(n2640) );
  OAI211_X1 U4056 ( .C1(n5654), .C2(n1328), .A(n6203), .B(n6204), .ZN(n2639)
         );
  OAI222_X1 U4058 ( .A1(n5652), .A2(n1300), .B1(n7518), .B2(n1156), .C1(n7484), 
        .C2(n1184), .ZN(n2638) );
  OAI221_X1 U4062 ( .B1(n5646), .B2(n1356), .C1(n5647), .C2(n1212), .A(n2641), 
        .ZN(n2637) );
  AOI22_X1 U4063 ( .A1(\regfile/reg_out[2][2] ), .A2(n7642), .B1(
        \regfile/reg_out[3][2] ), .B2(n2323), .ZN(n2641) );
  AOI211_X1 U4066 ( .C1(\regfile/reg_out[16][2] ), .C2(n2324), .A(n2642), .B(
        n2643), .ZN(n2635) );
  OAI22_X1 U4067 ( .A1(n5624), .A2(n1286), .B1(n1342), .B2(n2327), .ZN(n2643)
         );
  OAI221_X1 U4070 ( .B1(n1392), .B2(n2328), .C1(n1198), .C2(n2329), .A(n2644), 
        .ZN(n2642) );
  AOI22_X1 U4071 ( .A1(n2331), .A2(\regfile/reg_out[12][2] ), .B1(n2332), .B2(
        \regfile/reg_out[13][2] ), .ZN(n2644) );
  AOI222_X1 U4074 ( .A1(\regfile/reg_out[27][2] ), .A2(n2333), .B1(
        \regfile/reg_out[23][2] ), .B2(n2334), .C1(\regfile/reg_out[22][2] ), 
        .C2(n2335), .ZN(n2634) );
  AOI222_X1 U4075 ( .A1(\regfile/reg_out[30][2] ), .A2(n2336), .B1(
        \regfile/reg_out[26][2] ), .B2(n2337), .C1(\regfile/reg_out[31][2] ), 
        .C2(n2338), .ZN(n2633) );
  AOI221_X1 U4080 ( .B1(\Mcontrol/d_instr [7]), .B2(n333), .C1(n6214), .C2(
        n331), .A(n330), .ZN(n1623) );
  OAI222_X1 U4083 ( .A1(n5623), .A2(n5575), .B1(n7487), .B2(n2649), .C1(n5621), 
        .C2(n5573), .ZN(branch_rega[23]) );
  INV_X1 U4084 ( .A(n1081), .ZN(n2649) );
  NAND4_X1 U4085 ( .A1(n2650), .A2(n2651), .A3(n2652), .A4(n2653), .ZN(n1081)
         );
  NAND3_X1 U4087 ( .A1(n6218), .A2(n6217), .A3(n6219), .ZN(n2657) );
  OAI211_X1 U4088 ( .C1(n5654), .C2(n1333), .A(n6215), .B(n6216), .ZN(n2656)
         );
  OAI222_X1 U4090 ( .A1(n5652), .A2(n1305), .B1(n7519), .B2(n1161), .C1(n7482), 
        .C2(n1189), .ZN(n2655) );
  OAI221_X1 U4094 ( .B1(n5646), .B2(n1361), .C1(n5647), .C2(n1217), .A(n2658), 
        .ZN(n2654) );
  AOI22_X1 U4095 ( .A1(\regfile/reg_out[2][23] ), .A2(n7641), .B1(
        \regfile/reg_out[3][23] ), .B2(n2323), .ZN(n2658) );
  AOI211_X1 U4098 ( .C1(\regfile/reg_out[16][23] ), .C2(n2324), .A(n2659), .B(
        n2660), .ZN(n2652) );
  OAI22_X1 U4099 ( .A1(n5624), .A2(n1291), .B1(n1347), .B2(n2327), .ZN(n2660)
         );
  OAI221_X1 U4102 ( .B1(n1403), .B2(n2328), .C1(n1203), .C2(n2329), .A(n2661), 
        .ZN(n2659) );
  AOI22_X1 U4103 ( .A1(n2331), .A2(\regfile/reg_out[12][23] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][23] ), .ZN(n2661) );
  AOI222_X1 U4106 ( .A1(\regfile/reg_out[27][23] ), .A2(n2333), .B1(
        \regfile/reg_out[23][23] ), .B2(n2334), .C1(\regfile/reg_out[22][23] ), 
        .C2(n2335), .ZN(n2651) );
  AOI222_X1 U4107 ( .A1(\regfile/reg_out[30][23] ), .A2(n2336), .B1(
        \regfile/reg_out[26][23] ), .B2(n2337), .C1(\regfile/reg_out[31][23] ), 
        .C2(n2338), .ZN(n2650) );
  INV_X1 U4116 ( .A(n379), .ZN(n2666) );
  NAND4_X1 U4117 ( .A1(n2670), .A2(n2668), .A3(n2669), .A4(n2667), .ZN(n379)
         );
  NAND3_X1 U4119 ( .A1(n6231), .A2(n6230), .A3(n6232), .ZN(n2674) );
  OAI211_X1 U4120 ( .C1(n5654), .C2(n381), .A(n6228), .B(n6229), .ZN(n2673) );
  OAI222_X1 U4122 ( .A1(n5652), .A2(n385), .B1(n7518), .B2(n384), .C1(n7484), 
        .C2(n380), .ZN(n2672) );
  OAI221_X1 U4126 ( .B1(n5646), .B2(n398), .C1(n5647), .C2(n397), .A(n2675), 
        .ZN(n2671) );
  AOI22_X1 U4127 ( .A1(\regfile/reg_out[2][22] ), .A2(n7641), .B1(
        \regfile/reg_out[3][22] ), .B2(n2323), .ZN(n2675) );
  AOI211_X1 U4130 ( .C1(\regfile/reg_out[16][22] ), .C2(n2324), .A(n2676), .B(
        n2677), .ZN(n2669) );
  OAI22_X1 U4131 ( .A1(n5624), .A2(n387), .B1(n400), .B2(n2327), .ZN(n2677) );
  OAI221_X1 U4134 ( .B1(n388), .B2(n2328), .C1(n399), .C2(n2329), .A(n2678), 
        .ZN(n2676) );
  AOI22_X1 U4135 ( .A1(n2331), .A2(\regfile/reg_out[12][22] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][22] ), .ZN(n2678) );
  AOI222_X1 U4138 ( .A1(\regfile/reg_out[27][22] ), .A2(n2333), .B1(
        \regfile/reg_out[23][22] ), .B2(n2334), .C1(\regfile/reg_out[22][22] ), 
        .C2(n2335), .ZN(n2668) );
  AOI222_X1 U4139 ( .A1(\regfile/reg_out[30][22] ), .A2(n2336), .B1(
        \regfile/reg_out[26][22] ), .B2(n2337), .C1(\regfile/reg_out[31][22] ), 
        .C2(n2338), .ZN(n2667) );
  OAI211_X1 U4140 ( .C1(n2679), .C2(n1557), .A(n2681), .B(n2680), .ZN(n7871)
         );
  AOI22_X1 U4142 ( .A1(n1562), .A2(n2682), .B1(n1563), .B2(break_code[21]), 
        .ZN(n2680) );
  INV_X1 U4143 ( .A(n410), .ZN(break_code[21]) );
  INV_X1 U4145 ( .A(n6246), .ZN(n2682) );
  INV_X1 U4146 ( .A(branch_rega[21]), .ZN(n2679) );
  INV_X1 U4148 ( .A(n415), .ZN(n2683) );
  NAND4_X1 U4149 ( .A1(n2684), .A2(n2685), .A3(n2686), .A4(n2687), .ZN(n415)
         );
  NOR4_X1 U4150 ( .A1(n2688), .A2(n2689), .A3(n2690), .A4(n2691), .ZN(n2687)
         );
  NAND3_X1 U4151 ( .A1(n6243), .A2(n6242), .A3(n6244), .ZN(n2691) );
  OAI211_X1 U4152 ( .C1(n5654), .C2(n417), .A(n6240), .B(n6241), .ZN(n2690) );
  OAI222_X1 U4154 ( .A1(n5652), .A2(n421), .B1(n7518), .B2(n420), .C1(n7484), 
        .C2(n416), .ZN(n2689) );
  OAI221_X1 U4158 ( .B1(n5646), .B2(n434), .C1(n5647), .C2(n433), .A(n2692), 
        .ZN(n2688) );
  AOI22_X1 U4159 ( .A1(\regfile/reg_out[2][21] ), .A2(n7642), .B1(
        \regfile/reg_out[3][21] ), .B2(n2323), .ZN(n2692) );
  AOI211_X1 U4162 ( .C1(\regfile/reg_out[16][21] ), .C2(n2324), .A(n2693), .B(
        n2694), .ZN(n2686) );
  OAI22_X1 U4163 ( .A1(n5624), .A2(n423), .B1(n436), .B2(n2327), .ZN(n2694) );
  OAI221_X1 U4166 ( .B1(n424), .B2(n2328), .C1(n435), .C2(n2329), .A(n2695), 
        .ZN(n2693) );
  AOI22_X1 U4167 ( .A1(n2331), .A2(\regfile/reg_out[12][21] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][21] ), .ZN(n2695) );
  AOI222_X1 U4170 ( .A1(\regfile/reg_out[27][21] ), .A2(n2333), .B1(
        \regfile/reg_out[23][21] ), .B2(n2334), .C1(\regfile/reg_out[22][21] ), 
        .C2(n2335), .ZN(n2685) );
  AOI222_X1 U4171 ( .A1(\regfile/reg_out[30][21] ), .A2(n2336), .B1(
        \regfile/reg_out[26][21] ), .B2(n2337), .C1(\regfile/reg_out[31][21] ), 
        .C2(n2338), .ZN(n2684) );
  OAI211_X1 U4172 ( .C1(n2696), .C2(n1557), .A(n2697), .B(n2698), .ZN(n7872)
         );
  AOI22_X1 U4174 ( .A1(n1562), .A2(n2699), .B1(n1563), .B2(break_code[20]), 
        .ZN(n2697) );
  INV_X1 U4175 ( .A(n445), .ZN(break_code[20]) );
  OAI21_X1 U4177 ( .B1(n5880), .B2(n1523), .A(n213), .ZN(n330) );
  INV_X1 U4178 ( .A(n1663), .ZN(n213) );
  AND2_X1 U4179 ( .A1(n5847), .A2(n215), .ZN(n331) );
  AND2_X1 U4180 ( .A1(n7159), .A2(n215), .ZN(n333) );
  INV_X1 U4181 ( .A(n6262), .ZN(n2699) );
  INV_X1 U4182 ( .A(branch_rega[20]), .ZN(n2696) );
  INV_X1 U4184 ( .A(n450), .ZN(n2700) );
  NAND4_X1 U4185 ( .A1(n2701), .A2(n2702), .A3(n2703), .A4(n2704), .ZN(n450)
         );
  NOR4_X1 U4186 ( .A1(n2705), .A2(n2706), .A3(n2707), .A4(n2708), .ZN(n2704)
         );
  NAND3_X1 U4187 ( .A1(n6259), .A2(n6258), .A3(n6260), .ZN(n2708) );
  OAI211_X1 U4188 ( .C1(n5654), .C2(n452), .A(n6256), .B(n6257), .ZN(n2707) );
  OAI222_X1 U4190 ( .A1(n5652), .A2(n456), .B1(n7519), .B2(n455), .C1(n7484), 
        .C2(n451), .ZN(n2706) );
  OAI221_X1 U4194 ( .B1(n5646), .B2(n469), .C1(n5647), .C2(n468), .A(n2709), 
        .ZN(n2705) );
  AOI22_X1 U4195 ( .A1(\regfile/reg_out[2][20] ), .A2(n7641), .B1(
        \regfile/reg_out[3][20] ), .B2(n2323), .ZN(n2709) );
  AOI211_X1 U4198 ( .C1(\regfile/reg_out[16][20] ), .C2(n2324), .A(n2710), .B(
        n2711), .ZN(n2703) );
  OAI22_X1 U4199 ( .A1(n5624), .A2(n458), .B1(n471), .B2(n2327), .ZN(n2711) );
  OAI221_X1 U4202 ( .B1(n459), .B2(n2328), .C1(n470), .C2(n2329), .A(n2712), 
        .ZN(n2710) );
  AOI22_X1 U4203 ( .A1(n2331), .A2(\regfile/reg_out[12][20] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][20] ), .ZN(n2712) );
  AOI222_X1 U4206 ( .A1(\regfile/reg_out[27][20] ), .A2(n2333), .B1(
        \regfile/reg_out[23][20] ), .B2(n2334), .C1(\regfile/reg_out[22][20] ), 
        .C2(n2335), .ZN(n2702) );
  AOI222_X1 U4207 ( .A1(\regfile/reg_out[30][20] ), .A2(n2336), .B1(
        \regfile/reg_out[26][20] ), .B2(n2337), .C1(\regfile/reg_out[31][20] ), 
        .C2(n2338), .ZN(n2701) );
  OAI211_X1 U4208 ( .C1(n2713), .C2(n1557), .A(n2714), .B(n2715), .ZN(
        I_ADDR_OUTBUS[19]) );
  AOI22_X1 U4210 ( .A1(n1562), .A2(n2716), .B1(n1563), .B2(break_code[19]), 
        .ZN(n2714) );
  INV_X1 U4213 ( .A(n6267), .ZN(n2717) );
  INV_X1 U4214 ( .A(n6275), .ZN(n2716) );
  INV_X1 U4215 ( .A(branch_rega[19]), .ZN(n2713) );
  INV_X1 U4217 ( .A(n485), .ZN(n2720) );
  NAND4_X1 U4218 ( .A1(n2721), .A2(n2722), .A3(n2723), .A4(n2724), .ZN(n485)
         );
  NOR4_X1 U4219 ( .A1(n2725), .A2(n2726), .A3(n2727), .A4(n2728), .ZN(n2724)
         );
  NAND3_X1 U4220 ( .A1(n6272), .A2(n6271), .A3(n6273), .ZN(n2728) );
  OAI211_X1 U4221 ( .C1(n5654), .C2(n487), .A(n6269), .B(n6270), .ZN(n2727) );
  OAI222_X1 U4223 ( .A1(n5652), .A2(n491), .B1(n7519), .B2(n490), .C1(n7484), 
        .C2(n486), .ZN(n2726) );
  OAI221_X1 U4227 ( .B1(n5646), .B2(n504), .C1(n5647), .C2(n503), .A(n2729), 
        .ZN(n2725) );
  AOI22_X1 U4228 ( .A1(\regfile/reg_out[2][19] ), .A2(n7642), .B1(
        \regfile/reg_out[3][19] ), .B2(n2323), .ZN(n2729) );
  AOI211_X1 U4231 ( .C1(\regfile/reg_out[16][19] ), .C2(n2324), .A(n2730), .B(
        n2731), .ZN(n2723) );
  OAI22_X1 U4232 ( .A1(n5624), .A2(n493), .B1(n506), .B2(n2327), .ZN(n2731) );
  OAI221_X1 U4235 ( .B1(n494), .B2(n2328), .C1(n505), .C2(n2329), .A(n2732), 
        .ZN(n2730) );
  AOI22_X1 U4236 ( .A1(n2331), .A2(\regfile/reg_out[12][19] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][19] ), .ZN(n2732) );
  AOI222_X1 U4239 ( .A1(\regfile/reg_out[27][19] ), .A2(n2333), .B1(
        \regfile/reg_out[23][19] ), .B2(n2334), .C1(\regfile/reg_out[22][19] ), 
        .C2(n2335), .ZN(n2722) );
  AOI222_X1 U4240 ( .A1(\regfile/reg_out[30][19] ), .A2(n2336), .B1(
        \regfile/reg_out[26][19] ), .B2(n2337), .C1(\regfile/reg_out[31][19] ), 
        .C2(n2338), .ZN(n2721) );
  OAI211_X1 U4241 ( .C1(n2733), .C2(n1557), .A(n2734), .B(n2735), .ZN(n7873)
         );
  AOI22_X1 U4243 ( .A1(n1562), .A2(n2736), .B1(n1563), .B2(break_code[18]), 
        .ZN(n2734) );
  NAND2_X1 U4245 ( .A1(\Mcontrol/d_sampled_finstr [2]), .A2(n7278), .ZN(n5518)
         );
  INV_X1 U4246 ( .A(n6280), .ZN(n2737) );
  INV_X1 U4247 ( .A(n6290), .ZN(n2736) );
  INV_X1 U4248 ( .A(branch_rega[18]), .ZN(n2733) );
  OAI222_X1 U4249 ( .A1(n5623), .A2(n5593), .B1(n7487), .B2(n2738), .C1(n5621), 
        .C2(n5591), .ZN(branch_rega[18]) );
  INV_X1 U4250 ( .A(n520), .ZN(n2738) );
  NAND4_X1 U4251 ( .A1(n2739), .A2(n2740), .A3(n2741), .A4(n2742), .ZN(n520)
         );
  NOR4_X1 U4252 ( .A1(n2743), .A2(n2744), .A3(n2745), .A4(n2746), .ZN(n2742)
         );
  NAND3_X1 U4253 ( .A1(n6287), .A2(n6286), .A3(n6288), .ZN(n2746) );
  OAI211_X1 U4254 ( .C1(n5654), .C2(n522), .A(n6284), .B(n6285), .ZN(n2745) );
  OAI222_X1 U4256 ( .A1(n5652), .A2(n526), .B1(n7518), .B2(n525), .C1(n7482), 
        .C2(n521), .ZN(n2744) );
  OAI221_X1 U4260 ( .B1(n5646), .B2(n539), .C1(n5647), .C2(n538), .A(n2747), 
        .ZN(n2743) );
  AOI22_X1 U4261 ( .A1(\regfile/reg_out[2][18] ), .A2(n7642), .B1(
        \regfile/reg_out[3][18] ), .B2(n2323), .ZN(n2747) );
  AOI211_X1 U4264 ( .C1(\regfile/reg_out[16][18] ), .C2(n2324), .A(n2748), .B(
        n2749), .ZN(n2741) );
  OAI22_X1 U4265 ( .A1(n5624), .A2(n528), .B1(n541), .B2(n2327), .ZN(n2749) );
  OAI221_X1 U4268 ( .B1(n529), .B2(n2328), .C1(n540), .C2(n2329), .A(n2750), 
        .ZN(n2748) );
  AOI22_X1 U4269 ( .A1(n2331), .A2(\regfile/reg_out[12][18] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][18] ), .ZN(n2750) );
  AOI222_X1 U4272 ( .A1(\regfile/reg_out[27][18] ), .A2(n2333), .B1(
        \regfile/reg_out[23][18] ), .B2(n2334), .C1(\regfile/reg_out[22][18] ), 
        .C2(n2335), .ZN(n2740) );
  AOI222_X1 U4273 ( .A1(\regfile/reg_out[30][18] ), .A2(n2336), .B1(
        \regfile/reg_out[26][18] ), .B2(n2337), .C1(\regfile/reg_out[31][18] ), 
        .C2(n2338), .ZN(n2739) );
  OAI211_X1 U4274 ( .C1(n2751), .C2(n1557), .A(n2752), .B(n2753), .ZN(n7874)
         );
  AOI22_X1 U4276 ( .A1(n1562), .A2(n2754), .B1(n1563), .B2(break_code[17]), 
        .ZN(n2752) );
  OAI221_X1 U4277 ( .B1(n2500), .B2(n2755), .C1(n5519), .C2(n2718), .A(n2719), 
        .ZN(break_code[17]) );
  NAND2_X1 U4278 ( .A1(\Mcontrol/d_sampled_finstr [1]), .A2(n7278), .ZN(n5519)
         );
  INV_X1 U4279 ( .A(n6295), .ZN(n2755) );
  INV_X1 U4280 ( .A(n6304), .ZN(n2754) );
  INV_X1 U4281 ( .A(branch_rega[17]), .ZN(n2751) );
  OAI222_X1 U4282 ( .A1(n5623), .A2(n5596), .B1(n7487), .B2(n2756), .C1(n5621), 
        .C2(n5594), .ZN(branch_rega[17]) );
  INV_X1 U4283 ( .A(n555), .ZN(n2756) );
  NAND4_X1 U4284 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .ZN(n555)
         );
  NOR4_X1 U4285 ( .A1(n2761), .A2(n2762), .A3(n2763), .A4(n2764), .ZN(n2760)
         );
  NAND3_X1 U4286 ( .A1(n6301), .A2(n6300), .A3(n6302), .ZN(n2764) );
  OAI211_X1 U4287 ( .C1(n5654), .C2(n557), .A(n6298), .B(n6299), .ZN(n2763) );
  OAI222_X1 U4289 ( .A1(n5652), .A2(n561), .B1(n7519), .B2(n560), .C1(n7482), 
        .C2(n556), .ZN(n2762) );
  OAI221_X1 U4293 ( .B1(n5646), .B2(n574), .C1(n5647), .C2(n573), .A(n2765), 
        .ZN(n2761) );
  AOI22_X1 U4294 ( .A1(\regfile/reg_out[2][17] ), .A2(n7642), .B1(
        \regfile/reg_out[3][17] ), .B2(n2323), .ZN(n2765) );
  AOI211_X1 U4297 ( .C1(\regfile/reg_out[16][17] ), .C2(n2324), .A(n2766), .B(
        n2767), .ZN(n2759) );
  OAI22_X1 U4298 ( .A1(n5624), .A2(n563), .B1(n576), .B2(n2327), .ZN(n2767) );
  OAI221_X1 U4301 ( .B1(n564), .B2(n2328), .C1(n575), .C2(n2329), .A(n2768), 
        .ZN(n2766) );
  AOI22_X1 U4302 ( .A1(n2331), .A2(\regfile/reg_out[12][17] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][17] ), .ZN(n2768) );
  AOI222_X1 U4305 ( .A1(\regfile/reg_out[27][17] ), .A2(n2333), .B1(
        \regfile/reg_out[23][17] ), .B2(n2334), .C1(\regfile/reg_out[22][17] ), 
        .C2(n2335), .ZN(n2758) );
  AOI222_X1 U4306 ( .A1(\regfile/reg_out[30][17] ), .A2(n2336), .B1(
        \regfile/reg_out[26][17] ), .B2(n2337), .C1(\regfile/reg_out[31][17] ), 
        .C2(n2338), .ZN(n2757) );
  OAI211_X1 U4307 ( .C1(n2769), .C2(n1557), .A(n2770), .B(n2771), .ZN(n7875)
         );
  AOI22_X1 U4309 ( .A1(n1562), .A2(n2772), .B1(n1563), .B2(break_code[16]), 
        .ZN(n2770) );
  OAI221_X1 U4310 ( .B1(n2500), .B2(n2773), .C1(n5520), .C2(n2718), .A(n2719), 
        .ZN(break_code[16]) );
  AOI21_X1 U4311 ( .B1(n1533), .B2(n6268), .A(n1663), .ZN(n2719) );
  NOR3_X1 U4312 ( .A1(net56846), .A2(n5846), .A3(n1434), .ZN(n1663) );
  NAND2_X1 U4313 ( .A1(n215), .A2(n2774), .ZN(n2718) );
  INV_X1 U4314 ( .A(n1523), .ZN(n215) );
  NAND2_X1 U4315 ( .A1(\Mcontrol/d_sampled_finstr [0]), .A2(n7278), .ZN(n5520)
         );
  INV_X1 U4316 ( .A(n6309), .ZN(n2773) );
  INV_X1 U4320 ( .A(n6316), .ZN(n2772) );
  INV_X1 U4321 ( .A(branch_rega[16]), .ZN(n2769) );
  OAI222_X1 U4322 ( .A1(n5623), .A2(n5599), .B1(n7486), .B2(n2775), .C1(n5621), 
        .C2(n5597), .ZN(branch_rega[16]) );
  INV_X1 U4323 ( .A(n590), .ZN(n2775) );
  NAND4_X1 U4324 ( .A1(n2776), .A2(n2777), .A3(n2778), .A4(n2779), .ZN(n590)
         );
  NOR4_X1 U4325 ( .A1(n2780), .A2(n2781), .A3(n2782), .A4(n2783), .ZN(n2779)
         );
  NAND3_X1 U4326 ( .A1(n6313), .A2(n6312), .A3(n6314), .ZN(n2783) );
  OAI211_X1 U4327 ( .C1(n5654), .C2(n592), .A(n6310), .B(n6311), .ZN(n2782) );
  OAI222_X1 U4329 ( .A1(n5652), .A2(n596), .B1(n7518), .B2(n595), .C1(n7484), 
        .C2(n591), .ZN(n2781) );
  OAI221_X1 U4333 ( .B1(n5646), .B2(n609), .C1(n5647), .C2(n608), .A(n2784), 
        .ZN(n2780) );
  AOI22_X1 U4334 ( .A1(\regfile/reg_out[2][16] ), .A2(n7641), .B1(
        \regfile/reg_out[3][16] ), .B2(n2323), .ZN(n2784) );
  AOI211_X1 U4337 ( .C1(\regfile/reg_out[16][16] ), .C2(n2324), .A(n2785), .B(
        n2786), .ZN(n2778) );
  OAI22_X1 U4338 ( .A1(n5624), .A2(n598), .B1(n611), .B2(n2327), .ZN(n2786) );
  OAI221_X1 U4341 ( .B1(n599), .B2(n2328), .C1(n610), .C2(n2329), .A(n2787), 
        .ZN(n2785) );
  AOI22_X1 U4342 ( .A1(n2331), .A2(\regfile/reg_out[12][16] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][16] ), .ZN(n2787) );
  AOI222_X1 U4345 ( .A1(\regfile/reg_out[27][16] ), .A2(n2333), .B1(
        \regfile/reg_out[23][16] ), .B2(n2334), .C1(\regfile/reg_out[22][16] ), 
        .C2(n2335), .ZN(n2777) );
  AOI222_X1 U4346 ( .A1(\regfile/reg_out[30][16] ), .A2(n2336), .B1(
        \regfile/reg_out[26][16] ), .B2(n2337), .C1(\regfile/reg_out[31][16] ), 
        .C2(n2338), .ZN(n2776) );
  OAI211_X1 U4347 ( .C1(n2788), .C2(n1557), .A(n2789), .B(n2790), .ZN(n7876)
         );
  AOI222_X1 U4348 ( .A1(n6102), .A2(n6546), .B1(
        \Mcontrol/Nextpc_decoding/Bta [15]), .B2(n7356), .C1(jar_in[15]), .C2(
        net57184), .ZN(n2790) );
  AOI22_X1 U4349 ( .A1(epc[15]), .A2(n1562), .B1(n1563), .B2(break_code[15]), 
        .ZN(n2789) );
  OAI33_X1 U4350 ( .A1(n1474), .A2(n5846), .A3(net57323), .B1(n2774), .B2(
        n2791), .B3(n1523), .ZN(break_code[15]) );
  AOI21_X1 U4357 ( .B1(n6322), .B2(n7434), .A(n6268), .ZN(n2791) );
  INV_X1 U4358 ( .A(n7436), .ZN(n2774) );
  NAND2_X1 U4359 ( .A1(n7207), .A2(\Mcontrol/d_sampled_finstr [15]), .ZN(n5846) );
  INV_X1 U4361 ( .A(branch_rega[15]), .ZN(n2788) );
  INV_X1 U4363 ( .A(n631), .ZN(n2793) );
  NAND4_X1 U4364 ( .A1(n2794), .A2(n2795), .A3(n2796), .A4(n2797), .ZN(n631)
         );
  NAND3_X1 U4366 ( .A1(n6326), .A2(n6325), .A3(n6327), .ZN(n2801) );
  OAI211_X1 U4367 ( .C1(n5654), .C2(n633), .A(n6323), .B(n6324), .ZN(n2800) );
  OAI222_X1 U4369 ( .A1(n5652), .A2(n637), .B1(n7518), .B2(n636), .C1(n7482), 
        .C2(n632), .ZN(n2799) );
  OAI221_X1 U4373 ( .B1(n5646), .B2(n650), .C1(n5647), .C2(n649), .A(n2802), 
        .ZN(n2798) );
  AOI22_X1 U4374 ( .A1(\regfile/reg_out[2][15] ), .A2(n7641), .B1(
        \regfile/reg_out[3][15] ), .B2(n2323), .ZN(n2802) );
  AOI211_X1 U4377 ( .C1(\regfile/reg_out[16][15] ), .C2(n2324), .A(n2803), .B(
        n2804), .ZN(n2796) );
  OAI22_X1 U4378 ( .A1(n5624), .A2(n639), .B1(n652), .B2(n2327), .ZN(n2804) );
  OAI221_X1 U4381 ( .B1(n640), .B2(n2328), .C1(n651), .C2(n2329), .A(n2805), 
        .ZN(n2803) );
  AOI22_X1 U4382 ( .A1(n2331), .A2(\regfile/reg_out[12][15] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][15] ), .ZN(n2805) );
  AOI222_X1 U4385 ( .A1(\regfile/reg_out[27][15] ), .A2(n2333), .B1(
        \regfile/reg_out[23][15] ), .B2(n2334), .C1(\regfile/reg_out[22][15] ), 
        .C2(n2335), .ZN(n2795) );
  AOI222_X1 U4386 ( .A1(\regfile/reg_out[30][15] ), .A2(n2336), .B1(
        \regfile/reg_out[26][15] ), .B2(n2337), .C1(\regfile/reg_out[31][15] ), 
        .C2(n2338), .ZN(n2794) );
  OAI211_X1 U4387 ( .C1(n2806), .C2(n1557), .A(n2807), .B(n2808), .ZN(n7877)
         );
  AOI222_X1 U4388 ( .A1(n6102), .A2(n6523), .B1(
        \Mcontrol/Nextpc_decoding/Bta [14]), .B2(n7356), .C1(jar_in[14]), .C2(
        net57184), .ZN(n2808) );
  AOI22_X1 U4389 ( .A1(epc[14]), .A2(n1562), .B1(n1563), .B2(break_code[14]), 
        .ZN(n2807) );
  OAI22_X1 U4390 ( .A1(n2507), .A2(n2809), .B1(n6047), .B2(n2509), .ZN(
        break_code[14]) );
  NAND2_X1 U4391 ( .A1(\Mcontrol/d_sampled_finstr [14]), .A2(n7207), .ZN(n6047) );
  INV_X1 U4392 ( .A(n6334), .ZN(n2809) );
  INV_X1 U4393 ( .A(branch_rega[14]), .ZN(n2806) );
  INV_X1 U4395 ( .A(n1075), .ZN(n2810) );
  NAND4_X1 U4396 ( .A1(n2811), .A2(n2812), .A3(n2813), .A4(n2814), .ZN(n1075)
         );
  NOR4_X1 U4397 ( .A1(n2816), .A2(n2815), .A3(n2817), .A4(n2818), .ZN(n2814)
         );
  NAND3_X1 U4398 ( .A1(n6338), .A2(n6337), .A3(n6339), .ZN(n2818) );
  OAI211_X1 U4399 ( .C1(n5654), .C2(n1335), .A(n6335), .B(n6336), .ZN(n2817)
         );
  OAI222_X1 U4401 ( .A1(n5652), .A2(n1307), .B1(n7518), .B2(n1163), .C1(n7483), 
        .C2(n1191), .ZN(n2816) );
  OAI221_X1 U4405 ( .B1(n5646), .B2(n1363), .C1(n5647), .C2(n1219), .A(n2819), 
        .ZN(n2815) );
  AOI22_X1 U4406 ( .A1(\regfile/reg_out[2][14] ), .A2(n7642), .B1(
        \regfile/reg_out[3][14] ), .B2(n2323), .ZN(n2819) );
  AOI211_X1 U4409 ( .C1(\regfile/reg_out[16][14] ), .C2(n2324), .A(n2820), .B(
        n2821), .ZN(n2813) );
  OAI22_X1 U4410 ( .A1(n5624), .A2(n1293), .B1(n1349), .B2(n2327), .ZN(n2821)
         );
  OAI221_X1 U4413 ( .B1(n1407), .B2(n2328), .C1(n1205), .C2(n2329), .A(n2822), 
        .ZN(n2820) );
  AOI22_X1 U4414 ( .A1(n2331), .A2(\regfile/reg_out[12][14] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][14] ), .ZN(n2822) );
  AOI222_X1 U4417 ( .A1(\regfile/reg_out[27][14] ), .A2(n2333), .B1(
        \regfile/reg_out[23][14] ), .B2(n2334), .C1(\regfile/reg_out[22][14] ), 
        .C2(n2335), .ZN(n2812) );
  AOI222_X1 U4418 ( .A1(\regfile/reg_out[30][14] ), .A2(n2336), .B1(
        \regfile/reg_out[26][14] ), .B2(n2337), .C1(\regfile/reg_out[31][14] ), 
        .C2(n2338), .ZN(n2811) );
  OAI211_X1 U4419 ( .C1(n2823), .C2(n1557), .A(n2824), .B(n2825), .ZN(n7878)
         );
  AOI222_X1 U4420 ( .A1(n6102), .A2(n6521), .B1(
        \Mcontrol/Nextpc_decoding/Bta [13]), .B2(n7356), .C1(jar_in[13]), .C2(
        net57184), .ZN(n2825) );
  AOI22_X1 U4421 ( .A1(epc[13]), .A2(n1562), .B1(n1563), .B2(break_code[13]), 
        .ZN(n2824) );
  OAI22_X1 U4422 ( .A1(n2507), .A2(n2826), .B1(n6048), .B2(n2509), .ZN(
        break_code[13]) );
  NAND2_X1 U4423 ( .A1(\Mcontrol/d_sampled_finstr [13]), .A2(n7207), .ZN(n6048) );
  INV_X1 U4424 ( .A(n6346), .ZN(n2826) );
  INV_X1 U4425 ( .A(branch_rega[13]), .ZN(n2823) );
  INV_X1 U4427 ( .A(n794), .ZN(n2827) );
  NAND4_X1 U4428 ( .A1(n2828), .A2(n2829), .A3(n2830), .A4(n2831), .ZN(n794)
         );
  NOR4_X1 U4429 ( .A1(n2832), .A2(n2833), .A3(n2834), .A4(n2835), .ZN(n2831)
         );
  NAND3_X1 U4430 ( .A1(n6350), .A2(n6349), .A3(n6351), .ZN(n2835) );
  OAI211_X1 U4431 ( .C1(n5654), .C2(n796), .A(n6347), .B(n6348), .ZN(n2834) );
  OAI222_X1 U4433 ( .A1(n5652), .A2(n800), .B1(n7519), .B2(n799), .C1(n7482), 
        .C2(n795), .ZN(n2833) );
  OAI221_X1 U4437 ( .B1(n5646), .B2(n813), .C1(n5647), .C2(n812), .A(n2836), 
        .ZN(n2832) );
  AOI22_X1 U4438 ( .A1(\regfile/reg_out[2][13] ), .A2(n7642), .B1(
        \regfile/reg_out[3][13] ), .B2(n2323), .ZN(n2836) );
  AOI211_X1 U4441 ( .C1(\regfile/reg_out[16][13] ), .C2(n2324), .A(n2837), .B(
        n2838), .ZN(n2830) );
  OAI22_X1 U4442 ( .A1(n5624), .A2(n802), .B1(n815), .B2(n2327), .ZN(n2838) );
  OAI221_X1 U4445 ( .B1(n803), .B2(n2328), .C1(n814), .C2(n2329), .A(n2839), 
        .ZN(n2837) );
  AOI22_X1 U4446 ( .A1(n2331), .A2(\regfile/reg_out[12][13] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][13] ), .ZN(n2839) );
  AOI222_X1 U4449 ( .A1(\regfile/reg_out[27][13] ), .A2(n2333), .B1(
        \regfile/reg_out[23][13] ), .B2(n2334), .C1(\regfile/reg_out[22][13] ), 
        .C2(n2335), .ZN(n2829) );
  AOI222_X1 U4450 ( .A1(\regfile/reg_out[30][13] ), .A2(n2336), .B1(
        \regfile/reg_out[26][13] ), .B2(n2337), .C1(\regfile/reg_out[31][13] ), 
        .C2(n2338), .ZN(n2828) );
  OAI211_X1 U4451 ( .C1(n2840), .C2(n1557), .A(n2841), .B(n2842), .ZN(n7879)
         );
  AOI222_X1 U4452 ( .A1(n6102), .A2(n6519), .B1(
        \Mcontrol/Nextpc_decoding/Bta [12]), .B2(n7356), .C1(jar_in[12]), .C2(
        net57184), .ZN(n2842) );
  AOI22_X1 U4453 ( .A1(epc[12]), .A2(n1562), .B1(n1563), .B2(break_code[12]), 
        .ZN(n2841) );
  OAI22_X1 U4454 ( .A1(n2507), .A2(n2843), .B1(n6050), .B2(n2509), .ZN(
        break_code[12]) );
  NAND2_X1 U4455 ( .A1(\Mcontrol/d_sampled_finstr [12]), .A2(n7207), .ZN(n6050) );
  INV_X1 U4456 ( .A(n6358), .ZN(n2843) );
  INV_X1 U4457 ( .A(branch_rega[12]), .ZN(n2840) );
  INV_X1 U4459 ( .A(n756), .ZN(n2844) );
  NAND4_X1 U4460 ( .A1(n2845), .A2(n2846), .A3(n2847), .A4(n2848), .ZN(n756)
         );
  NAND3_X1 U4462 ( .A1(n6362), .A2(n6361), .A3(n6363), .ZN(n2852) );
  OAI211_X1 U4463 ( .C1(n5654), .C2(n758), .A(n6359), .B(n6360), .ZN(n2851) );
  OAI222_X1 U4465 ( .A1(n5652), .A2(n762), .B1(n7518), .B2(n761), .C1(n7484), 
        .C2(n757), .ZN(n2850) );
  OAI221_X1 U4469 ( .B1(n5646), .B2(n775), .C1(n5647), .C2(n774), .A(n2853), 
        .ZN(n2849) );
  AOI22_X1 U4470 ( .A1(\regfile/reg_out[2][12] ), .A2(n7641), .B1(
        \regfile/reg_out[3][12] ), .B2(n2323), .ZN(n2853) );
  AOI211_X1 U4473 ( .C1(\regfile/reg_out[16][12] ), .C2(n2324), .A(n2854), .B(
        n2855), .ZN(n2847) );
  OAI22_X1 U4474 ( .A1(n5624), .A2(n764), .B1(n777), .B2(n2327), .ZN(n2855) );
  OAI221_X1 U4477 ( .B1(n765), .B2(n2328), .C1(n776), .C2(n2329), .A(n2856), 
        .ZN(n2854) );
  AOI22_X1 U4478 ( .A1(n2331), .A2(\regfile/reg_out[12][12] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][12] ), .ZN(n2856) );
  AOI222_X1 U4481 ( .A1(\regfile/reg_out[27][12] ), .A2(n2333), .B1(
        \regfile/reg_out[23][12] ), .B2(n2334), .C1(\regfile/reg_out[22][12] ), 
        .C2(n2335), .ZN(n2846) );
  AOI222_X1 U4482 ( .A1(\regfile/reg_out[30][12] ), .A2(n2336), .B1(
        \regfile/reg_out[26][12] ), .B2(n2337), .C1(\regfile/reg_out[31][12] ), 
        .C2(n2338), .ZN(n2845) );
  OAI211_X1 U4483 ( .C1(n2857), .C2(n1557), .A(n2858), .B(n2859), .ZN(n7880)
         );
  AOI22_X1 U4485 ( .A1(epc[11]), .A2(n1562), .B1(n1563), .B2(break_code[11]), 
        .ZN(n2858) );
  NAND2_X1 U4487 ( .A1(\Mcontrol/d_sampled_finstr [11]), .A2(n7207), .ZN(n6051) );
  INV_X1 U4488 ( .A(n6370), .ZN(n2860) );
  INV_X1 U4489 ( .A(branch_rega[11]), .ZN(n2857) );
  INV_X1 U4491 ( .A(n718), .ZN(n2861) );
  NAND4_X1 U4492 ( .A1(n2862), .A2(n2863), .A3(n2864), .A4(n2865), .ZN(n718)
         );
  NAND3_X1 U4494 ( .A1(n6374), .A2(n6373), .A3(n6375), .ZN(n2869) );
  OAI211_X1 U4495 ( .C1(n5654), .C2(n720), .A(n6371), .B(n6372), .ZN(n2868) );
  OAI222_X1 U4497 ( .A1(n5652), .A2(n724), .B1(n7519), .B2(n723), .C1(n7484), 
        .C2(n719), .ZN(n2867) );
  OAI221_X1 U4501 ( .B1(n5646), .B2(n737), .C1(n5647), .C2(n736), .A(n2870), 
        .ZN(n2866) );
  AOI22_X1 U4502 ( .A1(\regfile/reg_out[2][11] ), .A2(n7642), .B1(
        \regfile/reg_out[3][11] ), .B2(n2323), .ZN(n2870) );
  AOI211_X1 U4505 ( .C1(\regfile/reg_out[16][11] ), .C2(n2324), .A(n2871), .B(
        n2872), .ZN(n2864) );
  OAI22_X1 U4506 ( .A1(n5624), .A2(n726), .B1(n739), .B2(n2327), .ZN(n2872) );
  OAI221_X1 U4509 ( .B1(n727), .B2(n2328), .C1(n738), .C2(n2329), .A(n2873), 
        .ZN(n2871) );
  AOI22_X1 U4510 ( .A1(n2331), .A2(\regfile/reg_out[12][11] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][11] ), .ZN(n2873) );
  AOI222_X1 U4513 ( .A1(\regfile/reg_out[27][11] ), .A2(n2333), .B1(
        \regfile/reg_out[23][11] ), .B2(n2334), .C1(\regfile/reg_out[22][11] ), 
        .C2(n2335), .ZN(n2863) );
  AOI222_X1 U4514 ( .A1(\regfile/reg_out[30][11] ), .A2(n2336), .B1(
        \regfile/reg_out[26][11] ), .B2(n2337), .C1(\regfile/reg_out[31][11] ), 
        .C2(n2338), .ZN(n2862) );
  OAI211_X1 U4515 ( .C1(n2874), .C2(n1557), .A(n2875), .B(n2876), .ZN(n7881)
         );
  AOI22_X1 U4519 ( .A1(epc[10]), .A2(n1562), .B1(n1563), .B2(break_code[10]), 
        .ZN(n2875) );
  OAI22_X1 U4520 ( .A1(n2507), .A2(n2879), .B1(n5894), .B2(n2509), .ZN(
        break_code[10]) );
  AOI21_X1 U4522 ( .B1(n7450), .B2(n6105), .A(n2792), .ZN(n2880) );
  NAND2_X1 U4534 ( .A1(\Mcontrol/d_sampled_finstr [10]), .A2(n7207), .ZN(n5894) );
  INV_X1 U4535 ( .A(n6383), .ZN(n2879) );
  NAND3_X1 U4536 ( .A1(net57341), .A2(n7430), .A3(n6105), .ZN(n2507) );
  INV_X1 U4538 ( .A(n7505), .ZN(\Mcontrol/Operation_decoding32/N1982 ) );
  INV_X1 U4542 ( .A(\Mcontrol/Nextpc_decoding/N171 ), .ZN(n2878) );
  INV_X1 U4543 ( .A(n6397), .ZN(n2877) );
  INV_X1 U4548 ( .A(branch_rega[10]), .ZN(n2874) );
  OAI222_X1 U4549 ( .A1(n5623), .A2(n5617), .B1(n7486), .B2(n2883), .C1(n5621), 
        .C2(n5615), .ZN(branch_rega[10]) );
  INV_X1 U4550 ( .A(n680), .ZN(n2883) );
  NAND4_X1 U4551 ( .A1(n2884), .A2(n2885), .A3(n2886), .A4(n2887), .ZN(n680)
         );
  NOR4_X1 U4552 ( .A1(n2888), .A2(n2889), .A3(n2890), .A4(n2891), .ZN(n2887)
         );
  NAND3_X1 U4553 ( .A1(n6388), .A2(n6387), .A3(n6389), .ZN(n2891) );
  OAI211_X1 U4554 ( .C1(n5654), .C2(n682), .A(n6385), .B(n6386), .ZN(n2890) );
  OAI222_X1 U4556 ( .A1(n5652), .A2(n686), .B1(n7518), .B2(n685), .C1(n7482), 
        .C2(n681), .ZN(n2889) );
  OAI221_X1 U4560 ( .B1(n5646), .B2(n699), .C1(n5647), .C2(n698), .A(n2892), 
        .ZN(n2888) );
  AOI22_X1 U4561 ( .A1(\regfile/reg_out[2][10] ), .A2(n7642), .B1(
        \regfile/reg_out[3][10] ), .B2(n2323), .ZN(n2892) );
  AOI211_X1 U4566 ( .C1(\regfile/reg_out[16][10] ), .C2(n2324), .A(n2893), .B(
        n2894), .ZN(n2886) );
  OAI22_X1 U4567 ( .A1(n5624), .A2(n688), .B1(n701), .B2(n2327), .ZN(n2894) );
  OAI221_X1 U4571 ( .B1(n689), .B2(n2328), .C1(n700), .C2(n2329), .A(n2895), 
        .ZN(n2893) );
  AOI22_X1 U4572 ( .A1(n2331), .A2(\regfile/reg_out[12][10] ), .B1(n2332), 
        .B2(\regfile/reg_out[13][10] ), .ZN(n2895) );
  INV_X1 U4576 ( .A(rs1_addr[4]), .ZN(n2896) );
  AOI222_X1 U4582 ( .A1(\regfile/reg_out[27][10] ), .A2(n2333), .B1(
        \regfile/reg_out[23][10] ), .B2(n2334), .C1(\regfile/reg_out[22][10] ), 
        .C2(n2335), .ZN(n2885) );
  AOI222_X1 U4586 ( .A1(\regfile/reg_out[30][10] ), .A2(n2336), .B1(
        \regfile/reg_out[26][10] ), .B2(n2337), .C1(\regfile/reg_out[31][10] ), 
        .C2(n2338), .ZN(n2884) );
  INV_X1 U4613 ( .A(\Scc_coproc/interrupt[2] ), .ZN(n6492) );
  INV_X1 U4614 ( .A(n4506), .ZN(\x_mem_command[MW] ) );
  AND2_X1 U4618 ( .A1(\Mcontrol/m_sampled_xrd[1] ), .A2(n5503), .ZN(rd_addr[1]) );
  OAI21_X1 U4620 ( .B1(n4506), .B2(n7109), .A(n5504), .ZN(mem_write) );
  NOR2_X1 U4621 ( .A1(\Mcontrol/x_sampled_dmem_command[MW] ), .A2(
        \Mcontrol/x_sampled_dwe ), .ZN(n4506) );
  NOR2_X1 U4622 ( .A1(n4507), .A2(n7109), .ZN(mem_read) );
  OAI21_X1 U4623 ( .B1(n4508), .B2(n7109), .A(n5504), .ZN(mem_ishalf) );
  OAI21_X1 U4624 ( .B1(n5505), .B2(n7109), .A(n5504), .ZN(mem_isbyte) );
  INV_X1 U4625 ( .A(N80), .ZN(dcheck_enable) );
  OR2_X1 U4626 ( .A1(\Mcontrol/bp_logicB/memory_main ), .A2(
        \Mcontrol/bp_logicB/exec_main ), .ZN(byp_controlB[2]) );
  OAI222_X1 U4628 ( .A1(n5522), .A2(n5523), .B1(n5524), .B2(n5525), .C1(n5526), 
        .C2(n5527), .ZN(branch_regb[9]) );
  OAI222_X1 U4629 ( .A1(n5528), .A2(n5523), .B1(n5529), .B2(n5525), .C1(n5530), 
        .C2(n5527), .ZN(branch_regb[8]) );
  OAI222_X1 U4630 ( .A1(n5531), .A2(n5523), .B1(n5532), .B2(n5525), .C1(n5533), 
        .C2(n5527), .ZN(branch_regb[7]) );
  OAI222_X1 U4632 ( .A1(n5537), .A2(n5523), .B1(n5538), .B2(n5525), .C1(n5539), 
        .C2(n5527), .ZN(branch_regb[5]) );
  OAI222_X1 U4633 ( .A1(n5540), .A2(n5523), .B1(n5541), .B2(n5525), .C1(n5542), 
        .C2(n5527), .ZN(branch_regb[4]) );
  OAI222_X1 U4634 ( .A1(n5543), .A2(n5523), .B1(n5544), .B2(n5525), .C1(n5545), 
        .C2(n5527), .ZN(branch_regb[3]) );
  OAI222_X1 U4637 ( .A1(n5552), .A2(n5523), .B1(n5553), .B2(n5525), .C1(n5554), 
        .C2(n5527), .ZN(branch_regb[2]) );
  OAI222_X1 U4638 ( .A1(n5555), .A2(n5523), .B1(n5556), .B2(n5525), .C1(n5557), 
        .C2(n5527), .ZN(branch_regb[29]) );
  OAI222_X1 U4642 ( .A1(n5567), .A2(n5523), .B1(n5568), .B2(n5525), .C1(n5569), 
        .C2(n5527), .ZN(branch_regb[25]) );
  OAI222_X1 U4643 ( .A1(n5570), .A2(n5523), .B1(n5571), .B2(n5525), .C1(n5572), 
        .C2(n5527), .ZN(branch_regb[24]) );
  OAI222_X1 U4644 ( .A1(n5573), .A2(n5523), .B1(n5574), .B2(n5525), .C1(n5575), 
        .C2(n5527), .ZN(branch_regb[23]) );
  OAI222_X1 U4646 ( .A1(n5579), .A2(n5523), .B1(n5580), .B2(n5525), .C1(n5581), 
        .C2(n5527), .ZN(branch_regb[21]) );
  OAI222_X1 U4647 ( .A1(n5582), .A2(n5523), .B1(n5583), .B2(n5525), .C1(n5584), 
        .C2(n5527), .ZN(branch_regb[20]) );
  OAI222_X1 U4648 ( .A1(n5585), .A2(n5523), .B1(n5586), .B2(n5525), .C1(n5587), 
        .C2(n5527), .ZN(branch_regb[1]) );
  OAI222_X1 U4649 ( .A1(n5588), .A2(n5523), .B1(n5589), .B2(n5525), .C1(n5590), 
        .C2(n5527), .ZN(branch_regb[19]) );
  OAI222_X1 U4650 ( .A1(n5591), .A2(n5523), .B1(n5592), .B2(n5525), .C1(n5593), 
        .C2(n5527), .ZN(branch_regb[18]) );
  OAI222_X1 U4651 ( .A1(n5594), .A2(n5523), .B1(n5595), .B2(n5525), .C1(n5596), 
        .C2(n5527), .ZN(branch_regb[17]) );
  OAI222_X1 U4652 ( .A1(n5597), .A2(n5523), .B1(n5598), .B2(n5525), .C1(n5599), 
        .C2(n5527), .ZN(branch_regb[16]) );
  OAI222_X1 U4653 ( .A1(n5600), .A2(n5523), .B1(n5601), .B2(n5525), .C1(n5602), 
        .C2(n5527), .ZN(branch_regb[15]) );
  OAI222_X1 U4654 ( .A1(n5603), .A2(n5523), .B1(n5604), .B2(n5525), .C1(n5605), 
        .C2(n5527), .ZN(branch_regb[14]) );
  OAI222_X1 U4655 ( .A1(n5606), .A2(n5523), .B1(n5607), .B2(n5525), .C1(n5608), 
        .C2(n5527), .ZN(branch_regb[13]) );
  OAI222_X1 U4656 ( .A1(n5609), .A2(n5523), .B1(n5610), .B2(n5525), .C1(n5611), 
        .C2(n5527), .ZN(branch_regb[12]) );
  OAI222_X1 U4657 ( .A1(n5612), .A2(n5523), .B1(n5613), .B2(n5525), .C1(n5614), 
        .C2(n5527), .ZN(branch_regb[11]) );
  OAI222_X1 U4659 ( .A1(n5618), .A2(n5523), .B1(n5619), .B2(n5525), .C1(n5620), 
        .C2(n5527), .ZN(branch_regb[0]) );
  AOI22_X1 U4664 ( .A1(n5627), .A2(\regfile/reg_out[19][30] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][30] ), .ZN(n5626) );
  AOI22_X1 U4665 ( .A1(n7501), .A2(\regfile/reg_out[21][30] ), .B1(n5633), 
        .B2(\regfile/reg_out[20][30] ), .ZN(n5631) );
  AOI22_X1 U4666 ( .A1(n5637), .A2(\regfile/reg_out[25][30] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][30] ), .ZN(n5636) );
  AOI22_X1 U4667 ( .A1(n5642), .A2(\regfile/reg_out[29][30] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][30] ), .ZN(n5641) );
  AOI22_X1 U4668 ( .A1(n5649), .A2(\regfile/reg_out[5][30] ), .B1(n5650), .B2(
        \regfile/reg_out[4][30] ), .ZN(n5648) );
  OAI222_X1 U4671 ( .A1(n5555), .A2(n5621), .B1(n5508), .B2(n7487), .C1(n5557), 
        .C2(n5623), .ZN(branch_rega[29]) );
  AOI22_X1 U4672 ( .A1(n7603), .A2(\regfile/reg_out[19][29] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][29] ), .ZN(n5660) );
  AOI22_X1 U4673 ( .A1(n7502), .A2(\regfile/reg_out[21][29] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][29] ), .ZN(n5661) );
  AOI22_X1 U4674 ( .A1(n5637), .A2(\regfile/reg_out[25][29] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][29] ), .ZN(n5662) );
  AOI22_X1 U4675 ( .A1(n5642), .A2(\regfile/reg_out[29][29] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][29] ), .ZN(n5663) );
  AOI22_X1 U4676 ( .A1(n5649), .A2(\regfile/reg_out[5][29] ), .B1(n5650), .B2(
        \regfile/reg_out[4][29] ), .ZN(n5664) );
  INV_X1 U4677 ( .A(n5665), .ZN(n5555) );
  OAI22_X1 U4678 ( .A1(n5666), .A2(n5657), .B1(n5667), .B2(n5659), .ZN(n5665)
         );
  AOI22_X1 U4680 ( .A1(n7603), .A2(\regfile/reg_out[19][28] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][28] ), .ZN(n5668) );
  AOI22_X1 U4681 ( .A1(n7502), .A2(\regfile/reg_out[21][28] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][28] ), .ZN(n5669) );
  AOI22_X1 U4682 ( .A1(n5637), .A2(\regfile/reg_out[25][28] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][28] ), .ZN(n5670) );
  AOI22_X1 U4683 ( .A1(n5642), .A2(\regfile/reg_out[29][28] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][28] ), .ZN(n5671) );
  AOI22_X1 U4684 ( .A1(n5649), .A2(\regfile/reg_out[5][28] ), .B1(n5650), .B2(
        \regfile/reg_out[4][28] ), .ZN(n5672) );
  INV_X1 U4685 ( .A(n5673), .ZN(n5558) );
  OAI22_X1 U4686 ( .A1(n5674), .A2(n5657), .B1(n5675), .B2(n5659), .ZN(n5673)
         );
  AOI22_X1 U4688 ( .A1(n7603), .A2(\regfile/reg_out[19][27] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][27] ), .ZN(n5676) );
  AOI22_X1 U4689 ( .A1(n7503), .A2(\regfile/reg_out[21][27] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][27] ), .ZN(n5677) );
  AOI22_X1 U4690 ( .A1(n5637), .A2(\regfile/reg_out[25][27] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][27] ), .ZN(n5678) );
  AOI22_X1 U4691 ( .A1(n5642), .A2(\regfile/reg_out[29][27] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][27] ), .ZN(n5679) );
  AOI22_X1 U4692 ( .A1(n5649), .A2(\regfile/reg_out[5][27] ), .B1(n5650), .B2(
        \regfile/reg_out[4][27] ), .ZN(n5680) );
  INV_X1 U4693 ( .A(n5681), .ZN(n5561) );
  OAI22_X1 U4694 ( .A1(n5682), .A2(n5657), .B1(n5683), .B2(n5659), .ZN(n5681)
         );
  OAI222_X1 U4695 ( .A1(n5564), .A2(n5621), .B1(n5511), .B2(n7486), .C1(n5566), 
        .C2(n5623), .ZN(branch_rega[26]) );
  AOI22_X1 U4696 ( .A1(n7603), .A2(\regfile/reg_out[19][26] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][26] ), .ZN(n5684) );
  AOI22_X1 U4697 ( .A1(n7502), .A2(\regfile/reg_out[21][26] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][26] ), .ZN(n5685) );
  AOI22_X1 U4698 ( .A1(n5637), .A2(\regfile/reg_out[25][26] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][26] ), .ZN(n5686) );
  AOI22_X1 U4699 ( .A1(n5642), .A2(\regfile/reg_out[29][26] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][26] ), .ZN(n5687) );
  AOI22_X1 U4700 ( .A1(n5649), .A2(\regfile/reg_out[5][26] ), .B1(n5650), .B2(
        \regfile/reg_out[4][26] ), .ZN(n5688) );
  INV_X1 U4701 ( .A(n5689), .ZN(n5564) );
  OAI22_X1 U4702 ( .A1(n5690), .A2(n5657), .B1(n5691), .B2(n5659), .ZN(n5689)
         );
  AOI22_X1 U4704 ( .A1(n7603), .A2(\regfile/reg_out[19][25] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][25] ), .ZN(n5692) );
  AOI22_X1 U4705 ( .A1(n7503), .A2(\regfile/reg_out[21][25] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][25] ), .ZN(n5693) );
  AOI22_X1 U4706 ( .A1(n5637), .A2(\regfile/reg_out[25][25] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][25] ), .ZN(n5694) );
  AOI22_X1 U4707 ( .A1(n5642), .A2(\regfile/reg_out[29][25] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][25] ), .ZN(n5695) );
  AOI22_X1 U4708 ( .A1(n5649), .A2(\regfile/reg_out[5][25] ), .B1(n5650), .B2(
        \regfile/reg_out[4][25] ), .ZN(n5696) );
  INV_X1 U4709 ( .A(n5697), .ZN(n5567) );
  OAI22_X1 U4710 ( .A1(n5698), .A2(n5657), .B1(n5699), .B2(n5659), .ZN(n5697)
         );
  AOI22_X1 U4712 ( .A1(n7603), .A2(\regfile/reg_out[19][24] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][24] ), .ZN(n5700) );
  AOI22_X1 U4713 ( .A1(n7503), .A2(\regfile/reg_out[21][24] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][24] ), .ZN(n5701) );
  AOI22_X1 U4714 ( .A1(n5637), .A2(\regfile/reg_out[25][24] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][24] ), .ZN(n5702) );
  AOI22_X1 U4715 ( .A1(n5642), .A2(\regfile/reg_out[29][24] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][24] ), .ZN(n5703) );
  AOI22_X1 U4716 ( .A1(n5649), .A2(\regfile/reg_out[5][24] ), .B1(n5650), .B2(
        \regfile/reg_out[4][24] ), .ZN(n5704) );
  INV_X1 U4717 ( .A(n5705), .ZN(n5570) );
  OAI22_X1 U4718 ( .A1(n5706), .A2(n5657), .B1(n5707), .B2(n5659), .ZN(n5705)
         );
  AOI22_X1 U4720 ( .A1(n7603), .A2(\regfile/reg_out[19][0] ), .B1(n7621), .B2(
        \regfile/reg_out[18][0] ), .ZN(n5708) );
  AOI22_X1 U4721 ( .A1(n7503), .A2(\regfile/reg_out[21][0] ), .B1(n5633), .B2(
        \regfile/reg_out[20][0] ), .ZN(n5709) );
  AOI22_X1 U4722 ( .A1(n5637), .A2(\regfile/reg_out[25][0] ), .B1(n7096), .B2(
        \regfile/reg_out[24][0] ), .ZN(n5710) );
  AOI22_X1 U4723 ( .A1(n5642), .A2(\regfile/reg_out[29][0] ), .B1(n5643), .B2(
        \regfile/reg_out[28][0] ), .ZN(n5711) );
  AOI22_X1 U4724 ( .A1(n5649), .A2(\regfile/reg_out[5][0] ), .B1(n5650), .B2(
        \regfile/reg_out[4][0] ), .ZN(n5712) );
  INV_X1 U4725 ( .A(n5713), .ZN(n5618) );
  OAI221_X1 U4726 ( .B1(n5714), .B2(n5659), .C1(n5715), .C2(n5657), .A(n5716), 
        .ZN(n5713) );
  INV_X1 U4728 ( .A(n5720), .ZN(n5717) );
  AOI22_X1 U4729 ( .A1(n5752), .A2(\regfile/reg_out[19][9] ), .B1(n5753), .B2(
        \regfile/reg_out[18][9] ), .ZN(n5751) );
  AOI22_X1 U4730 ( .A1(n5757), .A2(\regfile/reg_out[21][9] ), .B1(n5758), .B2(
        \regfile/reg_out[20][9] ), .ZN(n5756) );
  AOI22_X1 U4731 ( .A1(n5762), .A2(\regfile/reg_out[25][9] ), .B1(n5763), .B2(
        \regfile/reg_out[24][9] ), .ZN(n5761) );
  AOI22_X1 U4732 ( .A1(n5767), .A2(\regfile/reg_out[29][9] ), .B1(n5768), .B2(
        \regfile/reg_out[28][9] ), .ZN(n5766) );
  AOI22_X1 U4733 ( .A1(n5774), .A2(\regfile/reg_out[5][9] ), .B1(n5775), .B2(
        \regfile/reg_out[4][9] ), .ZN(n5773) );
  AOI22_X1 U4734 ( .A1(n5752), .A2(\regfile/reg_out[19][8] ), .B1(n5753), .B2(
        \regfile/reg_out[18][8] ), .ZN(n5780) );
  AOI22_X1 U4735 ( .A1(n5757), .A2(\regfile/reg_out[21][8] ), .B1(n5758), .B2(
        \regfile/reg_out[20][8] ), .ZN(n5781) );
  AOI22_X1 U4736 ( .A1(n5762), .A2(\regfile/reg_out[25][8] ), .B1(n5763), .B2(
        \regfile/reg_out[24][8] ), .ZN(n5782) );
  AOI22_X1 U4737 ( .A1(n5767), .A2(\regfile/reg_out[29][8] ), .B1(n5768), .B2(
        \regfile/reg_out[28][8] ), .ZN(n5783) );
  AOI22_X1 U4738 ( .A1(n5774), .A2(\regfile/reg_out[5][8] ), .B1(n5775), .B2(
        \regfile/reg_out[4][8] ), .ZN(n5784) );
  OAI22_X1 U4739 ( .A1(n5789), .A2(n5790), .B1(n5791), .B2(n5792), .ZN(n5788)
         );
  AOI22_X1 U4740 ( .A1(n5752), .A2(\regfile/reg_out[19][7] ), .B1(n5753), .B2(
        \regfile/reg_out[18][7] ), .ZN(n5793) );
  AOI22_X1 U4741 ( .A1(n5757), .A2(\regfile/reg_out[21][7] ), .B1(n5758), .B2(
        \regfile/reg_out[20][7] ), .ZN(n5794) );
  AOI22_X1 U4742 ( .A1(n5762), .A2(\regfile/reg_out[25][7] ), .B1(n5763), .B2(
        \regfile/reg_out[24][7] ), .ZN(n5795) );
  AOI22_X1 U4743 ( .A1(n5767), .A2(\regfile/reg_out[29][7] ), .B1(n5768), .B2(
        \regfile/reg_out[28][7] ), .ZN(n5796) );
  AOI22_X1 U4744 ( .A1(n5774), .A2(\regfile/reg_out[5][7] ), .B1(n5775), .B2(
        \regfile/reg_out[4][7] ), .ZN(n5797) );
  OAI22_X1 U4745 ( .A1(n5790), .A2(n5799), .B1(n5792), .B2(n5800), .ZN(n5798)
         );
  OAI22_X1 U4746 ( .A1(n5802), .A2(n5803), .B1(n5804), .B2(n5799), .ZN(n5801)
         );
  AOI22_X1 U4747 ( .A1(n5752), .A2(\regfile/reg_out[19][6] ), .B1(n5753), .B2(
        \regfile/reg_out[18][6] ), .ZN(n5805) );
  AOI22_X1 U4748 ( .A1(n5757), .A2(\regfile/reg_out[21][6] ), .B1(n5758), .B2(
        \regfile/reg_out[20][6] ), .ZN(n5806) );
  AOI22_X1 U4749 ( .A1(n5762), .A2(\regfile/reg_out[25][6] ), .B1(n5763), .B2(
        \regfile/reg_out[24][6] ), .ZN(n5807) );
  AOI22_X1 U4750 ( .A1(n5767), .A2(\regfile/reg_out[29][6] ), .B1(n5768), .B2(
        \regfile/reg_out[28][6] ), .ZN(n5808) );
  AOI22_X1 U4751 ( .A1(n5774), .A2(\regfile/reg_out[5][6] ), .B1(n5775), .B2(
        \regfile/reg_out[4][6] ), .ZN(n5809) );
  OAI22_X1 U4752 ( .A1(n5790), .A2(n5811), .B1(n5792), .B2(n5812), .ZN(n5810)
         );
  OAI22_X1 U4753 ( .A1(n5802), .A2(n5814), .B1(n5804), .B2(n5811), .ZN(n5813)
         );
  AOI22_X1 U4754 ( .A1(n5752), .A2(\regfile/reg_out[19][5] ), .B1(n5753), .B2(
        \regfile/reg_out[18][5] ), .ZN(n5815) );
  AOI22_X1 U4755 ( .A1(n5757), .A2(\regfile/reg_out[21][5] ), .B1(n5758), .B2(
        \regfile/reg_out[20][5] ), .ZN(n5816) );
  AOI22_X1 U4756 ( .A1(n5762), .A2(\regfile/reg_out[25][5] ), .B1(n5763), .B2(
        \regfile/reg_out[24][5] ), .ZN(n5817) );
  AOI22_X1 U4757 ( .A1(n5767), .A2(\regfile/reg_out[29][5] ), .B1(n5768), .B2(
        \regfile/reg_out[28][5] ), .ZN(n5818) );
  AOI22_X1 U4758 ( .A1(n5774), .A2(\regfile/reg_out[5][5] ), .B1(n5775), .B2(
        \regfile/reg_out[4][5] ), .ZN(n5819) );
  OAI22_X1 U4759 ( .A1(n5790), .A2(n5821), .B1(n5792), .B2(n5822), .ZN(n5820)
         );
  OAI22_X1 U4760 ( .A1(n5802), .A2(n5824), .B1(n5804), .B2(n5821), .ZN(n5823)
         );
  AOI22_X1 U4761 ( .A1(n5752), .A2(\regfile/reg_out[19][4] ), .B1(n5753), .B2(
        \regfile/reg_out[18][4] ), .ZN(n5825) );
  AOI22_X1 U4762 ( .A1(n5757), .A2(\regfile/reg_out[21][4] ), .B1(n5758), .B2(
        \regfile/reg_out[20][4] ), .ZN(n5826) );
  AOI22_X1 U4763 ( .A1(n5762), .A2(\regfile/reg_out[25][4] ), .B1(n5763), .B2(
        \regfile/reg_out[24][4] ), .ZN(n5827) );
  AOI22_X1 U4764 ( .A1(n5767), .A2(\regfile/reg_out[29][4] ), .B1(n5768), .B2(
        \regfile/reg_out[28][4] ), .ZN(n5828) );
  AOI22_X1 U4765 ( .A1(n5774), .A2(\regfile/reg_out[5][4] ), .B1(n5775), .B2(
        \regfile/reg_out[4][4] ), .ZN(n5829) );
  OAI22_X1 U4766 ( .A1(n5790), .A2(n5831), .B1(n5792), .B2(n5832), .ZN(n5830)
         );
  OAI22_X1 U4767 ( .A1(n5802), .A2(n5834), .B1(n5804), .B2(n5831), .ZN(n5833)
         );
  AOI22_X1 U4768 ( .A1(n5752), .A2(\regfile/reg_out[19][3] ), .B1(n5753), .B2(
        \regfile/reg_out[18][3] ), .ZN(n5835) );
  AOI22_X1 U4769 ( .A1(n5757), .A2(\regfile/reg_out[21][3] ), .B1(n5758), .B2(
        \regfile/reg_out[20][3] ), .ZN(n5836) );
  AOI22_X1 U4770 ( .A1(n5762), .A2(\regfile/reg_out[25][3] ), .B1(n5763), .B2(
        \regfile/reg_out[24][3] ), .ZN(n5837) );
  AOI22_X1 U4771 ( .A1(n5767), .A2(\regfile/reg_out[29][3] ), .B1(n5768), .B2(
        \regfile/reg_out[28][3] ), .ZN(n5838) );
  AOI22_X1 U4772 ( .A1(n5774), .A2(\regfile/reg_out[5][3] ), .B1(n5775), .B2(
        \regfile/reg_out[4][3] ), .ZN(n5839) );
  AOI22_X1 U4773 ( .A1(n5752), .A2(\regfile/reg_out[19][31] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][31] ), .ZN(n5840) );
  AOI22_X1 U4774 ( .A1(n5757), .A2(\regfile/reg_out[21][31] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][31] ), .ZN(n5841) );
  AOI22_X1 U4775 ( .A1(n5762), .A2(\regfile/reg_out[25][31] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][31] ), .ZN(n5842) );
  AOI22_X1 U4776 ( .A1(n5767), .A2(\regfile/reg_out[29][31] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][31] ), .ZN(n5843) );
  AOI22_X1 U4777 ( .A1(n5774), .A2(\regfile/reg_out[5][31] ), .B1(n5775), .B2(
        \regfile/reg_out[4][31] ), .ZN(n5844) );
  OAI21_X1 U4778 ( .B1(n5846), .B2(n5847), .A(n5848), .ZN(n5845) );
  AOI22_X1 U4779 ( .A1(n5752), .A2(\regfile/reg_out[19][30] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][30] ), .ZN(n5849) );
  AOI22_X1 U4780 ( .A1(n5757), .A2(\regfile/reg_out[21][30] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][30] ), .ZN(n5850) );
  AOI22_X1 U4781 ( .A1(n5762), .A2(\regfile/reg_out[25][30] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][30] ), .ZN(n5851) );
  AOI22_X1 U4782 ( .A1(n5767), .A2(\regfile/reg_out[29][30] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][30] ), .ZN(n5852) );
  AOI22_X1 U4783 ( .A1(n5774), .A2(\regfile/reg_out[5][30] ), .B1(n5775), .B2(
        \regfile/reg_out[4][30] ), .ZN(n5853) );
  OAI22_X1 U4784 ( .A1(n5790), .A2(n5856), .B1(n5792), .B2(n5857), .ZN(n5855)
         );
  OAI22_X1 U4785 ( .A1(n5802), .A2(n5859), .B1(n5804), .B2(n5856), .ZN(n5858)
         );
  INV_X1 U4786 ( .A(\Mpath/the_memhandle/N38 ), .ZN(n5804) );
  AOI22_X1 U4787 ( .A1(n5752), .A2(\regfile/reg_out[19][2] ), .B1(n5753), .B2(
        \regfile/reg_out[18][2] ), .ZN(n5860) );
  AOI22_X1 U4788 ( .A1(n5757), .A2(\regfile/reg_out[21][2] ), .B1(n5758), .B2(
        \regfile/reg_out[20][2] ), .ZN(n5861) );
  AOI22_X1 U4789 ( .A1(n5762), .A2(\regfile/reg_out[25][2] ), .B1(n5763), .B2(
        \regfile/reg_out[24][2] ), .ZN(n5862) );
  AOI22_X1 U4790 ( .A1(n5767), .A2(\regfile/reg_out[29][2] ), .B1(n5768), .B2(
        \regfile/reg_out[28][2] ), .ZN(n5863) );
  AOI22_X1 U4791 ( .A1(n5774), .A2(\regfile/reg_out[5][2] ), .B1(n5775), .B2(
        \regfile/reg_out[4][2] ), .ZN(n5864) );
  AOI22_X1 U4792 ( .A1(n5752), .A2(\regfile/reg_out[19][29] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][29] ), .ZN(n5865) );
  AOI22_X1 U4793 ( .A1(n5757), .A2(\regfile/reg_out[21][29] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][29] ), .ZN(n5866) );
  AOI22_X1 U4794 ( .A1(n5762), .A2(\regfile/reg_out[25][29] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][29] ), .ZN(n5867) );
  AOI22_X1 U4795 ( .A1(n5767), .A2(\regfile/reg_out[29][29] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][29] ), .ZN(n5868) );
  AOI22_X1 U4796 ( .A1(n5774), .A2(\regfile/reg_out[5][29] ), .B1(n5775), .B2(
        \regfile/reg_out[4][29] ), .ZN(n5869) );
  AOI22_X1 U4797 ( .A1(n5752), .A2(\regfile/reg_out[19][28] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][28] ), .ZN(n5870) );
  AOI22_X1 U4798 ( .A1(n5757), .A2(\regfile/reg_out[21][28] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][28] ), .ZN(n5871) );
  AOI22_X1 U4799 ( .A1(n5762), .A2(\regfile/reg_out[25][28] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][28] ), .ZN(n5872) );
  AOI22_X1 U4800 ( .A1(n5767), .A2(\regfile/reg_out[29][28] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][28] ), .ZN(n5873) );
  AOI22_X1 U4801 ( .A1(n5774), .A2(\regfile/reg_out[5][28] ), .B1(n5775), .B2(
        \regfile/reg_out[4][28] ), .ZN(n5874) );
  AOI22_X1 U4802 ( .A1(n5752), .A2(\regfile/reg_out[19][27] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][27] ), .ZN(n5875) );
  AOI22_X1 U4803 ( .A1(n5757), .A2(\regfile/reg_out[21][27] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][27] ), .ZN(n5876) );
  AOI22_X1 U4804 ( .A1(n5762), .A2(\regfile/reg_out[25][27] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][27] ), .ZN(n5877) );
  AOI22_X1 U4805 ( .A1(n5767), .A2(\regfile/reg_out[29][27] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][27] ), .ZN(n5878) );
  AOI22_X1 U4806 ( .A1(n5774), .A2(\regfile/reg_out[5][27] ), .B1(n5775), .B2(
        \regfile/reg_out[4][27] ), .ZN(n5879) );
  NAND2_X1 U4807 ( .A1(n5880), .A2(n5848), .ZN(n5854) );
  OAI21_X1 U4808 ( .B1(n5881), .B2(n5882), .A(n5847), .ZN(n5848) );
  NOR2_X1 U4809 ( .A1(n5883), .A2(n5884), .ZN(n5881) );
  AOI22_X1 U4810 ( .A1(n5752), .A2(\regfile/reg_out[19][26] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][26] ), .ZN(n5885) );
  AOI22_X1 U4811 ( .A1(n5757), .A2(\regfile/reg_out[21][26] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][26] ), .ZN(n5886) );
  AOI22_X1 U4812 ( .A1(n5762), .A2(\regfile/reg_out[25][26] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][26] ), .ZN(n5887) );
  AOI22_X1 U4813 ( .A1(n5767), .A2(\regfile/reg_out[29][26] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][26] ), .ZN(n5888) );
  AOI22_X1 U4814 ( .A1(n5774), .A2(\regfile/reg_out[5][26] ), .B1(n5775), .B2(
        \regfile/reg_out[4][26] ), .ZN(n5889) );
  OAI21_X1 U4815 ( .B1(n5892), .B2(n5884), .A(n5893), .ZN(n5891) );
  INV_X1 U4816 ( .A(n5894), .ZN(n5890) );
  AOI22_X1 U4817 ( .A1(n5752), .A2(\regfile/reg_out[19][25] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][25] ), .ZN(n5896) );
  AOI22_X1 U4818 ( .A1(n5757), .A2(\regfile/reg_out[21][25] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][25] ), .ZN(n5897) );
  AOI22_X1 U4819 ( .A1(n5762), .A2(\regfile/reg_out[25][25] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][25] ), .ZN(n5898) );
  AOI22_X1 U4820 ( .A1(n5767), .A2(\regfile/reg_out[29][25] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][25] ), .ZN(n5899) );
  AOI22_X1 U4821 ( .A1(n5774), .A2(\regfile/reg_out[5][25] ), .B1(n5775), .B2(
        \regfile/reg_out[4][25] ), .ZN(n5900) );
  OAI21_X1 U4822 ( .B1(n5884), .B2(n5903), .A(n5893), .ZN(n5902) );
  INV_X1 U4823 ( .A(n5904), .ZN(n5901) );
  AOI22_X1 U4824 ( .A1(n5752), .A2(\regfile/reg_out[19][24] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][24] ), .ZN(n5906) );
  AOI22_X1 U4825 ( .A1(n5757), .A2(\regfile/reg_out[21][24] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][24] ), .ZN(n5907) );
  AOI22_X1 U4826 ( .A1(n5762), .A2(\regfile/reg_out[25][24] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][24] ), .ZN(n5908) );
  AOI22_X1 U4827 ( .A1(n5767), .A2(\regfile/reg_out[29][24] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][24] ), .ZN(n5909) );
  AOI22_X1 U4828 ( .A1(n5774), .A2(\regfile/reg_out[5][24] ), .B1(n5775), .B2(
        \regfile/reg_out[4][24] ), .ZN(n5910) );
  OAI21_X1 U4829 ( .B1(n5913), .B2(n5884), .A(n5893), .ZN(n5912) );
  INV_X1 U4830 ( .A(n5914), .ZN(n5911) );
  AOI22_X1 U4831 ( .A1(n5752), .A2(\regfile/reg_out[19][23] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][23] ), .ZN(n5915) );
  AOI22_X1 U4832 ( .A1(n5757), .A2(\regfile/reg_out[21][23] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][23] ), .ZN(n5916) );
  AOI22_X1 U4833 ( .A1(n5762), .A2(\regfile/reg_out[25][23] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][23] ), .ZN(n5917) );
  AOI22_X1 U4834 ( .A1(n5767), .A2(\regfile/reg_out[29][23] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][23] ), .ZN(n5918) );
  AOI22_X1 U4835 ( .A1(n5774), .A2(\regfile/reg_out[5][23] ), .B1(n5775), .B2(
        \regfile/reg_out[4][23] ), .ZN(n5919) );
  AOI22_X1 U4836 ( .A1(n5752), .A2(\regfile/reg_out[19][22] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][22] ), .ZN(n5920) );
  AOI22_X1 U4837 ( .A1(n5757), .A2(\regfile/reg_out[21][22] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][22] ), .ZN(n5921) );
  AOI22_X1 U4838 ( .A1(n5762), .A2(\regfile/reg_out[25][22] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][22] ), .ZN(n5922) );
  AOI22_X1 U4839 ( .A1(n5767), .A2(\regfile/reg_out[29][22] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][22] ), .ZN(n5923) );
  AOI22_X1 U4840 ( .A1(n5774), .A2(\regfile/reg_out[5][22] ), .B1(n5775), .B2(
        \regfile/reg_out[4][22] ), .ZN(n5924) );
  AOI22_X1 U4841 ( .A1(n5752), .A2(\regfile/reg_out[19][21] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][21] ), .ZN(n5925) );
  AOI22_X1 U4842 ( .A1(n5757), .A2(\regfile/reg_out[21][21] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][21] ), .ZN(n5926) );
  AOI22_X1 U4843 ( .A1(n5762), .A2(\regfile/reg_out[25][21] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][21] ), .ZN(n5927) );
  AOI22_X1 U4844 ( .A1(n5767), .A2(\regfile/reg_out[29][21] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][21] ), .ZN(n5928) );
  AOI22_X1 U4845 ( .A1(n5774), .A2(\regfile/reg_out[5][21] ), .B1(n5775), .B2(
        \regfile/reg_out[4][21] ), .ZN(n5929) );
  AOI22_X1 U4846 ( .A1(n5752), .A2(\regfile/reg_out[19][20] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][20] ), .ZN(n5930) );
  AOI22_X1 U4847 ( .A1(n5757), .A2(\regfile/reg_out[21][20] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][20] ), .ZN(n5931) );
  AOI22_X1 U4848 ( .A1(n5762), .A2(\regfile/reg_out[25][20] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][20] ), .ZN(n5932) );
  AOI22_X1 U4849 ( .A1(n5767), .A2(\regfile/reg_out[29][20] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][20] ), .ZN(n5933) );
  AOI22_X1 U4850 ( .A1(n5774), .A2(\regfile/reg_out[5][20] ), .B1(n5775), .B2(
        \regfile/reg_out[4][20] ), .ZN(n5934) );
  OAI22_X1 U4851 ( .A1(n5936), .A2(n5790), .B1(n5895), .B2(n5792), .ZN(n5935)
         );
  OAI22_X1 U4852 ( .A1(n5938), .A2(n5939), .B1(n5802), .B2(n5940), .ZN(n5937)
         );
  AOI22_X1 U4853 ( .A1(n5752), .A2(\regfile/reg_out[19][1] ), .B1(n5753), .B2(
        \regfile/reg_out[18][1] ), .ZN(n5941) );
  AOI22_X1 U4854 ( .A1(n5757), .A2(\regfile/reg_out[21][1] ), .B1(n5758), .B2(
        \regfile/reg_out[20][1] ), .ZN(n5942) );
  AOI22_X1 U4855 ( .A1(n5762), .A2(\regfile/reg_out[25][1] ), .B1(n5763), .B2(
        \regfile/reg_out[24][1] ), .ZN(n5943) );
  AOI22_X1 U4856 ( .A1(n5767), .A2(\regfile/reg_out[29][1] ), .B1(n5768), .B2(
        \regfile/reg_out[28][1] ), .ZN(n5944) );
  AOI22_X1 U4857 ( .A1(n5774), .A2(\regfile/reg_out[5][1] ), .B1(n5775), .B2(
        \regfile/reg_out[4][1] ), .ZN(n5945) );
  AOI22_X1 U4858 ( .A1(n5752), .A2(\regfile/reg_out[19][19] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][19] ), .ZN(n5946) );
  AOI22_X1 U4859 ( .A1(n5757), .A2(\regfile/reg_out[21][19] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][19] ), .ZN(n5947) );
  AOI22_X1 U4860 ( .A1(n5762), .A2(\regfile/reg_out[25][19] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][19] ), .ZN(n5948) );
  AOI22_X1 U4861 ( .A1(n5767), .A2(\regfile/reg_out[29][19] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][19] ), .ZN(n5949) );
  AOI22_X1 U4862 ( .A1(n5774), .A2(\regfile/reg_out[5][19] ), .B1(n5775), .B2(
        \regfile/reg_out[4][19] ), .ZN(n5950) );
  AOI22_X1 U4863 ( .A1(n5752), .A2(\regfile/reg_out[19][18] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][18] ), .ZN(n5951) );
  AOI22_X1 U4864 ( .A1(n5757), .A2(\regfile/reg_out[21][18] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][18] ), .ZN(n5952) );
  AOI22_X1 U4865 ( .A1(n5762), .A2(\regfile/reg_out[25][18] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][18] ), .ZN(n5953) );
  AOI22_X1 U4866 ( .A1(n5767), .A2(\regfile/reg_out[29][18] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][18] ), .ZN(n5954) );
  AOI22_X1 U4867 ( .A1(n5774), .A2(\regfile/reg_out[5][18] ), .B1(n5775), .B2(
        \regfile/reg_out[4][18] ), .ZN(n5955) );
  AOI22_X1 U4868 ( .A1(n5752), .A2(\regfile/reg_out[19][17] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][17] ), .ZN(n5956) );
  AOI22_X1 U4869 ( .A1(n5757), .A2(\regfile/reg_out[21][17] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][17] ), .ZN(n5957) );
  AOI22_X1 U4870 ( .A1(n5762), .A2(\regfile/reg_out[25][17] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][17] ), .ZN(n5958) );
  AOI22_X1 U4871 ( .A1(n5767), .A2(\regfile/reg_out[29][17] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][17] ), .ZN(n5959) );
  AOI22_X1 U4872 ( .A1(n5774), .A2(\regfile/reg_out[5][17] ), .B1(n5775), .B2(
        \regfile/reg_out[4][17] ), .ZN(n5960) );
  NOR3_X1 U4873 ( .A1(n5963), .A2(n5964), .A3(n5965), .ZN(n5962) );
  AOI22_X1 U4874 ( .A1(n6546), .A2(n5966), .B1(\Mpath/the_memhandle/N239 ), 
        .B2(n6541), .ZN(n5964) );
  INV_X1 U4875 ( .A(\Mpath/the_memhandle/N86 ), .ZN(n5963) );
  AOI22_X1 U4876 ( .A1(n5752), .A2(\regfile/reg_out[19][16] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][16] ), .ZN(n5969) );
  AOI22_X1 U4877 ( .A1(n5757), .A2(\regfile/reg_out[21][16] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][16] ), .ZN(n5970) );
  AOI22_X1 U4878 ( .A1(n5762), .A2(\regfile/reg_out[25][16] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][16] ), .ZN(n5971) );
  AOI22_X1 U4879 ( .A1(n5767), .A2(\regfile/reg_out[29][16] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][16] ), .ZN(n5972) );
  AOI22_X1 U4880 ( .A1(n5774), .A2(\regfile/reg_out[5][16] ), .B1(n5775), .B2(
        \regfile/reg_out[4][16] ), .ZN(n5973) );
  AOI22_X1 U4881 ( .A1(n5752), .A2(\regfile/reg_out[19][15] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][15] ), .ZN(n5974) );
  AOI22_X1 U4882 ( .A1(n5757), .A2(\regfile/reg_out[21][15] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][15] ), .ZN(n5975) );
  AOI22_X1 U4883 ( .A1(n5762), .A2(\regfile/reg_out[25][15] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][15] ), .ZN(n5976) );
  AOI22_X1 U4884 ( .A1(n5767), .A2(\regfile/reg_out[29][15] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][15] ), .ZN(n5977) );
  AOI22_X1 U4885 ( .A1(n5774), .A2(\regfile/reg_out[5][15] ), .B1(n5775), .B2(
        \regfile/reg_out[4][15] ), .ZN(n5978) );
  AOI22_X1 U4886 ( .A1(n5752), .A2(\regfile/reg_out[19][14] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][14] ), .ZN(n5979) );
  AOI22_X1 U4887 ( .A1(n5757), .A2(\regfile/reg_out[21][14] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][14] ), .ZN(n5980) );
  AOI22_X1 U4888 ( .A1(n5762), .A2(\regfile/reg_out[25][14] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][14] ), .ZN(n5981) );
  AOI22_X1 U4889 ( .A1(n5767), .A2(\regfile/reg_out[29][14] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][14] ), .ZN(n5982) );
  AOI22_X1 U4890 ( .A1(n5774), .A2(\regfile/reg_out[5][14] ), .B1(n5775), .B2(
        \regfile/reg_out[4][14] ), .ZN(n5983) );
  AOI22_X1 U4891 ( .A1(n5752), .A2(\regfile/reg_out[19][13] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][13] ), .ZN(n5984) );
  AOI22_X1 U4892 ( .A1(n5757), .A2(\regfile/reg_out[21][13] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][13] ), .ZN(n5985) );
  AOI22_X1 U4893 ( .A1(n5762), .A2(\regfile/reg_out[25][13] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][13] ), .ZN(n5986) );
  AOI22_X1 U4894 ( .A1(n5767), .A2(\regfile/reg_out[29][13] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][13] ), .ZN(n5987) );
  AOI22_X1 U4895 ( .A1(n5774), .A2(\regfile/reg_out[5][13] ), .B1(n5775), .B2(
        \regfile/reg_out[4][13] ), .ZN(n5988) );
  AOI22_X1 U4896 ( .A1(n5752), .A2(\regfile/reg_out[19][12] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][12] ), .ZN(n5989) );
  AOI22_X1 U4897 ( .A1(n5757), .A2(\regfile/reg_out[21][12] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][12] ), .ZN(n5990) );
  AOI22_X1 U4898 ( .A1(n5762), .A2(\regfile/reg_out[25][12] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][12] ), .ZN(n5991) );
  AOI22_X1 U4899 ( .A1(n5767), .A2(\regfile/reg_out[29][12] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][12] ), .ZN(n5992) );
  AOI22_X1 U4900 ( .A1(n5774), .A2(\regfile/reg_out[5][12] ), .B1(n5775), .B2(
        \regfile/reg_out[4][12] ), .ZN(n5993) );
  AOI22_X1 U4901 ( .A1(n5752), .A2(\regfile/reg_out[19][11] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][11] ), .ZN(n5994) );
  AOI22_X1 U4902 ( .A1(n5757), .A2(\regfile/reg_out[21][11] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][11] ), .ZN(n5995) );
  AOI22_X1 U4903 ( .A1(n5762), .A2(\regfile/reg_out[25][11] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][11] ), .ZN(n5996) );
  AOI22_X1 U4904 ( .A1(n5767), .A2(\regfile/reg_out[29][11] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][11] ), .ZN(n5997) );
  AOI22_X1 U4905 ( .A1(n5774), .A2(\regfile/reg_out[5][11] ), .B1(n5775), .B2(
        \regfile/reg_out[4][11] ), .ZN(n5998) );
  INV_X1 U4906 ( .A(n5785), .ZN(n5748) );
  OAI221_X1 U4907 ( .B1(n5791), .B2(n6000), .C1(n6001), .C2(n5938), .A(n6002), 
        .ZN(n5999) );
  AOI22_X1 U4908 ( .A1(\Mpath/the_memhandle/N38 ), .A2(n6546), .B1(
        \Mpath/the_memhandle/N37 ), .B2(n6544), .ZN(n6002) );
  INV_X1 U4909 ( .A(\Mpath/the_memhandle/N36 ), .ZN(n6000) );
  NOR2_X1 U4910 ( .A1(n5965), .A2(n6003), .ZN(n5747) );
  NOR2_X1 U4911 ( .A1(n6004), .A2(n5965), .ZN(n5746) );
  INV_X1 U4912 ( .A(n5967), .ZN(n5965) );
  NOR2_X1 U4913 ( .A1(\Mpath/the_memhandle/N34 ), .A2(
        \Mpath/the_memhandle/N72 ), .ZN(n5967) );
  AOI22_X1 U4914 ( .A1(n5752), .A2(\regfile/reg_out[19][10] ), .B1(n5753), 
        .B2(\regfile/reg_out[18][10] ), .ZN(n6005) );
  AOI22_X1 U4915 ( .A1(n5757), .A2(\regfile/reg_out[21][10] ), .B1(n5758), 
        .B2(\regfile/reg_out[20][10] ), .ZN(n6006) );
  AOI22_X1 U4916 ( .A1(n5762), .A2(\regfile/reg_out[25][10] ), .B1(n5763), 
        .B2(\regfile/reg_out[24][10] ), .ZN(n6007) );
  AOI22_X1 U4917 ( .A1(n5767), .A2(\regfile/reg_out[29][10] ), .B1(n5768), 
        .B2(\regfile/reg_out[28][10] ), .ZN(n6008) );
  AOI22_X1 U4918 ( .A1(n5774), .A2(\regfile/reg_out[5][10] ), .B1(n5775), .B2(
        \regfile/reg_out[4][10] ), .ZN(n6009) );
  OAI22_X1 U4919 ( .A1(n6011), .A2(n5790), .B1(n5905), .B2(n5792), .ZN(n6010)
         );
  NAND2_X1 U4920 ( .A1(\Mpath/the_memhandle/N74 ), .A2(
        \Mpath/the_memhandle/N72 ), .ZN(n5792) );
  NAND2_X1 U4921 ( .A1(\Mpath/the_memhandle/N76 ), .A2(
        \Mpath/the_memhandle/N72 ), .ZN(n5790) );
  OAI22_X1 U4922 ( .A1(n6012), .A2(\Mpath/the_memhandle/N243 ), .B1(
        \Mpath/the_memhandle/N72 ), .B2(n6004), .ZN(n5787) );
  INV_X1 U4923 ( .A(n6003), .ZN(n6004) );
  INV_X1 U4924 ( .A(\Mpath/the_memhandle/N72 ), .ZN(n6012) );
  OAI21_X1 U4925 ( .B1(\Mpath/the_memhandle/N72 ), .B2(n6003), .A(n6013), .ZN(
        n5786) );
  NAND2_X1 U4926 ( .A1(\Mpath/the_memhandle/N77 ), .A2(
        \Mpath/the_memhandle/N72 ), .ZN(n6013) );
  NOR2_X1 U4927 ( .A1(n5966), .A2(n5968), .ZN(n6003) );
  NOR2_X1 U4928 ( .A1(\Mpath/the_memhandle/N120 ), .A2(
        \Mpath/the_memhandle/N86 ), .ZN(n5968) );
  INV_X1 U4929 ( .A(\Mpath/the_memhandle/N239 ), .ZN(n5966) );
  OAI22_X1 U4930 ( .A1(n5802), .A2(n5961), .B1(n5938), .B2(n6015), .ZN(n6014)
         );
  INV_X1 U4931 ( .A(D_DATA_INBUS[0]), .ZN(n6015) );
  INV_X1 U4932 ( .A(\Mpath/the_memhandle/N39 ), .ZN(n5938) );
  INV_X1 U4933 ( .A(\Mpath/the_memhandle/N37 ), .ZN(n5802) );
  AOI22_X1 U4934 ( .A1(n5752), .A2(\regfile/reg_out[19][0] ), .B1(n5753), .B2(
        \regfile/reg_out[18][0] ), .ZN(n6016) );
  NAND3_X1 U4937 ( .A1(n6019), .A2(n6020), .A3(n6017), .ZN(n5750) );
  AOI22_X1 U4940 ( .A1(n5757), .A2(\regfile/reg_out[21][0] ), .B1(n5758), .B2(
        \regfile/reg_out[20][0] ), .ZN(n6023) );
  AOI22_X1 U4946 ( .A1(n5762), .A2(\regfile/reg_out[25][0] ), .B1(n5763), .B2(
        \regfile/reg_out[24][0] ), .ZN(n6027) );
  AOI22_X1 U4951 ( .A1(n5767), .A2(\regfile/reg_out[29][0] ), .B1(n5768), .B2(
        \regfile/reg_out[28][0] ), .ZN(n6031) );
  NAND3_X1 U4954 ( .A1(n6032), .A2(rs2_addr[4]), .A3(n6018), .ZN(n5765) );
  NAND3_X1 U4955 ( .A1(n6029), .A2(n6032), .A3(rs2_addr[1]), .ZN(n5764) );
  NAND3_X1 U4957 ( .A1(rs2_addr[1]), .A2(n6022), .A3(n6033), .ZN(n5770) );
  NAND3_X1 U4958 ( .A1(n6022), .A2(n6034), .A3(n6035), .ZN(n5769) );
  AOI22_X1 U4959 ( .A1(n5774), .A2(\regfile/reg_out[5][0] ), .B1(n5775), .B2(
        \regfile/reg_out[4][0] ), .ZN(n6036) );
  NAND3_X1 U4963 ( .A1(rs2_addr[1]), .A2(rs2_addr[2]), .A3(n6033), .ZN(n5771)
         );
  NAND2_X1 U4966 ( .A1(n6035), .A2(n6032), .ZN(n5776) );
  INV_X1 U4987 ( .A(\Mcontrol/st_logic/N2 ), .ZN(
        \Mcontrol/st_logic/load_stall ) );
  INV_X1 U4988 ( .A(\Mcontrol/st_logic/N8 ), .ZN(
        \Mcontrol/st_logic/branchmul_stall ) );
  INV_X1 U4989 ( .A(\Mcontrol/st_logic/N6 ), .ZN(
        \Mcontrol/st_logic/branchlw_stall ) );
  INV_X1 U4990 ( .A(\Mcontrol/st_logic/N4 ), .ZN(
        \Mcontrol/st_logic/branch_uses_regb ) );
  INV_X1 U4991 ( .A(\Mcontrol/st_logic/N3 ), .ZN(
        \Mcontrol/st_logic/branch_uses_rega ) );
  INV_X1 U4992 ( .A(\Mcontrol/st_logic/N5 ), .ZN(
        \Mcontrol/st_logic/branch_uses_main_mem_result ) );
  INV_X1 U4993 ( .A(\Mcontrol/st_logic/N7 ), .ZN(
        \Mcontrol/st_logic/branch_uses_main_exe_result ) );
  OAI21_X1 U4994 ( .B1(\Mcontrol/st_logic/N10 ), .B2(n7109), .A(n5504), .ZN(
        \Mcontrol/stall_decode ) );
  AOI21_X1 U4995 ( .B1(n7218), .B2(\Mcontrol/Operation_decoding32/N1952 ), .A(
        \Mcontrol/Operation_decoding32/N1964 ), .ZN(n6053) );
  NAND4_X1 U4996 ( .A1(\Mcontrol/Operation_decoding32/N1907 ), .A2(n6058), 
        .A3(\Mcontrol/Operation_decoding32/N89 ), .A4(net56977), .ZN(n6055) );
  NOR3_X1 U4997 ( .A1(\Mcontrol/Operation_decoding32/N1958 ), .A2(
        \Mcontrol/Operation_decoding32/N1970 ), .A3(n6054), .ZN(n6058) );
  AOI21_X1 U4998 ( .B1(\Mcontrol/Operation_decoding32/N62 ), .B2(
        \Mcontrol/Operation_decoding32/N89 ), .A(n7416), .ZN(n6069) );
  INV_X1 U5005 ( .A(n7227), .ZN(n6076) );
  OAI211_X1 U5006 ( .C1(n6077), .C2(n6054), .A(n7598), .B(n6065), .ZN(n6078)
         );
  INV_X1 U5007 ( .A(n5519), .ZN(\Mcontrol/d_instr [1]) );
  AOI22_X1 U5008 ( .A1(n7603), .A2(\regfile/reg_out[19][1] ), .B1(n7621), .B2(
        \regfile/reg_out[18][1] ), .ZN(n6081) );
  AOI22_X1 U5009 ( .A1(n7502), .A2(\regfile/reg_out[21][1] ), .B1(n7514), .B2(
        \regfile/reg_out[20][1] ), .ZN(n6082) );
  AOI22_X1 U5010 ( .A1(n5637), .A2(\regfile/reg_out[25][1] ), .B1(n5638), .B2(
        \regfile/reg_out[24][1] ), .ZN(n6083) );
  AOI22_X1 U5011 ( .A1(n5642), .A2(\regfile/reg_out[29][1] ), .B1(n5643), .B2(
        \regfile/reg_out[28][1] ), .ZN(n6084) );
  AOI22_X1 U5012 ( .A1(n5649), .A2(\regfile/reg_out[5][1] ), .B1(n5650), .B2(
        \regfile/reg_out[4][1] ), .ZN(n6085) );
  INV_X1 U5013 ( .A(n6086), .ZN(n5585) );
  AOI22_X1 U5015 ( .A1(n6091), .A2(n6968), .B1(\Mpath/N190 ), .B2(n6092), .ZN(
        n6090) );
  OAI22_X1 U5016 ( .A1(net56668), .A2(n6093), .B1(n6095), .B2(n7442), .ZN(
        n6080) );
  NAND2_X1 U5017 ( .A1(n6097), .A2(n6096), .ZN(n6095) );
  AOI22_X1 U5028 ( .A1(n7603), .A2(\regfile/reg_out[19][9] ), .B1(n7592), .B2(
        \regfile/reg_out[18][9] ), .ZN(n6108) );
  AOI22_X1 U5029 ( .A1(n7503), .A2(\regfile/reg_out[21][9] ), .B1(n5633), .B2(
        \regfile/reg_out[20][9] ), .ZN(n6109) );
  AOI22_X1 U5030 ( .A1(n5637), .A2(\regfile/reg_out[25][9] ), .B1(n5638), .B2(
        \regfile/reg_out[24][9] ), .ZN(n6110) );
  AOI22_X1 U5031 ( .A1(n5642), .A2(\regfile/reg_out[29][9] ), .B1(n5643), .B2(
        \regfile/reg_out[28][9] ), .ZN(n6111) );
  AOI22_X1 U5032 ( .A1(n5649), .A2(\regfile/reg_out[5][9] ), .B1(n5650), .B2(
        \regfile/reg_out[4][9] ), .ZN(n6112) );
  INV_X1 U5033 ( .A(n6113), .ZN(n5522) );
  AOI22_X1 U5035 ( .A1(n6091), .A2(n6117), .B1(\Mpath/N190 ), .B2(n6118), .ZN(
        n6116) );
  OAI222_X1 U5036 ( .A1(n7255), .A2(n6047), .B1(n7176), .B2(n6120), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n5914), .ZN(n6119) );
  AOI22_X1 U5037 ( .A1(n7603), .A2(\regfile/reg_out[19][8] ), .B1(n7592), .B2(
        \regfile/reg_out[18][8] ), .ZN(n6121) );
  AOI22_X1 U5038 ( .A1(n7502), .A2(\regfile/reg_out[21][8] ), .B1(n7612), .B2(
        \regfile/reg_out[20][8] ), .ZN(n6122) );
  AOI22_X1 U5039 ( .A1(n5637), .A2(\regfile/reg_out[25][8] ), .B1(n5638), .B2(
        \regfile/reg_out[24][8] ), .ZN(n6123) );
  AOI22_X1 U5040 ( .A1(n5642), .A2(\regfile/reg_out[29][8] ), .B1(n5643), .B2(
        \regfile/reg_out[28][8] ), .ZN(n6124) );
  AOI22_X1 U5041 ( .A1(n5649), .A2(\regfile/reg_out[5][8] ), .B1(n5650), .B2(
        \regfile/reg_out[4][8] ), .ZN(n6125) );
  INV_X1 U5042 ( .A(n6126), .ZN(n5528) );
  AOI22_X1 U5044 ( .A1(n6091), .A2(n6130), .B1(\Mpath/N190 ), .B2(n6131), .ZN(
        n6129) );
  AOI22_X1 U5046 ( .A1(n7603), .A2(\regfile/reg_out[19][7] ), .B1(n7461), .B2(
        \regfile/reg_out[18][7] ), .ZN(n6133) );
  AOI22_X1 U5047 ( .A1(n7502), .A2(\regfile/reg_out[21][7] ), .B1(n7514), .B2(
        \regfile/reg_out[20][7] ), .ZN(n6134) );
  AOI22_X1 U5048 ( .A1(n5637), .A2(\regfile/reg_out[25][7] ), .B1(n5638), .B2(
        \regfile/reg_out[24][7] ), .ZN(n6135) );
  AOI22_X1 U5049 ( .A1(n5642), .A2(\regfile/reg_out[29][7] ), .B1(n5643), .B2(
        \regfile/reg_out[28][7] ), .ZN(n6136) );
  AOI22_X1 U5050 ( .A1(n5649), .A2(\regfile/reg_out[5][7] ), .B1(n5650), .B2(
        \regfile/reg_out[4][7] ), .ZN(n6137) );
  INV_X1 U5051 ( .A(n6138), .ZN(n5531) );
  AOI22_X1 U5053 ( .A1(n6091), .A2(n6142), .B1(\Mpath/N190 ), .B2(n6143), .ZN(
        n6141) );
  AOI22_X1 U5055 ( .A1(n7603), .A2(\regfile/reg_out[19][6] ), .B1(n7592), .B2(
        \regfile/reg_out[18][6] ), .ZN(n6145) );
  AOI22_X1 U5056 ( .A1(n7502), .A2(\regfile/reg_out[21][6] ), .B1(n5633), .B2(
        \regfile/reg_out[20][6] ), .ZN(n6146) );
  AOI22_X1 U5057 ( .A1(n5637), .A2(\regfile/reg_out[25][6] ), .B1(n5638), .B2(
        \regfile/reg_out[24][6] ), .ZN(n6147) );
  AOI22_X1 U5058 ( .A1(n5642), .A2(\regfile/reg_out[29][6] ), .B1(n5643), .B2(
        \regfile/reg_out[28][6] ), .ZN(n6148) );
  AOI22_X1 U5059 ( .A1(n5649), .A2(\regfile/reg_out[5][6] ), .B1(n5650), .B2(
        \regfile/reg_out[4][6] ), .ZN(n6149) );
  INV_X1 U5060 ( .A(n6150), .ZN(n5534) );
  AOI22_X1 U5062 ( .A1(n6091), .A2(n6154), .B1(\Mpath/N190 ), .B2(n6155), .ZN(
        n6153) );
  AOI22_X1 U5064 ( .A1(n7603), .A2(\regfile/reg_out[19][5] ), .B1(n5628), .B2(
        \regfile/reg_out[18][5] ), .ZN(n6157) );
  AOI22_X1 U5065 ( .A1(n7502), .A2(\regfile/reg_out[21][5] ), .B1(n7514), .B2(
        \regfile/reg_out[20][5] ), .ZN(n6158) );
  AOI22_X1 U5066 ( .A1(n5637), .A2(\regfile/reg_out[25][5] ), .B1(n5638), .B2(
        \regfile/reg_out[24][5] ), .ZN(n6159) );
  AOI22_X1 U5067 ( .A1(n5642), .A2(\regfile/reg_out[29][5] ), .B1(n5643), .B2(
        \regfile/reg_out[28][5] ), .ZN(n6160) );
  AOI22_X1 U5068 ( .A1(n5649), .A2(\regfile/reg_out[5][5] ), .B1(n5650), .B2(
        \regfile/reg_out[4][5] ), .ZN(n6161) );
  INV_X1 U5069 ( .A(n6162), .ZN(n5537) );
  AOI22_X1 U5071 ( .A1(n6091), .A2(n6166), .B1(\Mpath/N190 ), .B2(n6167), .ZN(
        n6165) );
  OAI22_X1 U5072 ( .A1(n6093), .A2(n5894), .B1(n6170), .B2(n6171), .ZN(n6169)
         );
  AOI22_X1 U5073 ( .A1(n6103), .A2(n6172), .B1(n7351), .B2(n7450), .ZN(n6170)
         );
  OAI222_X1 U5074 ( .A1(n7250), .A2(n5894), .B1(n7279), .B2(n5518), .C1(n5516), 
        .C2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n6172) );
  AOI22_X1 U5075 ( .A1(n7603), .A2(\regfile/reg_out[19][4] ), .B1(n7592), .B2(
        \regfile/reg_out[18][4] ), .ZN(n6174) );
  AOI22_X1 U5076 ( .A1(n7503), .A2(\regfile/reg_out[21][4] ), .B1(n5633), .B2(
        \regfile/reg_out[20][4] ), .ZN(n6175) );
  AOI22_X1 U5077 ( .A1(n5637), .A2(\regfile/reg_out[25][4] ), .B1(n7096), .B2(
        \regfile/reg_out[24][4] ), .ZN(n6176) );
  AOI22_X1 U5078 ( .A1(n5642), .A2(\regfile/reg_out[29][4] ), .B1(n5643), .B2(
        \regfile/reg_out[28][4] ), .ZN(n6177) );
  AOI22_X1 U5079 ( .A1(n5649), .A2(\regfile/reg_out[5][4] ), .B1(n5650), .B2(
        \regfile/reg_out[4][4] ), .ZN(n6178) );
  INV_X1 U5080 ( .A(n6179), .ZN(n5540) );
  AOI22_X1 U5082 ( .A1(n6091), .A2(n6183), .B1(\Mpath/N190 ), .B2(n6184), .ZN(
        n6182) );
  OAI22_X1 U5083 ( .A1(n6093), .A2(n5904), .B1(n6186), .B2(n6171), .ZN(n6185)
         );
  AOI22_X1 U5084 ( .A1(n6103), .A2(n6187), .B1(\Mcontrol/d_instr [3]), .B2(
        n6173), .ZN(n6186) );
  INV_X1 U5085 ( .A(n5517), .ZN(\Mcontrol/d_instr [3]) );
  OAI222_X1 U5086 ( .A1(n7250), .A2(n5904), .B1(n5519), .B2(n7279), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n5517), .ZN(n6187) );
  AOI22_X1 U5087 ( .A1(n7603), .A2(\regfile/reg_out[19][3] ), .B1(n5628), .B2(
        \regfile/reg_out[18][3] ), .ZN(n6188) );
  AOI22_X1 U5088 ( .A1(n7503), .A2(\regfile/reg_out[21][3] ), .B1(n5633), .B2(
        \regfile/reg_out[20][3] ), .ZN(n6189) );
  AOI22_X1 U5089 ( .A1(n5637), .A2(\regfile/reg_out[25][3] ), .B1(n7096), .B2(
        \regfile/reg_out[24][3] ), .ZN(n6190) );
  AOI22_X1 U5090 ( .A1(n5642), .A2(\regfile/reg_out[29][3] ), .B1(n5643), .B2(
        \regfile/reg_out[28][3] ), .ZN(n6191) );
  AOI22_X1 U5091 ( .A1(n5649), .A2(\regfile/reg_out[5][3] ), .B1(n5650), .B2(
        \regfile/reg_out[4][3] ), .ZN(n6192) );
  INV_X1 U5092 ( .A(n6193), .ZN(n5543) );
  AOI22_X1 U5094 ( .A1(n6091), .A2(n6197), .B1(\Mpath/N190 ), .B2(n6198), .ZN(
        n6196) );
  NOR2_X1 U5097 ( .A1(n7037), .A2(n6063), .ZN(n6101) );
  INV_X1 U5099 ( .A(n5518), .ZN(\Mcontrol/d_instr [2]) );
  OAI222_X1 U5100 ( .A1(n6094), .A2(n5914), .B1(n7262), .B2(n5520), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n5518), .ZN(n6201) );
  NOR2_X1 U5103 ( .A1(n7587), .A2(net57236), .ZN(n6168) );
  AOI22_X1 U5104 ( .A1(n7603), .A2(\regfile/reg_out[19][2] ), .B1(n7621), .B2(
        \regfile/reg_out[18][2] ), .ZN(n6203) );
  AOI22_X1 U5105 ( .A1(n7502), .A2(\regfile/reg_out[21][2] ), .B1(n5633), .B2(
        \regfile/reg_out[20][2] ), .ZN(n6204) );
  AOI22_X1 U5106 ( .A1(n5637), .A2(\regfile/reg_out[25][2] ), .B1(n5638), .B2(
        \regfile/reg_out[24][2] ), .ZN(n6205) );
  AOI22_X1 U5107 ( .A1(n5642), .A2(\regfile/reg_out[29][2] ), .B1(n5643), .B2(
        \regfile/reg_out[28][2] ), .ZN(n6206) );
  AOI22_X1 U5108 ( .A1(n5649), .A2(\regfile/reg_out[5][2] ), .B1(n5650), .B2(
        \regfile/reg_out[4][2] ), .ZN(n6207) );
  INV_X1 U5109 ( .A(n6208), .ZN(n5552) );
  AOI22_X1 U5111 ( .A1(n6091), .A2(n6212), .B1(\Mpath/N190 ), .B2(n6213), .ZN(
        n6211) );
  OAI21_X1 U5112 ( .B1(n6052), .B2(n5884), .A(n5893), .ZN(n6214) );
  AOI22_X1 U5114 ( .A1(n7603), .A2(\regfile/reg_out[19][23] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][23] ), .ZN(n6215) );
  AOI22_X1 U5115 ( .A1(n7503), .A2(\regfile/reg_out[21][23] ), .B1(n7611), 
        .B2(\regfile/reg_out[20][23] ), .ZN(n6216) );
  AOI22_X1 U5116 ( .A1(n5637), .A2(\regfile/reg_out[25][23] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][23] ), .ZN(n6217) );
  AOI22_X1 U5117 ( .A1(n5642), .A2(\regfile/reg_out[29][23] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][23] ), .ZN(n6218) );
  AOI22_X1 U5118 ( .A1(n5649), .A2(\regfile/reg_out[5][23] ), .B1(n5650), .B2(
        \regfile/reg_out[4][23] ), .ZN(n6219) );
  INV_X1 U5119 ( .A(n6220), .ZN(n5573) );
  AOI22_X1 U5121 ( .A1(n6091), .A2(n6225), .B1(\Mpath/N190 ), .B2(n6226), .ZN(
        n6224) );
  OAI21_X1 U5122 ( .B1(n6044), .B2(n5884), .A(n5893), .ZN(n6227) );
  AOI22_X1 U5124 ( .A1(n7603), .A2(\regfile/reg_out[19][22] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][22] ), .ZN(n6228) );
  AOI22_X1 U5126 ( .A1(n5637), .A2(\regfile/reg_out[25][22] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][22] ), .ZN(n6230) );
  AOI22_X1 U5127 ( .A1(n5642), .A2(\regfile/reg_out[29][22] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][22] ), .ZN(n6231) );
  AOI22_X1 U5128 ( .A1(n5649), .A2(\regfile/reg_out[5][22] ), .B1(n5650), .B2(
        \regfile/reg_out[4][22] ), .ZN(n6232) );
  INV_X1 U5129 ( .A(n6233), .ZN(n5576) );
  AOI22_X1 U5131 ( .A1(n6091), .A2(n6237), .B1(\Mpath/N190 ), .B2(n6238), .ZN(
        n6236) );
  OAI21_X1 U5132 ( .B1(n6046), .B2(n5884), .A(n5893), .ZN(n6239) );
  AOI22_X1 U5134 ( .A1(n7603), .A2(\regfile/reg_out[19][21] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][21] ), .ZN(n6240) );
  AOI22_X1 U5135 ( .A1(n7502), .A2(\regfile/reg_out[21][21] ), .B1(n7514), 
        .B2(\regfile/reg_out[20][21] ), .ZN(n6241) );
  AOI22_X1 U5136 ( .A1(n5637), .A2(\regfile/reg_out[25][21] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][21] ), .ZN(n6242) );
  AOI22_X1 U5137 ( .A1(n5642), .A2(\regfile/reg_out[29][21] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][21] ), .ZN(n6243) );
  AOI22_X1 U5138 ( .A1(n5649), .A2(\regfile/reg_out[5][21] ), .B1(n5650), .B2(
        \regfile/reg_out[4][21] ), .ZN(n6244) );
  INV_X1 U5139 ( .A(n6245), .ZN(n5579) );
  AOI22_X1 U5141 ( .A1(n6091), .A2(n6249), .B1(\Mpath/N190 ), .B2(n6250), .ZN(
        n6248) );
  NAND3_X1 U5142 ( .A1(n7506), .A2(n7436), .A3(n6045), .ZN(n5880) );
  OAI21_X1 U5143 ( .B1(n5884), .B2(n6039), .A(n5893), .ZN(n6251) );
  INV_X1 U5144 ( .A(n5882), .ZN(n5893) );
  OAI21_X1 U5145 ( .B1(n5846), .B2(n7510), .A(n6254), .ZN(n5882) );
  OR2_X1 U5146 ( .A1(n6255), .A2(\Mcontrol/Operation_decoding32/N1982 ), .ZN(
        n5884) );
  NOR2_X1 U5147 ( .A1(n7506), .A2(n7159), .ZN(n5847) );
  AOI22_X1 U5149 ( .A1(n7603), .A2(\regfile/reg_out[19][20] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][20] ), .ZN(n6256) );
  AOI22_X1 U5150 ( .A1(n7503), .A2(\regfile/reg_out[21][20] ), .B1(n5633), 
        .B2(\regfile/reg_out[20][20] ), .ZN(n6257) );
  AOI22_X1 U5151 ( .A1(n5637), .A2(\regfile/reg_out[25][20] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][20] ), .ZN(n6258) );
  AOI22_X1 U5152 ( .A1(n5642), .A2(\regfile/reg_out[29][20] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][20] ), .ZN(n6259) );
  AOI22_X1 U5153 ( .A1(n5649), .A2(\regfile/reg_out[5][20] ), .B1(n5650), .B2(
        \regfile/reg_out[4][20] ), .ZN(n6260) );
  INV_X1 U5154 ( .A(n6261), .ZN(n5582) );
  AOI22_X1 U5156 ( .A1(n6091), .A2(n6265), .B1(\Mpath/N190 ), .B2(n6266), .ZN(
        n6264) );
  OAI221_X1 U5157 ( .B1(n6049), .B2(n6255), .C1(n5883), .C2(n7255), .A(n6254), 
        .ZN(n6267) );
  AOI22_X1 U5158 ( .A1(n7603), .A2(\regfile/reg_out[19][19] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][19] ), .ZN(n6269) );
  AOI22_X1 U5159 ( .A1(n7502), .A2(\regfile/reg_out[21][19] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][19] ), .ZN(n6270) );
  AOI22_X1 U5160 ( .A1(n5637), .A2(\regfile/reg_out[25][19] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][19] ), .ZN(n6271) );
  AOI22_X1 U5161 ( .A1(n5642), .A2(\regfile/reg_out[29][19] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][19] ), .ZN(n6272) );
  AOI22_X1 U5162 ( .A1(n5649), .A2(\regfile/reg_out[5][19] ), .B1(n5650), .B2(
        \regfile/reg_out[4][19] ), .ZN(n6273) );
  INV_X1 U5163 ( .A(n6274), .ZN(n5588) );
  AOI22_X1 U5165 ( .A1(n6091), .A2(n6278), .B1(\Mpath/N190 ), .B2(n6279), .ZN(
        n6277) );
  OAI221_X1 U5166 ( .B1(n6255), .B2(n6042), .C1(n5892), .C2(n7454), .A(n6254), 
        .ZN(n6280) );
  AND2_X1 U5167 ( .A1(n6281), .A2(n6282), .ZN(n6254) );
  NAND3_X1 U5168 ( .A1(net56319), .A2(net57730), .A3(n6045), .ZN(n6282) );
  NAND2_X1 U5169 ( .A1(n6067), .A2(\Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n6255) );
  AOI22_X1 U5170 ( .A1(n7603), .A2(\regfile/reg_out[19][18] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][18] ), .ZN(n6284) );
  AOI22_X1 U5171 ( .A1(n7502), .A2(\regfile/reg_out[21][18] ), .B1(n7611), 
        .B2(\regfile/reg_out[20][18] ), .ZN(n6285) );
  AOI22_X1 U5172 ( .A1(n5637), .A2(\regfile/reg_out[25][18] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][18] ), .ZN(n6286) );
  AOI22_X1 U5173 ( .A1(n5642), .A2(\regfile/reg_out[29][18] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][18] ), .ZN(n6287) );
  AOI22_X1 U5174 ( .A1(n5649), .A2(\regfile/reg_out[5][18] ), .B1(n5650), .B2(
        \regfile/reg_out[4][18] ), .ZN(n6288) );
  INV_X1 U5175 ( .A(n6289), .ZN(n5591) );
  AOI22_X1 U5177 ( .A1(n6091), .A2(n6293), .B1(\Mpath/N190 ), .B2(n6294), .ZN(
        n6292) );
  OAI221_X1 U5178 ( .B1(n7255), .B2(n5903), .C1(n6296), .C2(n5846), .A(n6281), 
        .ZN(n6295) );
  INV_X1 U5179 ( .A(n7567), .ZN(n6296) );
  AOI22_X1 U5180 ( .A1(n7603), .A2(\regfile/reg_out[19][17] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][17] ), .ZN(n6298) );
  AOI22_X1 U5181 ( .A1(n7502), .A2(\regfile/reg_out[21][17] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][17] ), .ZN(n6299) );
  AOI22_X1 U5182 ( .A1(n5637), .A2(\regfile/reg_out[25][17] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][17] ), .ZN(n6300) );
  AOI22_X1 U5183 ( .A1(n5642), .A2(\regfile/reg_out[29][17] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][17] ), .ZN(n6301) );
  AOI22_X1 U5184 ( .A1(n5649), .A2(\regfile/reg_out[5][17] ), .B1(n5650), .B2(
        \regfile/reg_out[4][17] ), .ZN(n6302) );
  INV_X1 U5185 ( .A(n6303), .ZN(n5594) );
  AOI22_X1 U5187 ( .A1(n6091), .A2(n6307), .B1(\Mpath/N190 ), .B2(n6308), .ZN(
        n6306) );
  OAI221_X1 U5188 ( .B1(n7176), .B2(n6047), .C1(n5913), .C2(n7454), .A(n6281), 
        .ZN(n6309) );
  AOI22_X1 U5189 ( .A1(n7603), .A2(\regfile/reg_out[19][16] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][16] ), .ZN(n6310) );
  AOI22_X1 U5190 ( .A1(n7503), .A2(\regfile/reg_out[21][16] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][16] ), .ZN(n6311) );
  AOI22_X1 U5191 ( .A1(n5637), .A2(\regfile/reg_out[25][16] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][16] ), .ZN(n6312) );
  AOI22_X1 U5192 ( .A1(n5642), .A2(\regfile/reg_out[29][16] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][16] ), .ZN(n6313) );
  AOI22_X1 U5193 ( .A1(n5649), .A2(\regfile/reg_out[5][16] ), .B1(n5650), .B2(
        \regfile/reg_out[4][16] ), .ZN(n6314) );
  INV_X1 U5194 ( .A(n6315), .ZN(n5597) );
  AOI22_X1 U5196 ( .A1(n6091), .A2(n6319), .B1(\Mpath/N190 ), .B2(n6320), .ZN(
        n6318) );
  NOR2_X1 U5198 ( .A1(n5846), .A2(n7434), .ZN(n6268) );
  OAI221_X1 U5199 ( .B1(n7176), .B2(n6048), .C1(n6052), .C2(n7454), .A(n6281), 
        .ZN(n6322) );
  NAND2_X1 U5200 ( .A1(\Mcontrol/Operation_decoding32/N1976 ), .A2(n6045), 
        .ZN(n6281) );
  AOI22_X1 U5201 ( .A1(n7603), .A2(\regfile/reg_out[19][15] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][15] ), .ZN(n6323) );
  AOI22_X1 U5202 ( .A1(n7503), .A2(\regfile/reg_out[21][15] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][15] ), .ZN(n6324) );
  AOI22_X1 U5203 ( .A1(n5637), .A2(\regfile/reg_out[25][15] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][15] ), .ZN(n6325) );
  AOI22_X1 U5204 ( .A1(n5642), .A2(\regfile/reg_out[29][15] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][15] ), .ZN(n6326) );
  AOI22_X1 U5205 ( .A1(n5649), .A2(\regfile/reg_out[5][15] ), .B1(n5650), .B2(
        \regfile/reg_out[4][15] ), .ZN(n6327) );
  INV_X1 U5206 ( .A(n6328), .ZN(n5600) );
  AOI22_X1 U5208 ( .A1(n6091), .A2(n6332), .B1(\Mpath/N190 ), .B2(n6333), .ZN(
        n6331) );
  AOI22_X1 U5210 ( .A1(n7603), .A2(\regfile/reg_out[19][14] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][14] ), .ZN(n6335) );
  AOI22_X1 U5211 ( .A1(n7503), .A2(\regfile/reg_out[21][14] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][14] ), .ZN(n6336) );
  AOI22_X1 U5212 ( .A1(n5637), .A2(\regfile/reg_out[25][14] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][14] ), .ZN(n6337) );
  AOI22_X1 U5213 ( .A1(n5642), .A2(\regfile/reg_out[29][14] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][14] ), .ZN(n6338) );
  AOI22_X1 U5214 ( .A1(n5649), .A2(\regfile/reg_out[5][14] ), .B1(n5650), .B2(
        \regfile/reg_out[4][14] ), .ZN(n6339) );
  INV_X1 U5215 ( .A(n6340), .ZN(n5603) );
  AOI22_X1 U5217 ( .A1(n6091), .A2(n6344), .B1(\Mpath/N190 ), .B2(n6345), .ZN(
        n6343) );
  AOI22_X1 U5219 ( .A1(n7603), .A2(\regfile/reg_out[19][13] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][13] ), .ZN(n6347) );
  AOI22_X1 U5220 ( .A1(n7502), .A2(\regfile/reg_out[21][13] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][13] ), .ZN(n6348) );
  AOI22_X1 U5221 ( .A1(n5637), .A2(\regfile/reg_out[25][13] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][13] ), .ZN(n6349) );
  AOI22_X1 U5222 ( .A1(n5642), .A2(\regfile/reg_out[29][13] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][13] ), .ZN(n6350) );
  AOI22_X1 U5223 ( .A1(n5649), .A2(\regfile/reg_out[5][13] ), .B1(n5650), .B2(
        \regfile/reg_out[4][13] ), .ZN(n6351) );
  INV_X1 U5224 ( .A(n6352), .ZN(n5606) );
  AOI22_X1 U5226 ( .A1(n6091), .A2(n6356), .B1(\Mpath/N190 ), .B2(n6357), .ZN(
        n6355) );
  OAI222_X1 U5227 ( .A1(n7255), .A2(n6039), .B1(n7176), .B2(n5894), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n6050), .ZN(n6358) );
  AOI22_X1 U5228 ( .A1(n7603), .A2(\regfile/reg_out[19][12] ), .B1(n7592), 
        .B2(\regfile/reg_out[18][12] ), .ZN(n6359) );
  AOI22_X1 U5231 ( .A1(n5642), .A2(\regfile/reg_out[29][12] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][12] ), .ZN(n6362) );
  AOI22_X1 U5232 ( .A1(n5649), .A2(\regfile/reg_out[5][12] ), .B1(n5650), .B2(
        \regfile/reg_out[4][12] ), .ZN(n6363) );
  INV_X1 U5233 ( .A(n6364), .ZN(n5609) );
  AOI22_X1 U5235 ( .A1(n6091), .A2(n6368), .B1(\Mpath/N190 ), .B2(n6369), .ZN(
        n6367) );
  AOI22_X1 U5237 ( .A1(n7603), .A2(\regfile/reg_out[19][11] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][11] ), .ZN(n6371) );
  AOI22_X1 U5238 ( .A1(n7503), .A2(\regfile/reg_out[21][11] ), .B1(n5633), 
        .B2(\regfile/reg_out[20][11] ), .ZN(n6372) );
  AOI22_X1 U5239 ( .A1(n5637), .A2(\regfile/reg_out[25][11] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][11] ), .ZN(n6373) );
  AOI22_X1 U5240 ( .A1(n5642), .A2(\regfile/reg_out[29][11] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][11] ), .ZN(n6374) );
  AOI22_X1 U5241 ( .A1(n5649), .A2(\regfile/reg_out[5][11] ), .B1(n5650), .B2(
        \regfile/reg_out[4][11] ), .ZN(n6375) );
  INV_X1 U5242 ( .A(n6376), .ZN(n5612) );
  AOI22_X1 U5244 ( .A1(n6091), .A2(n6380), .B1(\Mpath/N190 ), .B2(n6381), .ZN(
        n6379) );
  OAI222_X1 U5245 ( .A1(n7255), .A2(n6042), .B1(n7176), .B2(n5914), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n5894), .ZN(n6383) );
  INV_X1 U5250 ( .A(n6321), .ZN(n6105) );
  AOI22_X1 U5251 ( .A1(n7603), .A2(\regfile/reg_out[19][10] ), .B1(n5628), 
        .B2(\regfile/reg_out[18][10] ), .ZN(n6385) );
  AOI22_X1 U5252 ( .A1(n7502), .A2(\regfile/reg_out[21][10] ), .B1(n7514), 
        .B2(\regfile/reg_out[20][10] ), .ZN(n6386) );
  AOI22_X1 U5253 ( .A1(n5637), .A2(\regfile/reg_out[25][10] ), .B1(n5638), 
        .B2(\regfile/reg_out[24][10] ), .ZN(n6387) );
  AOI22_X1 U5254 ( .A1(n5642), .A2(\regfile/reg_out[29][10] ), .B1(n5643), 
        .B2(\regfile/reg_out[28][10] ), .ZN(n6388) );
  AOI22_X1 U5255 ( .A1(n5649), .A2(\regfile/reg_out[5][10] ), .B1(n5650), .B2(
        \regfile/reg_out[4][10] ), .ZN(n6389) );
  INV_X1 U5256 ( .A(n6390), .ZN(n5615) );
  AOI22_X1 U5258 ( .A1(n6091), .A2(n6394), .B1(\Mpath/N190 ), .B2(n6395), .ZN(
        n6393) );
  NAND2_X1 U5261 ( .A1(\Mpath/N186 ), .A2(n5657), .ZN(n5720) );
  INV_X1 U5268 ( .A(\Mcontrol/Nextpc_decoding/N319 ), .ZN(n6402) );
  INV_X1 U5272 ( .A(\Mcontrol/Nextpc_decoding/N307 ), .ZN(n6407) );
  OAI22_X1 U5273 ( .A1(n7298), .A2(n6409), .B1(n6410), .B2(
        \Mcontrol/Nextpc_decoding/N301 ), .ZN(n6406) );
  INV_X1 U5276 ( .A(\Mcontrol/Nextpc_decoding/N301 ), .ZN(n6409) );
  NAND3_X1 U5289 ( .A1(n6414), .A2(rs1_addr[2]), .A3(n6417), .ZN(n5630) );
  NAND3_X1 U5296 ( .A1(rs1_addr[1]), .A2(n6425), .A3(n7327), .ZN(n5634) );
  NOR2_X1 U5302 ( .A1(n6422), .A2(n7675), .ZN(n6425) );
  INV_X1 U5323 ( .A(rs1_addr[1]), .ZN(n6416) );
  OAI22_X1 U5336 ( .A1(n6436), .A2(n5657), .B1(n6437), .B2(n5659), .ZN(n6435)
         );
  INV_X1 U5337 ( .A(n6091), .ZN(n5659) );
  INV_X1 U5339 ( .A(\Mpath/N190 ), .ZN(n5657) );
  INV_X1 U5340 ( .A(\Mcontrol/Nextpc_decoding/N313 ), .ZN(n6404) );
  INV_X1 U5341 ( .A(\Mcontrol/Nextpc_decoding/N325 ), .ZN(n6399) );
  OAI22_X1 U5342 ( .A1(n6438), .A2(n6439), .B1(n5505), .B2(n6440), .ZN(
        D_DATA_OUTBUS[9]) );
  OAI22_X1 U5343 ( .A1(n6439), .A2(n6441), .B1(n5505), .B2(n6442), .ZN(
        D_DATA_OUTBUS[8]) );
  OAI221_X1 U5344 ( .B1(n6443), .B2(n6444), .C1(n6439), .C2(n6445), .A(n6446), 
        .ZN(D_DATA_OUTBUS[31]) );
  NAND2_X1 U5345 ( .A1(\Mpath/the_memhandle/smdr_out[31] ), .A2(n6447), .ZN(
        n6446) );
  OAI221_X1 U5346 ( .B1(n6443), .B2(n6448), .C1(n6439), .C2(n6449), .A(n6450), 
        .ZN(D_DATA_OUTBUS[30]) );
  NAND2_X1 U5347 ( .A1(\Mpath/the_memhandle/smdr_out[30] ), .A2(n6447), .ZN(
        n6450) );
  OAI221_X1 U5348 ( .B1(n6443), .B2(n6451), .C1(n6439), .C2(n6452), .A(n6453), 
        .ZN(D_DATA_OUTBUS[29]) );
  NAND2_X1 U5349 ( .A1(\Mpath/the_memhandle/smdr_out[29] ), .A2(n6447), .ZN(
        n6453) );
  OAI221_X1 U5350 ( .B1(n6443), .B2(n6454), .C1(n6439), .C2(n6455), .A(n6456), 
        .ZN(D_DATA_OUTBUS[28]) );
  NAND2_X1 U5351 ( .A1(\Mpath/the_memhandle/smdr_out[28] ), .A2(n6447), .ZN(
        n6456) );
  OAI221_X1 U5352 ( .B1(n6443), .B2(n6457), .C1(n6439), .C2(n6458), .A(n6459), 
        .ZN(D_DATA_OUTBUS[27]) );
  NAND2_X1 U5353 ( .A1(\Mpath/the_memhandle/smdr_out[27] ), .A2(n6447), .ZN(
        n6459) );
  OAI221_X1 U5354 ( .B1(n6443), .B2(n6460), .C1(n6439), .C2(n6461), .A(n6462), 
        .ZN(D_DATA_OUTBUS[26]) );
  NAND2_X1 U5355 ( .A1(\Mpath/the_memhandle/smdr_out[26] ), .A2(n6447), .ZN(
        n6462) );
  OAI221_X1 U5356 ( .B1(n6443), .B2(n6440), .C1(n6438), .C2(n6439), .A(n6463), 
        .ZN(D_DATA_OUTBUS[25]) );
  NAND2_X1 U5357 ( .A1(\Mpath/the_memhandle/smdr_out[25] ), .A2(n6447), .ZN(
        n6463) );
  OAI221_X1 U5358 ( .B1(n6443), .B2(n6442), .C1(n6439), .C2(n6441), .A(n6464), 
        .ZN(D_DATA_OUTBUS[24]) );
  NAND2_X1 U5359 ( .A1(\Mpath/the_memhandle/smdr_out[24] ), .A2(n6447), .ZN(
        n6464) );
  OAI21_X1 U5360 ( .B1(n6465), .B2(n6445), .A(n6466), .ZN(D_DATA_OUTBUS[23])
         );
  NAND2_X1 U5361 ( .A1(\Mpath/the_memhandle/smdr_out[23] ), .A2(n6447), .ZN(
        n6466) );
  OAI21_X1 U5362 ( .B1(n6465), .B2(n6449), .A(n6467), .ZN(D_DATA_OUTBUS[22])
         );
  NAND2_X1 U5363 ( .A1(\Mpath/the_memhandle/smdr_out[22] ), .A2(n6447), .ZN(
        n6467) );
  OAI21_X1 U5364 ( .B1(n6465), .B2(n6452), .A(n6468), .ZN(D_DATA_OUTBUS[21])
         );
  NAND2_X1 U5365 ( .A1(\Mpath/the_memhandle/smdr_out[21] ), .A2(n6447), .ZN(
        n6468) );
  OAI21_X1 U5366 ( .B1(n6465), .B2(n6455), .A(n6469), .ZN(D_DATA_OUTBUS[20])
         );
  NAND2_X1 U5367 ( .A1(\Mpath/the_memhandle/smdr_out[20] ), .A2(n6447), .ZN(
        n6469) );
  OAI21_X1 U5368 ( .B1(n6465), .B2(n6458), .A(n6470), .ZN(D_DATA_OUTBUS[19])
         );
  NAND2_X1 U5369 ( .A1(\Mpath/the_memhandle/smdr_out[19] ), .A2(n6447), .ZN(
        n6470) );
  OAI21_X1 U5370 ( .B1(n6465), .B2(n6461), .A(n6471), .ZN(D_DATA_OUTBUS[18])
         );
  NAND2_X1 U5371 ( .A1(\Mpath/the_memhandle/smdr_out[18] ), .A2(n6447), .ZN(
        n6471) );
  OAI21_X1 U5372 ( .B1(n6465), .B2(n6438), .A(n6472), .ZN(D_DATA_OUTBUS[17])
         );
  NAND2_X1 U5373 ( .A1(\Mpath/the_memhandle/smdr_out[17] ), .A2(n6447), .ZN(
        n6472) );
  OAI21_X1 U5374 ( .B1(n6465), .B2(n6441), .A(n6473), .ZN(D_DATA_OUTBUS[16])
         );
  NAND2_X1 U5375 ( .A1(\Mpath/the_memhandle/smdr_out[16] ), .A2(n6447), .ZN(
        n6473) );
  NOR2_X1 U5376 ( .A1(\d_chk/N10 ), .A2(n6474), .ZN(n6465) );
  OAI22_X1 U5377 ( .A1(n6439), .A2(n6445), .B1(n5505), .B2(n6444), .ZN(
        D_DATA_OUTBUS[15]) );
  OAI22_X1 U5378 ( .A1(n6439), .A2(n6449), .B1(n5505), .B2(n6448), .ZN(
        D_DATA_OUTBUS[14]) );
  OAI22_X1 U5379 ( .A1(n6439), .A2(n6452), .B1(n5505), .B2(n6451), .ZN(
        D_DATA_OUTBUS[13]) );
  OAI22_X1 U5380 ( .A1(n6439), .A2(n6455), .B1(n5505), .B2(n6454), .ZN(
        D_DATA_OUTBUS[12]) );
  OAI22_X1 U5381 ( .A1(n6439), .A2(n6458), .B1(n5505), .B2(n6457), .ZN(
        D_DATA_OUTBUS[11]) );
  OAI22_X1 U5382 ( .A1(n6439), .A2(n6461), .B1(n5505), .B2(n6460), .ZN(
        D_DATA_OUTBUS[10]) );
  INV_X1 U5383 ( .A(\d_chk/N10 ), .ZN(n6439) );
  AND2_X1 U5384 ( .A1(n6117), .A2(n6475), .ZN(D_ADDR_OUTBUS[9]) );
  AND2_X1 U5385 ( .A1(n6130), .A2(n6475), .ZN(D_ADDR_OUTBUS[8]) );
  OAI22_X1 U5386 ( .A1(n4509), .A2(n5504), .B1(n6476), .B2(n6477), .ZN(
        D_ADDR_OUTBUS[7]) );
  INV_X1 U5387 ( .A(n6142), .ZN(n6476) );
  NAND2_X1 U5388 ( .A1(\Scc_coproc/ein_exc_word[5] ), .A2(n6479), .ZN(n6478)
         );
  OAI22_X1 U5389 ( .A1(n4510), .A2(n5504), .B1(n6480), .B2(n6477), .ZN(
        D_ADDR_OUTBUS[6]) );
  INV_X1 U5390 ( .A(n6154), .ZN(n6480) );
  INV_X1 U5391 ( .A(n6481), .ZN(D_ADDR_OUTBUS[5]) );
  AOI22_X1 U5392 ( .A1(serve_proc_addr[5]), .A2(n7109), .B1(n6166), .B2(n6475), 
        .ZN(n6481) );
  INV_X1 U5393 ( .A(n6483), .ZN(D_ADDR_OUTBUS[4]) );
  AOI22_X1 U5394 ( .A1(serve_proc_addr[4]), .A2(n7109), .B1(n6183), .B2(n6475), 
        .ZN(n6483) );
  INV_X1 U5395 ( .A(n6486), .ZN(D_ADDR_OUTBUS[3]) );
  AOI22_X1 U5396 ( .A1(serve_proc_addr[3]), .A2(n7109), .B1(n6197), .B2(n6475), 
        .ZN(n6486) );
  NOR2_X1 U5397 ( .A1(n6437), .A2(n6477), .ZN(D_ADDR_OUTBUS[31]) );
  NOR2_X1 U5398 ( .A1(n5658), .A2(n6477), .ZN(D_ADDR_OUTBUS[30]) );
  INV_X1 U5399 ( .A(n6488), .ZN(D_ADDR_OUTBUS[2]) );
  AOI22_X1 U5400 ( .A1(serve_proc_addr[2]), .A2(n7109), .B1(n6212), .B2(n6475), 
        .ZN(n6488) );
  AOI21_X1 U5401 ( .B1(n5741), .B2(n6491), .A(\Scc_coproc/interrupt[6] ), .ZN(
        n6490) );
  OAI21_X1 U5402 ( .B1(n6492), .B2(\Scc_coproc/interrupt[3] ), .A(n5742), .ZN(
        n6491) );
  INV_X1 U5403 ( .A(\Scc_coproc/interrupt[5] ), .ZN(n5741) );
  INV_X1 U5406 ( .A(\d_chk/N13 ), .ZN(n6495) );
  INV_X1 U5408 ( .A(n6443), .ZN(n6474) );
  NAND2_X1 U5409 ( .A1(\d_chk/N11 ), .A2(\x_mem_command[MB] ), .ZN(n6443) );
  NOR2_X1 U5414 ( .A1(n5667), .A2(n6477), .ZN(D_ADDR_OUTBUS[29]) );
  NOR2_X1 U5415 ( .A1(n5675), .A2(n6477), .ZN(D_ADDR_OUTBUS[28]) );
  NOR2_X1 U5416 ( .A1(n5683), .A2(n6477), .ZN(D_ADDR_OUTBUS[27]) );
  NOR2_X1 U5417 ( .A1(n5691), .A2(n6477), .ZN(D_ADDR_OUTBUS[26]) );
  NOR2_X1 U5418 ( .A1(n5699), .A2(n6477), .ZN(D_ADDR_OUTBUS[25]) );
  NOR2_X1 U5419 ( .A1(n5707), .A2(n6477), .ZN(D_ADDR_OUTBUS[24]) );
  AND2_X1 U5420 ( .A1(n6225), .A2(n6475), .ZN(D_ADDR_OUTBUS[23]) );
  AND2_X1 U5421 ( .A1(n6237), .A2(n6475), .ZN(D_ADDR_OUTBUS[22]) );
  AND2_X1 U5422 ( .A1(n6249), .A2(n6475), .ZN(D_ADDR_OUTBUS[21]) );
  AND2_X1 U5423 ( .A1(n6265), .A2(n6475), .ZN(D_ADDR_OUTBUS[20]) );
  AND2_X1 U5424 ( .A1(n6968), .A2(n6475), .ZN(D_ADDR_OUTBUS[1]) );
  AND2_X1 U5425 ( .A1(n6278), .A2(n6475), .ZN(D_ADDR_OUTBUS[19]) );
  AND2_X1 U5426 ( .A1(n6293), .A2(n6475), .ZN(D_ADDR_OUTBUS[18]) );
  AND2_X1 U5427 ( .A1(n6307), .A2(n6475), .ZN(D_ADDR_OUTBUS[17]) );
  AND2_X1 U5428 ( .A1(n6319), .A2(n6475), .ZN(D_ADDR_OUTBUS[16]) );
  AND2_X1 U5429 ( .A1(n6332), .A2(n6475), .ZN(D_ADDR_OUTBUS[15]) );
  OAI21_X1 U5430 ( .B1(n6498), .B2(n6477), .A(n5504), .ZN(D_ADDR_OUTBUS[14])
         );
  INV_X1 U5431 ( .A(n7110), .ZN(n5504) );
  INV_X1 U5432 ( .A(n6344), .ZN(n6498) );
  AND2_X1 U5433 ( .A1(n6356), .A2(n6475), .ZN(D_ADDR_OUTBUS[13]) );
  AND2_X1 U5434 ( .A1(n6368), .A2(n6475), .ZN(D_ADDR_OUTBUS[12]) );
  AND2_X1 U5435 ( .A1(n6380), .A2(n6475), .ZN(D_ADDR_OUTBUS[11]) );
  AND2_X1 U5436 ( .A1(n6394), .A2(n6475), .ZN(D_ADDR_OUTBUS[10]) );
  INV_X1 U5437 ( .A(n6477), .ZN(n6475) );
  NOR2_X1 U5438 ( .A1(n5714), .A2(n6477), .ZN(D_ADDR_OUTBUS[0]) );
  NAND2_X1 U5439 ( .A1(N5), .A2(serve_exception), .ZN(n6477) );
  INV_X1 U5441 ( .A(\Mpath/the_alu/N492 ), .ZN(n6501) );
  NOR3_X1 U5443 ( .A1(\Mpath/the_shift/N115 ), .A2(\Mpath/the_shift/N118 ), 
        .A3(\Mpath/the_shift/N111 ), .ZN(n6503) );
  OAI21_X1 U5444 ( .B1(\Mpath/the_alu/N492 ), .B2(n6505), .A(n6506), .ZN(n6504) );
  NAND2_X1 U5445 ( .A1(\Mpath/the_alu/N125 ), .A2(\Mpath/the_alu/N492 ), .ZN(
        n6506) );
  AOI22_X1 U5446 ( .A1(n6507), .A2(\Mpath/the_alu/N485 ), .B1(
        \Mpath/the_alu/N157 ), .B2(\Mpath/the_alu/N486 ), .ZN(n6505) );
  OAI21_X1 U5447 ( .B1(\Mpath/the_alu/N480 ), .B2(n6508), .A(n6509), .ZN(n6507) );
  NAND2_X1 U5448 ( .A1(\Mpath/the_alu/N189 ), .A2(\Mpath/the_alu/N480 ), .ZN(
        n6509) );
  AOI22_X1 U5449 ( .A1(\Mpath/the_alu/N221 ), .A2(\Mpath/the_alu/N474 ), .B1(
        \Mpath/the_alu/N473 ), .B2(\Mpath/out_regA[0] ), .ZN(n6508) );
  OAI21_X1 U5450 ( .B1(n6511), .B2(n6075), .A(n7552), .ZN(n6510) );
  AOI211_X1 U5452 ( .C1(n6060), .C2(n7576), .A(n7441), .B(n6067), .ZN(n6511)
         );
  CLKBUF_X2 U5455 ( .A(n6512), .Z(\Mpath/the_alu/N1 ) );
  Xi_core_DW01_add_0 \Mcontrol/Nextpc_decoding/bta_calc/add_391  ( .A({1'b0, 
        \Mcontrol/f_currpc[23] , \Mcontrol/f_currpc[22] , 
        \Mcontrol/f_currpc[21] , \Mcontrol/f_currpc[20] , 
        \Mcontrol/f_currpc[19] , \Mcontrol/f_currpc[18] , 
        \Mcontrol/f_currpc[17] , \Mcontrol/f_currpc[16] , 
        \Mcontrol/f_currpc[15] , \Mcontrol/f_currpc[14] , 
        \Mcontrol/f_currpc[13] , \Mcontrol/f_currpc[12] , 
        \Mcontrol/f_currpc[11] , \Mcontrol/f_currpc[10] , 
        \Mcontrol/f_currpc[9] , \Mcontrol/f_currpc[8] , \Mcontrol/f_currpc[7] , 
        \Mcontrol/f_currpc[6] , \Mcontrol/f_currpc[5] , \Mcontrol/f_currpc[4] , 
        \Mcontrol/f_currpc[3] , \Mcontrol/f_currpc[2] , \Mcontrol/f_currpc[1] , 
        \Mcontrol/f_currpc[0] }), .B({1'b0, break_code[23:16], n6551, 
        break_code[14:0]}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        \Mcontrol/Nextpc_decoding/Bta }) );
  Xi_core_DW01_add_1 \Mcontrol/Nextpc_decoding/incr/add_391  ( .A({1'b0, 
        \Mcontrol/f_currpc[23] , \Mcontrol/f_currpc[22] , 
        \Mcontrol/f_currpc[21] , \Mcontrol/f_currpc[20] , 
        \Mcontrol/f_currpc[19] , \Mcontrol/f_currpc[18] , 
        \Mcontrol/f_currpc[17] , \Mcontrol/f_currpc[16] , 
        \Mcontrol/f_currpc[15] , \Mcontrol/f_currpc[14] , 
        \Mcontrol/f_currpc[13] , \Mcontrol/f_currpc[12] , 
        \Mcontrol/f_currpc[11] , \Mcontrol/f_currpc[10] , 
        \Mcontrol/f_currpc[9] , \Mcontrol/f_currpc[8] , \Mcontrol/f_currpc[7] , 
        \Mcontrol/f_currpc[6] , \Mcontrol/f_currpc[5] , \Mcontrol/f_currpc[4] , 
        \Mcontrol/f_currpc[3] , \Mcontrol/f_currpc[2] , \Mcontrol/f_currpc[1] , 
        \Mcontrol/f_currpc[0] }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, jar_in}) );
  Xi_core_DW01_sub_1 \Mpath/the_alu/sub_96  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        \Mpath/out_regA[12] , \Mpath/out_regA[11] , \Mpath/out_regA[10] , 
        \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , 
        \Mpath/out_regA[5] , \Mpath/out_regA[4] , \Mpath/out_regA[3] , 
        \Mpath/out_regA[2] , \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .B({
        \Mpath/out_regB[31] , \Mpath/out_regB[30] , \Mpath/out_regB[29] , 
        \Mpath/out_regB[28] , \Mpath/out_regB[27] , \Mpath/out_regB[26] , 
        \Mpath/out_regB[25] , \Mpath/out_regB[24] , \Mpath/out_regB[23] , 
        \Mpath/out_regB[22] , \Mpath/out_regB[21] , \Mpath/out_regB[20] , 
        n7331, n7359, n7343, n7386, n7322, n7393, n7105, \Mpath/out_regB[12] , 
        \Mpath/out_regB[11] , \Mpath/out_regB[10] , \Mpath/out_regB[9] , n7614, 
        \Mpath/out_regB[7] , \Mpath/out_regB[6] , \Mpath/out_regB[5] , n7707, 
        n7708, n7711, n7713, n7715}), .DIFF({\Mpath/the_alu/diff[31] , 
        \Mpath/the_alu/diff[30] , \Mpath/the_alu/diff[29] , 
        \Mpath/the_alu/diff[28] , \Mpath/the_alu/diff[27] , 
        \Mpath/the_alu/diff[26] , \Mpath/the_alu/diff[25] , 
        \Mpath/the_alu/diff[24] , \Mpath/the_alu/diff[23] , 
        \Mpath/the_alu/diff[22] , \Mpath/the_alu/diff[21] , 
        \Mpath/the_alu/diff[20] , \Mpath/the_alu/diff[19] , 
        \Mpath/the_alu/diff[18] , \Mpath/the_alu/diff[17] , 
        \Mpath/the_alu/diff[16] , \Mpath/the_alu/diff[15] , 
        \Mpath/the_alu/diff[14] , \Mpath/the_alu/diff[13] , 
        \Mpath/the_alu/diff[12] , \Mpath/the_alu/diff[11] , 
        \Mpath/the_alu/diff[10] , \Mpath/the_alu/diff[9] , 
        \Mpath/the_alu/diff[8] , \Mpath/the_alu/diff[7] , 
        \Mpath/the_alu/diff[6] , \Mpath/the_alu/diff[5] , 
        \Mpath/the_alu/diff[4] , \Mpath/the_alu/diff[3] , 
        \Mpath/the_alu/diff[2] , \Mpath/the_alu/diff[1] , 
        \Mpath/the_alu/diff[0] }), .CI(1'b0) );
  Xi_core_DW01_add_3 \Mpath/the_alu/add_95  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        \Mpath/out_regA[12] , \Mpath/out_regA[11] , \Mpath/out_regA[10] , 
        \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , 
        \Mpath/out_regA[5] , \Mpath/out_regA[4] , \Mpath/out_regA[3] , 
        \Mpath/out_regA[2] , \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .B({
        \Mpath/out_regB[31] , \Mpath/out_regB[30] , \Mpath/out_regB[29] , 
        \Mpath/out_regB[28] , \Mpath/out_regB[27] , \Mpath/out_regB[26] , 
        \Mpath/out_regB[25] , \Mpath/out_regB[24] , \Mpath/out_regB[23] , 
        \Mpath/out_regB[22] , \Mpath/out_regB[21] , \Mpath/out_regB[20] , 
        n7332, n7360, n7344, n7387, n7323, n7394, n7106, \Mpath/out_regB[12] , 
        \Mpath/out_regB[11] , \Mpath/out_regB[10] , \Mpath/out_regB[9] , n7615, 
        \Mpath/out_regB[7] , \Mpath/out_regB[6] , \Mpath/out_regB[5] , n7706, 
        n7708, n7710, n7712, n7715}), .SUM({\Mpath/the_alu/sum[31] , 
        \Mpath/the_alu/sum[30] , \Mpath/the_alu/sum[29] , 
        \Mpath/the_alu/sum[28] , \Mpath/the_alu/sum[27] , 
        \Mpath/the_alu/sum[26] , \Mpath/the_alu/sum[25] , 
        \Mpath/the_alu/sum[24] , \Mpath/the_alu/sum[23] , 
        \Mpath/the_alu/sum[22] , \Mpath/the_alu/sum[21] , 
        \Mpath/the_alu/sum[20] , \Mpath/the_alu/sum[19] , 
        \Mpath/the_alu/sum[18] , \Mpath/the_alu/sum[17] , 
        \Mpath/the_alu/sum[16] , \Mpath/the_alu/sum[15] , 
        \Mpath/the_alu/sum[14] , \Mpath/the_alu/sum[13] , 
        \Mpath/the_alu/sum[12] , \Mpath/the_alu/sum[11] , 
        \Mpath/the_alu/sum[10] , \Mpath/the_alu/sum[9] , 
        \Mpath/the_alu/sum[8] , \Mpath/the_alu/sum[7] , \Mpath/the_alu/sum[6] , 
        \Mpath/the_alu/sum[5] , \Mpath/the_alu/sum[4] , \Mpath/the_alu/sum[3] , 
        \Mpath/the_alu/sum[2] , \Mpath/the_alu/sum[1] , \Mpath/the_alu/sum[0] }), .CI(1'b0) );
  Xi_core_DW_rightsh_1 \Mpath/the_shift/S_SRL/srl_128  ( .A({
        \Mpath/out_regA[31] , \Mpath/out_regA[30] , \Mpath/out_regA[29] , 
        \Mpath/out_regA[28] , \Mpath/out_regA[27] , \Mpath/out_regA[26] , 
        \Mpath/out_regA[25] , \Mpath/out_regA[24] , \Mpath/out_regA[23] , 
        \Mpath/out_regA[22] , \Mpath/out_regA[21] , \Mpath/out_regA[20] , 
        \Mpath/out_regA[19] , \Mpath/out_regA[18] , \Mpath/out_regA[17] , 
        \Mpath/out_regA[16] , \Mpath/out_regA[15] , \Mpath/out_regA[14] , 
        \Mpath/out_regA[13] , n7182, \Mpath/out_regA[11] , 
        \Mpath/out_regA[10] , \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , 
        \Mpath/out_regA[6] , \Mpath/out_regA[5] , \Mpath/out_regA[4] , 
        \Mpath/out_regA[3] , \Mpath/out_regA[2] , \Mpath/out_regA[1] , 
        \Mpath/out_regA[0] }), .SH({n7706, n7708, n7711, n7713, n7714}), .B(
        \Mpath/the_shift/sh_srl ), .DATA_TC(1'b0) );
  Xi_core_DW_sra_1 \Mpath/the_shift/S_SRA/sra_106  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        n7182, \Mpath/out_regA[11] , \Mpath/out_regA[10] , \Mpath/out_regA[9] , 
        n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , \Mpath/out_regA[5] , 
        \Mpath/out_regA[4] , \Mpath/out_regA[3] , \Mpath/out_regA[2] , 
        \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .SH({n7706, n7708, n7709, 
        n7712, n7715}), .B(\Mpath/the_shift/sh_sra ), .SH_TC(1'b0) );
  Xi_core_DW_rbsh_1 \Mpath/the_shift/S_ROR/ror_81  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        \Mpath/out_regA[12] , \Mpath/out_regA[11] , \Mpath/out_regA[10] , 
        \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , 
        \Mpath/out_regA[5] , \Mpath/out_regA[4] , \Mpath/out_regA[3] , 
        \Mpath/out_regA[2] , \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .SH({
        n7706, n7708, n7710, n7712, n7714}), .B(\Mpath/the_shift/sh_ror ), 
        .SH_TC(1'b0) );
  Xi_core_DW01_bsh_1 \Mpath/the_shift/S_ROL/rol_55  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        \Mpath/out_regA[12] , \Mpath/out_regA[11] , \Mpath/out_regA[10] , 
        \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , 
        \Mpath/out_regA[5] , \Mpath/out_regA[4] , \Mpath/out_regA[3] , 
        \Mpath/out_regA[2] , \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .SH({
        n7706, n7708, n7709, n7712, n7714}), .B(\Mpath/the_shift/sh_rol ) );
  Xi_core_DW_leftsh_1 \Mpath/the_shift/S_SLL/sll_150  ( .A({
        \Mpath/out_regA[31] , \Mpath/out_regA[30] , \Mpath/out_regA[29] , 
        \Mpath/out_regA[28] , \Mpath/out_regA[27] , \Mpath/out_regA[26] , 
        \Mpath/out_regA[25] , \Mpath/out_regA[24] , \Mpath/out_regA[23] , 
        \Mpath/out_regA[22] , \Mpath/out_regA[21] , \Mpath/out_regA[20] , 
        \Mpath/out_regA[19] , \Mpath/out_regA[18] , \Mpath/out_regA[17] , 
        \Mpath/out_regA[16] , \Mpath/out_regA[15] , \Mpath/out_regA[14] , 
        \Mpath/out_regA[13] , n7182, \Mpath/out_regA[11] , 
        \Mpath/out_regA[10] , \Mpath/out_regA[9] , n7185, \Mpath/out_regA[7] , 
        \Mpath/out_regA[6] , \Mpath/out_regA[5] , \Mpath/out_regA[4] , 
        \Mpath/out_regA[3] , \Mpath/out_regA[2] , \Mpath/out_regA[1] , 
        \Mpath/out_regA[0] }), .SH({n7707, n7708, n7711, n7712, n7714}), .B(
        \Mpath/the_shift/sh_sll ) );
  Xi_core_DW_cmp_0 \Mpath/the_alu/lt_114  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        n7182, \Mpath/out_regA[11] , \Mpath/out_regA[10] , \Mpath/out_regA[9] , 
        n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , \Mpath/out_regA[5] , 
        \Mpath/out_regA[4] , \Mpath/out_regA[3] , \Mpath/out_regA[2] , 
        \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .B({\Mpath/out_regB[31] , 
        \Mpath/out_regB[30] , \Mpath/out_regB[29] , \Mpath/out_regB[28] , 
        \Mpath/out_regB[27] , \Mpath/out_regB[26] , \Mpath/out_regB[25] , 
        \Mpath/out_regB[24] , \Mpath/out_regB[23] , \Mpath/out_regB[22] , 
        \Mpath/out_regB[21] , n7476, n7333, n7361, n7344, n7388, n7323, n7395, 
        n7106, \Mpath/out_regB[12] , \Mpath/out_regB[11] , n7192, 
        \Mpath/out_regB[9] , n7616, \Mpath/out_regB[7] , \Mpath/out_regB[6] , 
        \Mpath/out_regB[5] , n7706, n7708, n7710, n7712, n7715}), .TC(1'b1), 
        .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(\Mpath/the_alu/N91 ) );
  Xi_core_DW_cmp_1 \Mpath/the_alu/lt_120  ( .A({\Mpath/out_regA[31] , 
        \Mpath/out_regA[30] , \Mpath/out_regA[29] , \Mpath/out_regA[28] , 
        \Mpath/out_regA[27] , \Mpath/out_regA[26] , \Mpath/out_regA[25] , 
        \Mpath/out_regA[24] , \Mpath/out_regA[23] , \Mpath/out_regA[22] , 
        \Mpath/out_regA[21] , \Mpath/out_regA[20] , \Mpath/out_regA[19] , 
        \Mpath/out_regA[18] , \Mpath/out_regA[17] , \Mpath/out_regA[16] , 
        \Mpath/out_regA[15] , \Mpath/out_regA[14] , \Mpath/out_regA[13] , 
        n7182, \Mpath/out_regA[11] , \Mpath/out_regA[10] , \Mpath/out_regA[9] , 
        n7185, \Mpath/out_regA[7] , \Mpath/out_regA[6] , \Mpath/out_regA[5] , 
        \Mpath/out_regA[4] , \Mpath/out_regA[3] , \Mpath/out_regA[2] , 
        \Mpath/out_regA[1] , \Mpath/out_regA[0] }), .B({\Mpath/out_regB[31] , 
        \Mpath/out_regB[30] , \Mpath/out_regB[29] , \Mpath/out_regB[28] , 
        \Mpath/out_regB[27] , \Mpath/out_regB[26] , \Mpath/out_regB[25] , 
        \Mpath/out_regB[24] , \Mpath/out_regB[23] , \Mpath/out_regB[22] , 
        \Mpath/out_regB[21] , n7476, n7332, n7360, n7344, n7387, n7323, n7394, 
        n7106, \Mpath/out_regB[12] , \Mpath/out_regB[11] , n7192, 
        \Mpath/out_regB[9] , n7615, \Mpath/out_regB[7] , \Mpath/out_regB[6] , 
        \Mpath/out_regB[5] , n7706, n7708, n7710, n7712, n7715}), .TC(1'b0), 
        .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(\Mpath/the_alu/N93 ) );
  Xi_core_DW01_cmp6_1 r772 ( .A({n7298, branch_rega[30:23], n6952, 
        branch_rega[21:9], n6893, branch_rega[7:0]}), .B(branch_regb), .TC(
        1'b0), .EQ(\Mcontrol/Nextpc_decoding/N26 ), .NE(
        \Mcontrol/Nextpc_decoding/N29 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[7]  ( .D(n3809), .CK(CLK), .RN(n7817), .Q(
        \Mpath/out_regA[7] ), .QN(\Mpath/the_alu/N69 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[5]  ( .D(n3725), .CK(CLK), .RN(n7797), .Q(
        \Mpath/out_regA[5] ), .QN(\Mpath/the_alu/N73 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[6]  ( .D(n3767), .CK(CLK), .RN(n7738), .Q(
        \Mpath/out_regA[6] ), .QN(\Mpath/the_alu/N71 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[16]  ( .D(n3453), .CK(CLK), .RN(n7791), .Q(
        \Mpath/out_regA[16] ), .QN(\Mpath/the_alu/N51 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[21]  ( .D(n3258), .CK(CLK), .RN(n7758), .Q(
        \Mpath/out_regA[21] ), .QN(\Mpath/the_alu/N41 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[31]  ( .D(n3910), .CK(CLK), .RN(n7753), .Q(
        \Mpath/out_regA[31] ), .QN(\Mpath/the_alu/N21 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[23]  ( .D(n3908), .CK(CLK), .RN(n7754), .Q(
        \Mpath/out_regA[23] ), .QN(\Mpath/the_alu/N37 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[3]  ( .D(n3911), .CK(CLK), .RN(n7800), .Q(
        \Mpath/out_regA[3] ), .QN(\Mpath/the_alu/N77 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[27]  ( .D(n4455), .CK(CLK), .RN(n7806), .Q(
        \Mpath/out_regA[27] ), .QN(\Mpath/the_alu/N29 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[22]  ( .D(n3219), .CK(CLK), .RN(n7812), .Q(
        \Mpath/out_regA[22] ), .QN(\Mpath/the_alu/N39 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[2]  ( .D(n3909), .CK(CLK), .RN(n7748), .Q(
        \Mpath/out_regA[2] ), .QN(\Mpath/the_alu/N79 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[4]  ( .D(n3912), .CK(CLK), .RN(n7717), .Q(
        \Mpath/out_regA[4] ), .QN(\Mpath/the_alu/N75 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[25]  ( .D(n3146), .CK(CLK), .RN(n7729), .Q(
        \Mpath/out_regA[25] ), .QN(\Mpath/the_alu/N33 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[29]  ( .D(n4459), .CK(CLK), .RN(n7741), .Q(
        \Mpath/out_regA[29] ), .QN(\Mpath/the_alu/N25 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[0]  ( .D(n4494), .CK(CLK), .RN(n7750), .Q(
        \Mpath/out_regA[0] ), .QN(\Mpath/the_alu/N83 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[26]  ( .D(n4453), .CK(CLK), .RN(n7820), .Q(
        \Mpath/out_regA[26] ), .QN(\Mpath/the_alu/N31 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[30]  ( .D(n4461), .CK(CLK), .RN(n7763), .Q(
        \Mpath/out_regA[30] ), .QN(\Mpath/the_alu/N23 ) );
  DFFR_X2 \regfile/rx_24/data_out_reg[31]  ( .D(n3959), .CK(CLK), .RN(n7742), 
        .Q(\regfile/reg_out[24][31] ), .QN(n4998) );
  DFFR_X2 \regfile/rx_25/data_out_reg[31]  ( .D(n4169), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[25][31] ), .QN(n4966) );
  DFFR_X2 \Mpath/regA/data_out_reg[24]  ( .D(n3180), .CK(CLK), .RN(n7809), .Q(
        \Mpath/out_regA[24] ), .QN(\Mpath/the_alu/N35 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[28]  ( .D(n4457), .CK(CLK), .RN(n7803), .Q(
        \Mpath/out_regA[28] ), .QN(\Mpath/the_alu/N27 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[1]  ( .D(n3907), .CK(CLK), .RN(n7720), .Q(
        \Mpath/out_regA[1] ), .QN(\Mpath/the_alu/N81 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[11]  ( .D(n3575), .CK(CLK), .RN(n7735), .Q(
        \Mpath/out_regA[11] ), .QN(\Mpath/the_alu/N61 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[15]  ( .D(n3495), .CK(CLK), .RN(n7776), .Q(
        \Mpath/out_regA[15] ), .QN(\Mpath/the_alu/N53 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[17]  ( .D(n3414), .CK(CLK), .RN(n7761), .Q(
        \Mpath/out_regA[17] ), .QN(\Mpath/the_alu/N49 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[18]  ( .D(n3375), .CK(CLK), .RN(n7815), .Q(
        \Mpath/out_regA[18] ), .QN(\Mpath/the_alu/N47 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[20]  ( .D(n3297), .CK(CLK), .RN(n7793), .Q(
        \Mpath/out_regA[20] ), .QN(\Mpath/the_alu/N43 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[10]  ( .D(n3536), .CK(CLK), .RN(n7779), .Q(
        \Mpath/out_regA[10] ), .QN(\Mpath/the_alu/N63 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[13]  ( .D(n3653), .CK(CLK), .RN(n7723), .Q(
        \Mpath/out_regA[13] ), .QN(\Mpath/the_alu/N57 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[14]  ( .D(n3906), .CK(CLK), .RN(n7770), .Q(
        \Mpath/out_regA[14] ), .QN(\Mpath/the_alu/N55 ) );
  DFFR_X2 \regfile/rx_18/data_out_reg[31]  ( .D(n4001), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[18][31] ), .QN(n5222) );
  DFFR_X2 \regfile/rx_19/data_out_reg[31]  ( .D(n4211), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[19][31] ), .QN(n5190) );
  DFFR_X1 \Mpath/regB/data_out_reg[18]  ( .D(n3374), .CK(CLK), .RN(n7814), .Q(
        \Mpath/out_regB[18] ), .QN(\Mpath/the_alu/N48 ) );
  DFFR_X2 \regfile/rx_20/data_out_reg[31]  ( .D(n3987), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[20][31] ), .QN(n5126) );
  DFFR_X2 \regfile/rx_21/data_out_reg[31]  ( .D(n4197), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[21][31] ), .QN(n5094) );
  DFFR_X2 \regfile/rx_4/data_out_reg[31]  ( .D(n4099), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[4][31] ), .QN(n4678) );
  DFFR_X2 \regfile/rx_5/data_out_reg[31]  ( .D(n4309), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[5][31] ), .QN(n4646) );
  DFFR_X1 \Mpath/regB/data_out_reg[7]  ( .D(n3805), .CK(CLK), .RN(n7817), .Q(
        \Mpath/out_regB[7] ), .QN(\Mpath/the_alu/N70 ) );
  DFFR_X2 \Mpath/regA/data_out_reg[9]  ( .D(n3851), .CK(CLK), .RN(n7782), .Q(
        \Mpath/out_regA[9] ), .QN(\Mpath/the_alu/N65 ) );
  DFFR_X2 \regfile/rx_28/data_out_reg[31]  ( .D(n3931), .CK(CLK), .RN(n7742), 
        .Q(\regfile/reg_out[28][31] ), .QN(n4870) );
  DFFR_X2 \regfile/rx_29/data_out_reg[31]  ( .D(n4141), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[29][31] ), .QN(n4838) );
  DFFR_X1 \Mpath/regB/data_out_reg[16]  ( .D(n3452), .CK(CLK), .RN(n7791), .Q(
        \Mpath/out_regB[16] ), .QN(\Mpath/the_alu/N52 ) );
  DFFS_X2 \Mcontrol/ir_dx/out_mem_command_reg[MW]  ( .D(n4413), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_sampled_dmem_command[MW] ), .QN(
        n3083) );
  DFFR_X2 \Mpath/regA/data_out_reg[19]  ( .D(n3336), .CK(CLK), .RN(n7731), .Q(
        \Mpath/out_regA[19] ), .QN(\Mpath/the_alu/N45 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[17]  ( .D(n3413), .CK(CLK), .RN(n7751), .Q(
        \Mpath/out_regB[17] ), .QN(\Mpath/the_alu/N50 ) );
  DFFR_X2 \Mpath/regB/data_out_reg[6]  ( .D(n3763), .CK(CLK), .RN(n7738), .Q(
        \Mpath/out_regB[6] ), .QN(\Mpath/the_alu/N72 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[15]  ( .D(n3491), .CK(CLK), .RN(n7790), .Q(
        \Mpath/out_regB[15] ), .QN(\Mpath/the_alu/N54 ) );
  DFFR_X1 \Mpath/regB/data_out_reg[13]  ( .D(n3652), .CK(CLK), .RN(n7752), .Q(
        \Mpath/out_regB[13] ), .QN(\Mpath/the_alu/N58 ) );
  DFFR_X2 \Mcontrol/ir_fd/data_out_reg[3]  ( .D(n4372), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [3]), .QN(n7287)
         );
  DFFR_X1 \Mcontrol/irfd/q_reg  ( .D(n4424), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(n7673), .QN(n6073) );
  DFFR_X2 \Mpath/regB/data_out_reg[12]  ( .D(n3613), .CK(CLK), .RN(n7773), .Q(
        \Mpath/out_regB[12] ), .QN(\Mpath/the_alu/N60 ) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[4]  ( .D(n4375), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [4]), .QN(n7352)
         );
  DFFR_X1 \Mpath/regA/data_out_reg[12]  ( .D(n3614), .CK(CLK), .RN(n7773), .Q(
        \Mpath/out_regA[12] ), .QN(\Mpath/the_alu/N59 ) );
  DFFS_X2 \Mcontrol/ir_dx/out_mul_command_reg[3]  ( .D(n4371), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_mul_command [3]), .QN(n3052) );
  DFFR_X1 \Mcontrol/ir_dx/out_alu_command_reg[OP][3]  ( .D(n4370), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][3] ), .QN(n3051) );
  NAND2_X2 syn1837 ( .A1(n7013), .A2(\Mcontrol/d_jump_type[3] ), .ZN(n6993) );
  NAND2_X2 syn1835 ( .A1(n7015), .A2(n7014), .ZN(n6994) );
  INV_X2 syn1831 ( .A(n6998), .ZN(n7010) );
  INV_X2 syn1829 ( .A(n7008), .ZN(n6999) );
  INV_X2 syn1824 ( .A(n7007), .ZN(n7001) );
  INV_X2 syn1030 ( .A(n7016), .ZN(n6397) );
  NAND3_X1 syn1029 ( .A1(net59736), .A2(net59612), .A3(net59757), .ZN(n7016)
         );
  INV_X2 syn973 ( .A(\Mcontrol/bvgen/N2 ), .ZN(n7015) );
  INV_X2 syn960 ( .A(net55826), .ZN(n7014) );
  INV_X2 syn952 ( .A(net55912), .ZN(n7013) );
  NOR2_X2 syn918 ( .A1(n7006), .A2(n7011), .ZN(n7000) );
  OAI21_X2 syn917 ( .B1(n6221), .B2(net59734), .A(n7012), .ZN(n7011) );
  NOR2_X2 syn912 ( .A1(\Mcontrol/Nextpc_decoding/N182 ), .A2(
        \Mcontrol/d_jump_type[2] ), .ZN(n6996) );
  NOR2_X2 syn910 ( .A1(\Mcontrol/d_jump_type[1] ), .A2(
        \Mcontrol/Nextpc_decoding/N173 ), .ZN(n6997) );
  OAI21_X2 syn907 ( .B1(n7003), .B2(n6046), .A(net57730), .ZN(n6990) );
  NOR2_X2 syn865 ( .A1(n1557), .A2(n7005), .ZN(n7008) );
  NOR2_X2 syn863 ( .A1(net59767), .A2(n7004), .ZN(n7007) );
  NOR2_X2 syn860 ( .A1(n1623), .A2(net59732), .ZN(n7006) );
  INV_X2 syn856 ( .A(jar_in[23]), .ZN(n7004) );
  INV_X2 syn853 ( .A(n1562), .ZN(net59734) );
  INV_X2 syn852 ( .A(n1563), .ZN(net59732) );
  INV_X2 syn835 ( .A(net56319), .ZN(n6991) );
  INV_X2 syn830 ( .A(n2492), .ZN(n7003) );
  NAND3_X1 \I_ADDR_OUTBUS[23]_inst  ( .A1(n6999), .A2(n7000), .A3(n7001), .ZN(
        n6998) );
  INV_X2 net58775 ( .A(n1623), .ZN(break_code[23]) );
  NAND2_X2 \Mcontrol/Nextpc_decoding/N178  ( .A1(n6996), .A2(n6997), .ZN(
        net59612) );
  NAND2_X2 net58683 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(n6995), .ZN(
        \Mcontrol/Nextpc_decoding/N182 ) );
  NAND2_X2 net58986 ( .A1(n6993), .A2(n6994), .ZN(n4393) );
  OR3_X4 net58736 ( .A1(n6990), .A2(n6991), .A3(n6992), .ZN(
        \Mcontrol/d_jump_type[3] ) );
  INV_X2 net58991 ( .A(n6046), .ZN(n6040) );
  DFFR_X2 \Mcontrol/ir_dx/out_alu_command_reg[OP][2]  ( .D(n4366), .CK(CLK), 
        .RN(\Mcontrol/int_reset ), .Q(\Alu_command[OP][2] ), .QN(n3049) );
  NAND2_X2 syn674 ( .A1(n6949), .A2(n6948), .ZN(n6933) );
  INV_X2 syn670 ( .A(n6934), .ZN(n6949) );
  INV_X2 syn668 ( .A(n6947), .ZN(n6935) );
  NAND2_X2 syn665 ( .A1(net58826), .A2(\Mcontrol/Nextpc_decoding/Bta [22]), 
        .ZN(n6948) );
  INV_X2 syn661 ( .A(n6946), .ZN(n6938) );
  INV_X2 syn652 ( .A(net59757), .ZN(n6932) );
  INV_X2 syn512 ( .A(n6234), .ZN(n6950) );
  INV_X2 syn451 ( .A(n6942), .ZN(n1562) );
  INV_X2 syn433 ( .A(\Mcontrol/Nextpc_decoding/N182 ), .ZN(n6931) );
  INV_X2 syn393 ( .A(\Mcontrol/Nextpc_decoding/N286 ), .ZN(n6927) );
  INV_X2 syn391 ( .A(\Mcontrol/Nextpc_decoding/N292 ), .ZN(n6926) );
  AOI21_X2 syn355 ( .B1(n1562), .B2(n6950), .A(n6945), .ZN(n6937) );
  NOR2_X2 syn351 ( .A1(\Mcontrol/d_jump_type[2] ), .A2(n6939), .ZN(n6930) );
  NAND2_X2 syn345 ( .A1(n6948), .A2(n6949), .ZN(net57039) );
  NOR2_X2 syn303 ( .A1(n1557), .A2(n6944), .ZN(n6947) );
  NOR2_X2 syn300 ( .A1(n6951), .A2(n6943), .ZN(n6946) );
  NOR2_X2 syn298 ( .A1(n374), .A2(n6941), .ZN(n6945) );
  INV_X2 syn297 ( .A(n6952), .ZN(n6944) );
  INV_X2 syn293 ( .A(jar_in[22]), .ZN(n6943) );
  NAND2_X2 syn292 ( .A1(n6932), .A2(n6940), .ZN(n6942) );
  NAND4_X1 \I_ADDR_OUTBUS[22]_inst  ( .A1(n6935), .A2(n6936), .A3(n6937), .A4(
        n6938), .ZN(n6934) );
  NAND2_X2 net60658 ( .A1(n6933), .A2(n372), .ZN(net56784) );
  INV_X2 net60469 ( .A(n374), .ZN(break_code[22]) );
  INV_X2 net60510 ( .A(net55921), .ZN(n1561) );
  NAND3_X1 \Mcontrol/Nextpc_decoding/N185  ( .A1(n6929), .A2(n6930), .A3(n6931), .ZN(net59757) );
  NAND2_X2 net60408 ( .A1(n6928), .A2(n6953), .ZN(
        \Mcontrol/Nextpc_decoding/N299 ) );
  NAND2_X2 net60404 ( .A1(n6927), .A2(n6953), .ZN(
        \Mcontrol/Nextpc_decoding/N287 ) );
  NAND2_X2 net60406 ( .A1(n6926), .A2(n6953), .ZN(
        \Mcontrol/Nextpc_decoding/N293 ) );
  OAI21_X1 U5018 ( .B1(net57038), .B2(net57810), .A(n6100), .ZN(n6079) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2062  ( .A1(\Mcontrol/d_instr[0] ), 
        .A2(\Mcontrol/Operation_decoding32/N1886 ), .ZN(
        \Mcontrol/Operation_decoding32/N1887 ) );
  AND2_X2 \Mcontrol/Operation_decoding32/C2078  ( .A1(\Mcontrol/d_instr[0] ), 
        .A2(\Mcontrol/Operation_decoding32/N1897 ), .ZN(
        \Mcontrol/Operation_decoding32/N1898 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2092  ( .A1(\Mcontrol/d_instr[0] ), 
        .A2(\Mcontrol/Operation_decoding32/N1911 ), .ZN(
        \Mcontrol/Operation_decoding32/N1912 ) );
  INV_X1 U5026 ( .A(n5520), .ZN(\Mcontrol/d_instr[0] ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2086  ( .A1(
        \Mcontrol/Operation_decoding32/N1901 ), .A2(
        \Mcontrol/Operation_decoding32/N1905 ), .ZN(
        \Mcontrol/Operation_decoding32/N1906 ) );
  INV_X2 \Mcontrol/Operation_decoding32/I_8  ( .A(\Mcontrol/d_instr[0] ), .ZN(
        \Mcontrol/Operation_decoding32/N1901 ) );
  OR2_X2 \Mcontrol/Operation_decoding32/C2094  ( .A1(\Mcontrol/d_instr[6] ), 
        .A2(\Mcontrol/d_instr [7]), .ZN(\Mcontrol/Operation_decoding32/N1914 )
         );
  AOI221_X1 U4112 ( .B1(\Mcontrol/d_instr[6] ), .B2(n333), .C1(n6227), .C2(
        n331), .A(n330), .ZN(n374) );
  DFFS_X1 \Scc_coproc/dec_eword_reg/data_out_reg[4]  ( .D(n3896), .CK(CLK), 
        .SN(n7822), .Q(\Scc_coproc/din_exc_word[4] ), .QN(n1062) );
  DFFR_X1 \Mpath/regA/data_out_reg[8]  ( .D(n3913), .CK(CLK), .RN(n7726), .Q(
        n1834), .QN(n7184) );
  DFFS_X1 \Scc_coproc/dec_eword_reg/data_out_reg[5]  ( .D(n3897), .CK(CLK), 
        .SN(n7824), .Q(\Scc_coproc/din_exc_word[5] ), .QN(n1064) );
  DFFS_X1 \Scc_coproc/dec_eword_reg/data_out_reg[0]  ( .D(n4427), .CK(CLK), 
        .SN(n7822), .Q(\Scc_coproc/din_exc_word[0] ), .QN(n1552) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[4]  ( .D(n3696), .CK(CLK), .SN(
        n6550), .Q(\Mcontrol/f_currpc[4] ) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_e/data_out_reg[2]  ( .D(n4502), .CK(CLK), 
        .SN(n7849), .QN(n1682) );
  DFFS_X1 \Scc_coproc/Delay_ref_reg_e/data_out_reg[1]  ( .D(n4503), .CK(CLK), 
        .SN(n7850), .QN(n1683) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[4]  ( .D(n3892), .CK(CLK), .SN(
        n6550), .Q(\Scc_coproc/ein_exc_word[4] ), .QN(n1054) );
  DFFS_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[8]  ( .D(n3688), .CK(CLK), 
        .SN(n7786), .Q(\Mcontrol/bvgen/x_curr_pc [8]), .QN(n823) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[15]  ( .D(n3492), .CK(CLK), 
        .SN(n6550), .QN(n625) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[7]  ( .D(n3806), .CK(CLK), 
        .SN(n6550), .QN(n970) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[6]  ( .D(n3764), .CK(CLK), 
        .SN(n7845), .QN(n931) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[5]  ( .D(n3722), .CK(CLK), 
        .SN(n6550), .QN(n887) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[3]  ( .D(n4435), .CK(CLK), 
        .SN(n7808), .QN(n1582) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[4]  ( .D(n4440), .CK(CLK), 
        .SN(n6550), .QN(n1592) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[2]  ( .D(n4430), .CK(CLK), 
        .SN(n7787), .QN(n1575) );
  DFFS_X1 \Scc_coproc/X_status_reg/data_out_reg[14]  ( .D(n4449), .CK(CLK), 
        .SN(n7738), .Q(\Scc_coproc/x_status[14] ), .QN(n1603) );
  DFFS_X1 \Mcontrol/ir_dx/out_mem_command_reg[MB]  ( .D(n4408), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(n1519) );
  DFFS_X1 \Mcontrol/ir_dx/out_mem_command_reg[MR]  ( .D(n4412), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(n1530) );
  DFFS_X1 \Mcontrol/ir_dx/out_mem_command_reg[SIGN]  ( .D(n4415), .CK(CLK), 
        .SN(\Mcontrol/int_reset ), .Q(\Mcontrol/x_sampled_dmem_command[SIGN] )
         );
  DFFS_X1 \Mcontrol/ir_dx/out_mem_command_reg[MH]  ( .D(n4410), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(n1526) );
  DFFS_X1 \Mcontrol/ir_dx/out_alu_command_reg[HRDWIT]  ( .D(n4406), .CK(CLK), 
        .SN(\Mcontrol/int_reset ), .QN(n1515) );
  DFFS_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[8]  ( .D(n3687), .CK(CLK), 
        .SN(n7789), .QN(n820) );
  DFFS_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[2]  ( .D(n3705), .CK(CLK), 
        .SN(n7785), .QN(n853) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[0]  ( .D(n4426), .CK(CLK), .SN(
        n7818), .Q(\Scc_coproc/ein_exc_word[0] ), .QN(n1551) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[3]  ( .D(n3893), .CK(CLK), .SN(
        n6550), .Q(\Scc_coproc/ein_exc_word[3] ), .QN(n1057) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[2]  ( .D(n3894), .CK(CLK), .SN(
        n6550), .Q(\Scc_coproc/ein_exc_word[2] ), .QN(n1058) );
  DFFS_X1 \Scc_coproc/x_eword_reg/data_out_reg[1]  ( .D(n3891), .CK(CLK), .SN(
        n6550), .Q(\Scc_coproc/ein_exc_word[1] ), .QN(n1052) );
  DFFS_X1 \Scc_coproc/CAUSE_REG/data_out_reg[4]  ( .D(n4444), .CK(CLK), .SN(
        n7819), .Q(\Scc_coproc/cause[4] ) );
  DFFS_X1 \Mcontrol/ir_dx/out_rf_we_reg  ( .D(n4423), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_sampled_dwe ), .QN(n1546) );
  DFFS_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[8]  ( .D(n3689), .CK(CLK), 
        .SN(n7825), .Q(\Mcontrol/bvgen/d_curr_pc[8] ), .QN(n824) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[11]  ( .D(n3573), .CK(CLK), 
        .SN(n7851), .Q(\Mcontrol/f_currpc[11] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[9]  ( .D(n3846), .CK(CLK), .SN(
        n7848), .Q(\Mcontrol/f_currpc[9] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[2]  ( .D(n3708), .CK(CLK), .SN(
        n7847), .Q(\Mcontrol/f_currpc[2] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[7]  ( .D(n3804), .CK(CLK), .SN(
        n7846), .Q(\Mcontrol/f_currpc[7] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[6]  ( .D(n3762), .CK(CLK), .SN(
        n7814), .Q(\Mcontrol/f_currpc[6] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[3]  ( .D(n3702), .CK(CLK), .SN(
        n7742), .Q(\Mcontrol/f_currpc[3] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[5]  ( .D(n3719), .CK(CLK), .SN(
        n7788), .Q(\Mcontrol/f_currpc[5] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[10]  ( .D(n4490), .CK(CLK), 
        .SN(n6550), .Q(\Mcontrol/f_currpc[10] ) );
  DFFS_X1 \Mcontrol/Program_counter/out_pc_reg[8]  ( .D(n3690), .CK(CLK), .SN(
        n7816), .Q(\Mcontrol/f_currpc[8] ) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[13]  ( .D(n3649), .CK(CLK), 
        .RN(n7777), .Q(\Mcontrol/bvgen/x_curr_pc [13]), .QN(n785) );
  DFFR_X1 \Scc_coproc/X_status_reg/data_out_reg[9]  ( .D(n3848), .CK(CLK), 
        .RN(n6550), .QN(n1009) );
  DFFR_X1 \Scc_coproc/X_status_reg/data_out_reg[8]  ( .D(n4445), .CK(CLK), 
        .RN(n7735), .QN(n1597) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[20]  ( .D(n3293), .CK(CLK), 
        .RN(n7766), .Q(\Mcontrol/bvgen/x_curr_pc [20]), .QN(n441) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[19]  ( .D(n3332), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [19]), .QN(n476) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[18]  ( .D(n3371), .CK(CLK), 
        .RN(n7731), .Q(\Mcontrol/bvgen/x_curr_pc [18]), .QN(n511) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[17]  ( .D(n3410), .CK(CLK), 
        .RN(n7767), .Q(\Mcontrol/bvgen/x_curr_pc [17]), .QN(n546) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[16]  ( .D(n3449), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [16]), .QN(n581) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[15]  ( .D(n3488), .CK(CLK), 
        .RN(n7723), .Q(\Mcontrol/bvgen/x_curr_pc [15]), .QN(n617) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[14]  ( .D(n3530), .CK(CLK), 
        .RN(n7768), .Q(\Mcontrol/bvgen/x_curr_pc [14]), .QN(n664) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[12]  ( .D(n3610), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [12]), .QN(n747) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[11]  ( .D(n3571), .CK(CLK), 
        .RN(n7729), .Q(\Mcontrol/bvgen/x_curr_pc [11]), .QN(n709) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[10]  ( .D(n3899), .CK(CLK), 
        .RN(n7769), .Q(\Mcontrol/bvgen/x_curr_pc [10]), .QN(n1065) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[9]  ( .D(n3844), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [9]), .QN(n1001) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[7]  ( .D(n3802), .CK(CLK), 
        .RN(n7824), .Q(\Mcontrol/bvgen/x_curr_pc [7]), .QN(n962) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[6]  ( .D(n3760), .CK(CLK), 
        .RN(n7771), .Q(\Mcontrol/bvgen/x_curr_pc [6]), .QN(n923) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[5]  ( .D(n3717), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [5]), .QN(n875) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[4]  ( .D(n3694), .CK(CLK), 
        .RN(n7842), .Q(\Mcontrol/bvgen/x_curr_pc [4]), .QN(n834) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[2]  ( .D(n3706), .CK(CLK), 
        .RN(n7796), .Q(\Mcontrol/bvgen/x_curr_pc [2]), .QN(n856) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[1]  ( .D(n3712), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [1]), .QN(n867) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[0]  ( .D(n3886), .CK(CLK), 
        .RN(n7826), .Q(\Mcontrol/bvgen/x_curr_pc [0]), .QN(n1039) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[23]  ( .D(n3902), .CK(CLK), 
        .RN(n7798), .Q(\Mcontrol/bvgen/x_curr_pc [23]), .QN(n1068) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[3]  ( .D(n3700), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [3]), .QN(n845) );
  DFFR_X1 \Mcontrol/ir_xm/out_rd1_reg[0]  ( .D(n4348), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/m_sampled_xrd[0] ), .QN(n1412) );
  DFFR_X1 \Mpath/JAR/data_out_reg[0]  ( .D(n4488), .CK(CLK), .RN(n7829), .Q(
        \Mpath/out_jar[0] ), .QN(n1652) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[22]  ( .D(n3215), .CK(CLK), 
        .RN(n7799), .Q(\Mcontrol/bvgen/x_curr_pc [22]), .QN(n363) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg2/data_out_reg[21]  ( .D(n3254), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/x_curr_pc [21]), .QN(n406) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[23]  ( .D(n3901), .CK(CLK), 
        .RN(n7828), .QN(n1047) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[21]  ( .D(n3253), .CK(CLK), 
        .RN(n7801), .QN(n404) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[20]  ( .D(n3292), .CK(CLK), 
        .RN(n6550), .QN(n439) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[19]  ( .D(n3331), .CK(CLK), 
        .RN(n7827), .QN(n474) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[18]  ( .D(n3370), .CK(CLK), 
        .RN(n7790), .QN(n509) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[17]  ( .D(n3409), .CK(CLK), 
        .RN(n6550), .QN(n544) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[16]  ( .D(n3448), .CK(CLK), 
        .RN(n7832), .QN(n579) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[15]  ( .D(n3487), .CK(CLK), 
        .RN(n7794), .QN(n614) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[14]  ( .D(n3529), .CK(CLK), 
        .RN(n6550), .QN(n661) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[13]  ( .D(n3648), .CK(CLK), 
        .RN(n7831), .QN(n782) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[12]  ( .D(n3609), .CK(CLK), 
        .RN(n7795), .QN(n744) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[11]  ( .D(n3570), .CK(CLK), 
        .RN(n6550), .QN(n706) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[10]  ( .D(n3898), .CK(CLK), 
        .RN(n7830), .QN(n676) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[9]  ( .D(n3843), .CK(CLK), 
        .RN(n7784), .QN(n998) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[7]  ( .D(n3801), .CK(CLK), 
        .RN(n6550), .QN(n959) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[6]  ( .D(n3759), .CK(CLK), 
        .RN(n7835), .QN(n920) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[5]  ( .D(n3716), .CK(CLK), 
        .RN(n7785), .QN(n872) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[4]  ( .D(n3693), .CK(CLK), 
        .RN(n6550), .QN(n831) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[3]  ( .D(n3699), .CK(CLK), 
        .RN(n7834), .QN(n842) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[1]  ( .D(n3711), .CK(CLK), 
        .RN(n7786), .QN(n864) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[0]  ( .D(n3885), .CK(CLK), 
        .RN(n6550), .QN(n1041) );
  DFFR_X1 \Scc_coproc/x_basevalue_reg/data_out_reg[22]  ( .D(n3214), .CK(CLK), 
        .RN(n7833), .QN(n358) );
  DFFR_X1 \Mcontrol/ir_dx/out_rd1_reg[3]  ( .D(n4355), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_rd[3] ), .QN(n1424) );
  DFFR_X1 \Mcontrol/ir_dx/out_rd1_reg[2]  ( .D(n4353), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_rd[2] ), .QN(n1421) );
  DFFR_X1 \Mcontrol/ir_dx/out_rd1_reg[1]  ( .D(n4351), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_rd[1] ), .QN(n1419) );
  DFFR_X1 \Mcontrol/ir_dx/out_rd1_reg[0]  ( .D(n4349), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_rd[0] ), .QN(n1411) );
  DFFR_X1 \Mcontrol/ir_dx/out_rd1_reg[4]  ( .D(n4357), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/x_rd[4] ), .QN(n1426) );
  DFFR_X1 \Mcontrol/bvgen/jtype_reg1/data_out_reg[0]  ( .D(n3904), .CK(CLK), 
        .RN(n7787), .Q(\Mcontrol/bvgen/x_jump_type[0] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[31]  ( .D(n3108), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[31] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[30]  ( .D(n3109), .CK(CLK), 
        .RN(n7838), .Q(\Mpath/the_memhandle/smdr_out[30] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[29]  ( .D(n3110), .CK(CLK), 
        .RN(n7788), .Q(\Mpath/the_memhandle/smdr_out[29] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[28]  ( .D(n3111), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[28] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[27]  ( .D(n3112), .CK(CLK), 
        .RN(n7837), .Q(\Mpath/the_memhandle/smdr_out[27] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[26]  ( .D(n3113), .CK(CLK), 
        .RN(n7789), .Q(\Mpath/the_memhandle/smdr_out[26] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[25]  ( .D(n3114), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[25] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[24]  ( .D(n3115), .CK(CLK), 
        .RN(n7836), .Q(\Mpath/the_memhandle/smdr_out[24] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[23]  ( .D(n3116), .CK(CLK), 
        .RN(n7814), .Q(\Mpath/the_memhandle/smdr_out[23] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[22]  ( .D(n3117), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[22] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[21]  ( .D(n3118), .CK(CLK), 
        .RN(n7841), .Q(\Mpath/the_memhandle/smdr_out[21] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[20]  ( .D(n3119), .CK(CLK), 
        .RN(n7816), .Q(\Mpath/the_memhandle/smdr_out[20] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[19]  ( .D(n3120), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[19] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[18]  ( .D(n3121), .CK(CLK), 
        .RN(n7840), .Q(\Mpath/the_memhandle/smdr_out[18] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[17]  ( .D(n3122), .CK(CLK), 
        .RN(n7818), .Q(\Mpath/the_memhandle/smdr_out[17] ) );
  DFFR_X1 \Mpath/the_memhandle/SMDR/data_out_reg[16]  ( .D(n3123), .CK(CLK), 
        .RN(n6550), .Q(\Mpath/the_memhandle/smdr_out[16] ) );
  DFFR_X1 \Scc_coproc/CAUSE_REG/data_out_reg[5]  ( .D(n3884), .CK(CLK), .RN(
        n7839), .Q(\Scc_coproc/cause[5] ) );
  DFFR_X1 \regfile/rx_1/data_out_reg[29]  ( .D(n4340), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[1][29] ), .QN(n1399) );
  DFFR_X1 \regfile/rx_1/data_out_reg[27]  ( .D(n4342), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][27] ), .QN(n1401) );
  DFFR_X1 \regfile/rx_1/data_out_reg[24]  ( .D(n3191), .CK(CLK), .RN(n7843), 
        .Q(\regfile/reg_out[1][24] ), .QN(n344) );
  DFFR_X1 \regfile/rx_1/data_out_reg[23]  ( .D(n4344), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][23] ), .QN(n1403) );
  DFFR_X1 \regfile/rx_1/data_out_reg[18]  ( .D(n3386), .CK(CLK), .RN(n7775), 
        .Q(\regfile/reg_out[1][18] ), .QN(n529) );
  DFFR_X1 \regfile/rx_1/data_out_reg[16]  ( .D(n3464), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[1][16] ), .QN(n599) );
  DFFR_X1 \regfile/rx_1/data_out_reg[6]  ( .D(n3778), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][6] ), .QN(n942) );
  DFFR_X1 \regfile/rx_1/data_out_reg[4]  ( .D(n4335), .CK(CLK), .RN(n7774), 
        .Q(\regfile/reg_out[1][4] ), .QN(n1383) );
  DFFR_X1 \regfile/rx_1/data_out_reg[10]  ( .D(n3547), .CK(CLK), .RN(n7758), 
        .Q(\regfile/reg_out[1][10] ), .QN(n689) );
  DFFR_X1 \regfile/rx_1/data_out_reg[9]  ( .D(n3862), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][9] ), .QN(n1020) );
  DFFR_X1 \regfile/rx_2/data_out_reg[23]  ( .D(n4120), .CK(CLK), .RN(n7772), 
        .Q(\regfile/reg_out[2][23] ), .QN(n1233) );
  DFFR_X1 \regfile/rx_2/data_out_reg[30]  ( .D(n4114), .CK(CLK), .RN(n7750), 
        .Q(\regfile/reg_out[2][30] ), .QN(n1227) );
  DFFR_X1 \regfile/rx_2/data_out_reg[29]  ( .D(n4116), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][29] ), .QN(n1229) );
  DFFR_X1 \regfile/rx_2/data_out_reg[28]  ( .D(n4117), .CK(CLK), .RN(n7783), 
        .Q(\regfile/reg_out[2][28] ), .QN(n1230) );
  DFFR_X1 \regfile/rx_2/data_out_reg[27]  ( .D(n4118), .CK(CLK), .RN(n7779), 
        .Q(\regfile/reg_out[2][27] ), .QN(n1231) );
  DFFR_X1 \regfile/rx_2/data_out_reg[31]  ( .D(n4113), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][31] ), .QN(n1226) );
  DFFR_X1 \regfile/rx_2/data_out_reg[26]  ( .D(n4119), .CK(CLK), .RN(n7781), 
        .Q(\regfile/reg_out[2][26] ), .QN(n1232) );
  DFFR_X1 \regfile/rx_2/data_out_reg[25]  ( .D(n3168), .CK(CLK), .RN(n7776), 
        .Q(\regfile/reg_out[2][25] ), .QN(n293) );
  DFFR_X1 \regfile/rx_2/data_out_reg[24]  ( .D(n3202), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][24] ), .QN(n349) );
  DFFR_X1 \regfile/rx_2/data_out_reg[22]  ( .D(n3241), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[2][22] ), .QN(n393) );
  DFFR_X1 \regfile/rx_2/data_out_reg[21]  ( .D(n3280), .CK(CLK), .RN(n7797), 
        .Q(\regfile/reg_out[2][21] ), .QN(n429) );
  DFFR_X1 \regfile/rx_2/data_out_reg[20]  ( .D(n3319), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][20] ), .QN(n464) );
  DFFR_X1 \regfile/rx_2/data_out_reg[19]  ( .D(n3358), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[2][19] ), .QN(n499) );
  DFFR_X1 \regfile/rx_2/data_out_reg[18]  ( .D(n3397), .CK(CLK), .RN(n7791), 
        .Q(\regfile/reg_out[2][18] ), .QN(n534) );
  DFFR_X1 \regfile/rx_2/data_out_reg[17]  ( .D(n3436), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][17] ), .QN(n569) );
  DFFR_X1 \regfile/rx_2/data_out_reg[16]  ( .D(n3475), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[2][16] ), .QN(n604) );
  DFFR_X1 \regfile/rx_2/data_out_reg[7]  ( .D(n3831), .CK(CLK), .RN(n7793), 
        .Q(\regfile/reg_out[2][7] ), .QN(n986) );
  DFFR_X1 \regfile/rx_2/data_out_reg[1]  ( .D(n4121), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][1] ), .QN(n1234) );
  DFFR_X1 \regfile/rx_2/data_out_reg[0]  ( .D(n4123), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[2][0] ), .QN(n1236) );
  DFFR_X1 \regfile/rx_2/data_out_reg[14]  ( .D(n4122), .CK(CLK), .RN(n7815), 
        .Q(\regfile/reg_out[2][14] ), .QN(n1235) );
  DFFR_X1 \regfile/rx_2/data_out_reg[13]  ( .D(n3675), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][13] ), .QN(n808) );
  DFFR_X1 \regfile/rx_2/data_out_reg[12]  ( .D(n3636), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[2][12] ), .QN(n770) );
  DFFR_X1 \regfile/rx_2/data_out_reg[11]  ( .D(n3597), .CK(CLK), .RN(n7817), 
        .Q(\regfile/reg_out[2][11] ), .QN(n732) );
  DFFR_X1 \regfile/rx_2/data_out_reg[10]  ( .D(n3558), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][10] ), .QN(n694) );
  DFFR_X1 \regfile/rx_2/data_out_reg[6]  ( .D(n3789), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[2][6] ), .QN(n947) );
  DFFR_X1 \regfile/rx_2/data_out_reg[5]  ( .D(n3747), .CK(CLK), .RN(n7809), 
        .Q(\regfile/reg_out[2][5] ), .QN(n903) );
  DFFR_X1 \regfile/rx_2/data_out_reg[4]  ( .D(n4111), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][4] ), .QN(n1224) );
  DFFR_X1 \regfile/rx_2/data_out_reg[3]  ( .D(n4112), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[2][3] ), .QN(n1225) );
  DFFR_X1 \regfile/rx_2/data_out_reg[2]  ( .D(n4115), .CK(CLK), .RN(n7812), 
        .Q(\regfile/reg_out[2][2] ), .QN(n1228) );
  DFFR_X1 \regfile/rx_2/data_out_reg[15]  ( .D(n3517), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[2][15] ), .QN(n645) );
  DFFR_X1 \regfile/rx_2/data_out_reg[9]  ( .D(n3873), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[2][9] ), .QN(n1025) );
  DFFR_X1 \regfile/rx_2/data_out_reg[8]  ( .D(n4110), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[2][8] ), .QN(n1223) );
  DFFR_X1 \regfile/rx_1/data_out_reg[31]  ( .D(n4337), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][31] ), .QN(n1389) );
  DFFR_X1 \regfile/rx_1/data_out_reg[30]  ( .D(n4338), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[1][30] ), .QN(n1391) );
  DFFR_X1 \regfile/rx_1/data_out_reg[28]  ( .D(n4341), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[1][28] ), .QN(n1400) );
  DFFR_X1 \regfile/rx_1/data_out_reg[26]  ( .D(n4343), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][26] ), .QN(n1402) );
  DFFR_X1 \regfile/rx_1/data_out_reg[25]  ( .D(n3157), .CK(CLK), .RN(n7734), 
        .Q(\regfile/reg_out[1][25] ), .QN(n266) );
  DFFR_X1 \regfile/rx_1/data_out_reg[22]  ( .D(n3230), .CK(CLK), .RN(n7844), 
        .Q(\regfile/reg_out[1][22] ), .QN(n388) );
  DFFR_X1 \regfile/rx_1/data_out_reg[21]  ( .D(n3269), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][21] ), .QN(n424) );
  DFFR_X1 \regfile/rx_1/data_out_reg[20]  ( .D(n3308), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[1][20] ), .QN(n459) );
  DFFR_X1 \regfile/rx_1/data_out_reg[19]  ( .D(n3347), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[1][19] ), .QN(n494) );
  DFFR_X1 \regfile/rx_1/data_out_reg[17]  ( .D(n3425), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][17] ), .QN(n564) );
  DFFR_X1 \regfile/rx_1/data_out_reg[5]  ( .D(n3736), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[1][5] ), .QN(n898) );
  DFFR_X1 \regfile/rx_1/data_out_reg[3]  ( .D(n4336), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[1][3] ), .QN(n1386) );
  DFFR_X1 \regfile/rx_1/data_out_reg[2]  ( .D(n4339), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][2] ), .QN(n1392) );
  DFFR_X1 \regfile/rx_1/data_out_reg[15]  ( .D(n3506), .CK(CLK), .RN(n7730), 
        .Q(\regfile/reg_out[1][15] ), .QN(n640) );
  DFFR_X1 \regfile/rx_1/data_out_reg[14]  ( .D(n4346), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[1][14] ), .QN(n1407) );
  DFFR_X1 \regfile/rx_1/data_out_reg[13]  ( .D(n3664), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][13] ), .QN(n803) );
  DFFR_X1 \regfile/rx_1/data_out_reg[12]  ( .D(n3625), .CK(CLK), .RN(n7740), 
        .Q(\regfile/reg_out[1][12] ), .QN(n765) );
  DFFR_X1 \regfile/rx_1/data_out_reg[11]  ( .D(n3586), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[1][11] ), .QN(n727) );
  DFFR_X1 \regfile/rx_1/data_out_reg[8]  ( .D(n4334), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][8] ), .QN(n1380) );
  DFFR_X1 \regfile/rx_1/data_out_reg[7]  ( .D(n3820), .CK(CLK), .RN(n7737), 
        .Q(\regfile/reg_out[1][7] ), .QN(n981) );
  DFFR_X1 \regfile/rx_1/data_out_reg[1]  ( .D(n4345), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[1][1] ), .QN(n1405) );
  DFFR_X1 \regfile/rx_1/data_out_reg[0]  ( .D(n4347), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[1][0] ), .QN(n1410) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[1]  ( .D(n3713), .CK(CLK), 
        .RN(n7736), .Q(\Mcontrol/bvgen/d_curr_pc[1] ), .QN(n868) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[0]  ( .D(n3887), .CK(CLK), 
        .RN(n7721), .Q(\Mcontrol/bvgen/d_curr_pc[0] ), .QN(n1040) );
  DFFR_X1 \regfile/rx_22/data_out_reg[23]  ( .D(n3980), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][23] ), .QN(n1133) );
  DFFR_X1 \regfile/rx_22/data_out_reg[30]  ( .D(n3974), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[22][30] ), .QN(n1127) );
  DFFR_X1 \regfile/rx_22/data_out_reg[29]  ( .D(n3976), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[22][29] ), .QN(n1129) );
  DFFR_X1 \regfile/rx_22/data_out_reg[28]  ( .D(n3977), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][28] ), .QN(n1130) );
  DFFR_X1 \regfile/rx_22/data_out_reg[27]  ( .D(n3978), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[22][27] ), .QN(n1131) );
  DFFR_X1 \regfile/rx_22/data_out_reg[31]  ( .D(n3973), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[22][31] ), .QN(n1126) );
  DFFR_X1 \regfile/rx_22/data_out_reg[26]  ( .D(n3979), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][26] ), .QN(n1132) );
  DFFR_X1 \regfile/rx_22/data_out_reg[25]  ( .D(n3160), .CK(CLK), .RN(n7722), 
        .Q(\regfile/reg_out[22][25] ), .QN(n273) );
  DFFR_X1 \regfile/rx_22/data_out_reg[24]  ( .D(n3194), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[22][24] ), .QN(n345) );
  DFFR_X1 \regfile/rx_22/data_out_reg[22]  ( .D(n3233), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][22] ), .QN(n389) );
  DFFR_X1 \regfile/rx_22/data_out_reg[21]  ( .D(n3272), .CK(CLK), .RN(n7721), 
        .Q(\regfile/reg_out[22][21] ), .QN(n425) );
  DFFR_X1 \regfile/rx_22/data_out_reg[20]  ( .D(n3311), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[22][20] ), .QN(n460) );
  DFFR_X1 \regfile/rx_22/data_out_reg[19]  ( .D(n3350), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][19] ), .QN(n495) );
  DFFR_X1 \regfile/rx_22/data_out_reg[18]  ( .D(n3389), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[22][18] ), .QN(n530) );
  DFFR_X1 \regfile/rx_22/data_out_reg[17]  ( .D(n3428), .CK(CLK), .RN(n7737), 
        .Q(\regfile/reg_out[22][17] ), .QN(n565) );
  DFFR_X1 \regfile/rx_22/data_out_reg[16]  ( .D(n3467), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][16] ), .QN(n600) );
  DFFR_X1 \regfile/rx_22/data_out_reg[7]  ( .D(n3823), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[22][7] ), .QN(n982) );
  DFFR_X1 \regfile/rx_22/data_out_reg[1]  ( .D(n3981), .CK(CLK), .RN(n7740), 
        .Q(\regfile/reg_out[22][1] ), .QN(n1134) );
  DFFR_X1 \regfile/rx_22/data_out_reg[0]  ( .D(n3983), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][0] ), .QN(n1136) );
  DFFR_X1 \regfile/rx_22/data_out_reg[14]  ( .D(n3982), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[22][14] ), .QN(n1135) );
  DFFR_X1 \regfile/rx_22/data_out_reg[13]  ( .D(n3667), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[22][13] ), .QN(n804) );
  DFFR_X1 \regfile/rx_22/data_out_reg[12]  ( .D(n3628), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][12] ), .QN(n766) );
  DFFR_X1 \regfile/rx_22/data_out_reg[11]  ( .D(n3589), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[22][11] ), .QN(n728) );
  DFFR_X1 \regfile/rx_22/data_out_reg[10]  ( .D(n3550), .CK(CLK), .RN(n7733), 
        .Q(\regfile/reg_out[22][10] ), .QN(n690) );
  DFFR_X1 \regfile/rx_22/data_out_reg[6]  ( .D(n3781), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][6] ), .QN(n943) );
  DFFR_X1 \regfile/rx_22/data_out_reg[5]  ( .D(n3739), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[22][5] ), .QN(n899) );
  DFFR_X1 \regfile/rx_22/data_out_reg[4]  ( .D(n3971), .CK(CLK), .RN(n7734), 
        .Q(\regfile/reg_out[22][4] ), .QN(n1124) );
  DFFR_X1 \regfile/rx_22/data_out_reg[3]  ( .D(n3972), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][3] ), .QN(n1125) );
  DFFR_X1 \regfile/rx_22/data_out_reg[2]  ( .D(n3975), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[22][2] ), .QN(n1128) );
  DFFR_X1 \regfile/rx_22/data_out_reg[15]  ( .D(n3509), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[22][15] ), .QN(n641) );
  DFFR_X1 \regfile/rx_22/data_out_reg[9]  ( .D(n3865), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[22][9] ), .QN(n1021) );
  DFFR_X1 \regfile/rx_22/data_out_reg[8]  ( .D(n3970), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[22][8] ), .QN(n1123) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[23]  ( .D(n3903), .CK(CLK), 
        .RN(n7764), .Q(\Mcontrol/bvgen/d_curr_pc[23] ), .QN(n1069) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[22]  ( .D(n3216), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[22] ), .QN(n365) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[21]  ( .D(n3255), .CK(CLK), 
        .RN(n7716), .Q(\Mcontrol/bvgen/d_curr_pc[21] ), .QN(n407) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[20]  ( .D(n3294), .CK(CLK), 
        .RN(n7765), .Q(\Mcontrol/bvgen/d_curr_pc[20] ), .QN(n442) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[19]  ( .D(n3333), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[19] ), .QN(n477) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[18]  ( .D(n3372), .CK(CLK), 
        .RN(n7821), .Q(\Mcontrol/bvgen/d_curr_pc[18] ), .QN(n512) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[17]  ( .D(n3411), .CK(CLK), 
        .RN(n7757), .Q(\Mcontrol/bvgen/d_curr_pc[17] ), .QN(n547) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[16]  ( .D(n3450), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[16] ), .QN(n582) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[15]  ( .D(n3489), .CK(CLK), 
        .RN(n7845), .Q(\Mcontrol/bvgen/d_curr_pc[15] ), .QN(n618) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[14]  ( .D(n3531), .CK(CLK), 
        .RN(n7749), .Q(\Mcontrol/bvgen/d_curr_pc[14] ), .QN(n665) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[13]  ( .D(n3650), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[13] ), .QN(n786) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[12]  ( .D(n3611), .CK(CLK), 
        .RN(n7744), .Q(\Mcontrol/bvgen/d_curr_pc[12] ), .QN(n748) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[11]  ( .D(n3572), .CK(CLK), 
        .RN(n7778), .Q(\Mcontrol/bvgen/d_curr_pc[11] ), .QN(n710) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[10]  ( .D(n3900), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[10] ), .QN(n1066) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[9]  ( .D(n3845), .CK(CLK), 
        .RN(n7844), .Q(\Mcontrol/bvgen/d_curr_pc[9] ), .QN(n1002) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[7]  ( .D(n3803), .CK(CLK), 
        .RN(n7780), .Q(\Mcontrol/bvgen/d_curr_pc[7] ), .QN(n963) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[6]  ( .D(n3761), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[6] ), .QN(n924) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[5]  ( .D(n3718), .CK(CLK), 
        .RN(n7822), .Q(\Mcontrol/bvgen/d_curr_pc[5] ), .QN(n876) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[4]  ( .D(n3695), .CK(CLK), 
        .RN(n7781), .Q(\Mcontrol/bvgen/d_curr_pc[4] ), .QN(n835) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[3]  ( .D(n3701), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/bvgen/d_curr_pc[3] ), .QN(n846) );
  DFFR_X1 \Mcontrol/bvgen/pcbv_reg1/data_out_reg[2]  ( .D(n3707), .CK(CLK), 
        .RN(n7829), .Q(\Mcontrol/bvgen/d_curr_pc[2] ), .QN(n857) );
  DFFR_X1 \regfile/rx_10/data_out_reg[23]  ( .D(n4064), .CK(CLK), .RN(n7783), 
        .QN(n1189) );
  DFFR_X1 \regfile/rx_10/data_out_reg[30]  ( .D(n4058), .CK(CLK), .RN(n6550), 
        .QN(n1183) );
  DFFR_X1 \regfile/rx_10/data_out_reg[29]  ( .D(n4060), .CK(CLK), .RN(n7828), 
        .QN(n1185) );
  DFFR_X1 \regfile/rx_10/data_out_reg[28]  ( .D(n4061), .CK(CLK), .RN(n7772), 
        .QN(n1186) );
  DFFR_X1 \regfile/rx_10/data_out_reg[27]  ( .D(n4062), .CK(CLK), .RN(n6550), 
        .QN(n1187) );
  DFFR_X1 \regfile/rx_10/data_out_reg[31]  ( .D(n4057), .CK(CLK), .RN(n7827), 
        .QN(n1182) );
  DFFR_X1 \regfile/rx_10/data_out_reg[26]  ( .D(n4063), .CK(CLK), .RN(n7774), 
        .QN(n1188) );
  DFFR_X1 \regfile/rx_10/data_out_reg[25]  ( .D(n3147), .CK(CLK), .RN(n6550), 
        .QN(n238) );
  DFFR_X1 \regfile/rx_10/data_out_reg[24]  ( .D(n3181), .CK(CLK), .RN(n7832), 
        .QN(n336) );
  DFFR_X1 \regfile/rx_10/data_out_reg[22]  ( .D(n3220), .CK(CLK), .RN(n7775), 
        .QN(n380) );
  DFFR_X1 \regfile/rx_10/data_out_reg[21]  ( .D(n3259), .CK(CLK), .RN(n6550), 
        .QN(n416) );
  DFFR_X1 \regfile/rx_10/data_out_reg[20]  ( .D(n3298), .CK(CLK), .RN(n7831), 
        .QN(n451) );
  DFFR_X1 \regfile/rx_10/data_out_reg[19]  ( .D(n3337), .CK(CLK), .RN(n7766), 
        .QN(n486) );
  DFFR_X1 \regfile/rx_10/data_out_reg[18]  ( .D(n3376), .CK(CLK), .RN(n6550), 
        .QN(n521) );
  DFFR_X1 \regfile/rx_10/data_out_reg[17]  ( .D(n3415), .CK(CLK), .RN(n7830), 
        .QN(n556) );
  DFFR_X1 \regfile/rx_10/data_out_reg[16]  ( .D(n3454), .CK(CLK), .RN(n7767), 
        .QN(n591) );
  DFFR_X1 \regfile/rx_10/data_out_reg[7]  ( .D(n3810), .CK(CLK), .RN(n6550), 
        .QN(n973) );
  DFFR_X1 \regfile/rx_10/data_out_reg[1]  ( .D(n4065), .CK(CLK), .RN(n7835), 
        .QN(n1190) );
  DFFR_X1 \regfile/rx_14/data_out_reg[23]  ( .D(n4036), .CK(CLK), .RN(n7768), 
        .QN(n1161) );
  DFFR_X1 \regfile/rx_13/data_out_reg[23]  ( .D(n4260), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][23] ), .QN(n1319) );
  DFFR_X1 \regfile/rx_10/data_out_reg[0]  ( .D(n4067), .CK(CLK), .RN(n7834), 
        .QN(n1192) );
  DFFR_X1 \regfile/rx_14/data_out_reg[30]  ( .D(n4030), .CK(CLK), .RN(n7769), 
        .QN(n1155) );
  DFFR_X1 \regfile/rx_14/data_out_reg[29]  ( .D(n4032), .CK(CLK), .RN(n6550), 
        .QN(n1157) );
  DFFR_X1 \regfile/rx_14/data_out_reg[28]  ( .D(n4033), .CK(CLK), .RN(n7833), 
        .QN(n1158) );
  DFFR_X1 \regfile/rx_14/data_out_reg[27]  ( .D(n4034), .CK(CLK), .RN(n7771), 
        .QN(n1159) );
  DFFR_X1 \regfile/rx_13/data_out_reg[30]  ( .D(n4254), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][30] ), .QN(n1313) );
  DFFR_X1 \regfile/rx_13/data_out_reg[29]  ( .D(n4256), .CK(CLK), .RN(n7838), 
        .Q(\regfile/reg_out[13][29] ), .QN(n1315) );
  DFFR_X1 \regfile/rx_13/data_out_reg[28]  ( .D(n4257), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[13][28] ), .QN(n1316) );
  DFFR_X1 \regfile/rx_13/data_out_reg[27]  ( .D(n4258), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][27] ), .QN(n1317) );
  DFFR_X1 \regfile/rx_14/data_out_reg[31]  ( .D(n4029), .CK(CLK), .RN(n7837), 
        .QN(n1154) );
  DFFR_X1 \regfile/rx_13/data_out_reg[31]  ( .D(n4253), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[13][31] ), .QN(n1312) );
  DFFR_X1 \regfile/rx_14/data_out_reg[26]  ( .D(n4035), .CK(CLK), .RN(n6550), 
        .QN(n1160) );
  DFFR_X1 \regfile/rx_14/data_out_reg[25]  ( .D(n3151), .CK(CLK), .RN(n7836), 
        .QN(n250) );
  DFFR_X1 \regfile/rx_14/data_out_reg[24]  ( .D(n3185), .CK(CLK), .RN(n7799), 
        .QN(n340) );
  DFFR_X1 \regfile/rx_13/data_out_reg[26]  ( .D(n4259), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][26] ), .QN(n1318) );
  DFFR_X1 \regfile/rx_13/data_out_reg[25]  ( .D(n3150), .CK(CLK), .RN(n7841), 
        .Q(\regfile/reg_out[13][25] ), .QN(n247) );
  DFFR_X1 \regfile/rx_13/data_out_reg[24]  ( .D(n3184), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[13][24] ), .QN(n339) );
  DFFR_X1 \regfile/rx_14/data_out_reg[22]  ( .D(n3224), .CK(CLK), .RN(n6550), 
        .QN(n384) );
  DFFR_X1 \regfile/rx_14/data_out_reg[21]  ( .D(n3263), .CK(CLK), .RN(n7840), 
        .QN(n420) );
  DFFR_X1 \regfile/rx_14/data_out_reg[20]  ( .D(n3302), .CK(CLK), .RN(n7788), 
        .QN(n455) );
  DFFR_X1 \regfile/rx_14/data_out_reg[19]  ( .D(n3341), .CK(CLK), .RN(n6550), 
        .QN(n490) );
  DFFR_X1 \regfile/rx_14/data_out_reg[18]  ( .D(n3380), .CK(CLK), .RN(n7839), 
        .QN(n525) );
  DFFR_X1 \regfile/rx_14/data_out_reg[17]  ( .D(n3419), .CK(CLK), .RN(n7794), 
        .QN(n560) );
  DFFR_X1 \regfile/rx_14/data_out_reg[16]  ( .D(n3458), .CK(CLK), .RN(n6550), 
        .QN(n595) );
  DFFR_X1 \regfile/rx_13/data_out_reg[22]  ( .D(n3223), .CK(CLK), .RN(n7843), 
        .Q(\regfile/reg_out[13][22] ), .QN(n383) );
  DFFR_X1 \regfile/rx_13/data_out_reg[21]  ( .D(n3262), .CK(CLK), .RN(n7784), 
        .Q(\regfile/reg_out[13][21] ), .QN(n419) );
  DFFR_X1 \regfile/rx_13/data_out_reg[20]  ( .D(n3301), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][20] ), .QN(n454) );
  DFFR_X1 \regfile/rx_13/data_out_reg[19]  ( .D(n3340), .CK(CLK), .RN(n7842), 
        .Q(\regfile/reg_out[13][19] ), .QN(n489) );
  DFFR_X1 \regfile/rx_13/data_out_reg[18]  ( .D(n3379), .CK(CLK), .RN(n7785), 
        .Q(\regfile/reg_out[13][18] ), .QN(n524) );
  DFFR_X1 \regfile/rx_13/data_out_reg[17]  ( .D(n3418), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][17] ), .QN(n559) );
  DFFR_X1 \regfile/rx_13/data_out_reg[16]  ( .D(n3457), .CK(CLK), .RN(n7826), 
        .Q(\regfile/reg_out[13][16] ), .QN(n594) );
  DFFR_X1 \regfile/rx_14/data_out_reg[7]  ( .D(n3814), .CK(CLK), .RN(n7786), 
        .QN(n977) );
  DFFR_X1 \regfile/rx_14/data_out_reg[1]  ( .D(n4037), .CK(CLK), .RN(n6550), 
        .QN(n1162) );
  DFFR_X1 \regfile/rx_13/data_out_reg[7]  ( .D(n3813), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[13][7] ), .QN(n976) );
  DFFR_X1 \regfile/rx_13/data_out_reg[1]  ( .D(n4261), .CK(CLK), .RN(n7787), 
        .Q(\regfile/reg_out[13][1] ), .QN(n1320) );
  DFFR_X1 \regfile/rx_14/data_out_reg[0]  ( .D(n4039), .CK(CLK), .RN(n6550), 
        .QN(n1164) );
  DFFR_X1 \regfile/rx_13/data_out_reg[0]  ( .D(n4263), .CK(CLK), .RN(n7812), 
        .Q(\regfile/reg_out[13][0] ), .QN(n1322) );
  DFFR_X1 \regfile/rx_10/data_out_reg[14]  ( .D(n4066), .CK(CLK), .RN(n7788), 
        .QN(n1191) );
  DFFR_X1 \regfile/rx_10/data_out_reg[13]  ( .D(n3654), .CK(CLK), .RN(n6550), 
        .QN(n795) );
  DFFR_X1 \regfile/rx_10/data_out_reg[12]  ( .D(n3615), .CK(CLK), .RN(n7809), 
        .QN(n757) );
  DFFR_X1 \regfile/rx_10/data_out_reg[11]  ( .D(n3576), .CK(CLK), .RN(n7789), 
        .QN(n719) );
  DFFR_X1 \regfile/rx_10/data_out_reg[10]  ( .D(n3537), .CK(CLK), .RN(n6550), 
        .QN(n681) );
  DFFR_X1 \regfile/rx_10/data_out_reg[6]  ( .D(n3768), .CK(CLK), .RN(n7817), 
        .QN(n934) );
  DFFR_X1 \regfile/rx_10/data_out_reg[5]  ( .D(n3726), .CK(CLK), .RN(n7814), 
        .QN(n890) );
  DFFR_X1 \regfile/rx_10/data_out_reg[4]  ( .D(n4055), .CK(CLK), .RN(n6550), 
        .QN(n1180) );
  DFFR_X1 \regfile/rx_10/data_out_reg[3]  ( .D(n4056), .CK(CLK), .RN(n7815), 
        .QN(n1181) );
  DFFR_X1 \regfile/rx_10/data_out_reg[2]  ( .D(n4059), .CK(CLK), .RN(n7816), 
        .QN(n1184) );
  DFFR_X1 \regfile/rx_10/data_out_reg[15]  ( .D(n3496), .CK(CLK), .RN(n6550), 
        .QN(n632) );
  DFFR_X1 \regfile/rx_10/data_out_reg[9]  ( .D(n3852), .CK(CLK), .RN(n7793), 
        .QN(n1012) );
  DFFR_X1 \regfile/rx_10/data_out_reg[8]  ( .D(n4054), .CK(CLK), .RN(n7818), 
        .QN(n1179) );
  DFFR_X1 \regfile/rx_14/data_out_reg[14]  ( .D(n4038), .CK(CLK), .RN(n6550), 
        .QN(n1163) );
  DFFR_X1 \regfile/rx_14/data_out_reg[13]  ( .D(n3658), .CK(CLK), .RN(n7791), 
        .QN(n799) );
  DFFR_X1 \regfile/rx_14/data_out_reg[12]  ( .D(n3619), .CK(CLK), .RN(n7819), 
        .QN(n761) );
  DFFR_X1 \regfile/rx_14/data_out_reg[11]  ( .D(n3580), .CK(CLK), .RN(n6550), 
        .QN(n723) );
  DFFR_X1 \regfile/rx_14/data_out_reg[10]  ( .D(n3541), .CK(CLK), .RN(n7800), 
        .QN(n685) );
  DFFR_X1 \regfile/rx_13/data_out_reg[14]  ( .D(n4262), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[13][14] ), .QN(n1321) );
  DFFR_X1 \regfile/rx_13/data_out_reg[13]  ( .D(n3657), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][13] ), .QN(n798) );
  DFFR_X1 \regfile/rx_13/data_out_reg[12]  ( .D(n3618), .CK(CLK), .RN(n7797), 
        .Q(\regfile/reg_out[13][12] ), .QN(n760) );
  DFFR_X1 \regfile/rx_13/data_out_reg[11]  ( .D(n3579), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[13][11] ), .QN(n722) );
  DFFR_X1 \regfile/rx_13/data_out_reg[10]  ( .D(n3540), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][10] ), .QN(n684) );
  DFFR_X1 \regfile/rx_14/data_out_reg[6]  ( .D(n3772), .CK(CLK), .RN(n7776), 
        .QN(n938) );
  DFFR_X1 \regfile/rx_14/data_out_reg[5]  ( .D(n3730), .CK(CLK), .RN(n7802), 
        .QN(n894) );
  DFFR_X1 \regfile/rx_14/data_out_reg[4]  ( .D(n4027), .CK(CLK), .RN(n6550), 
        .QN(n1152) );
  DFFR_X1 \regfile/rx_14/data_out_reg[3]  ( .D(n4028), .CK(CLK), .RN(n7779), 
        .QN(n1153) );
  DFFR_X1 \regfile/rx_14/data_out_reg[2]  ( .D(n4031), .CK(CLK), .RN(n7804), 
        .QN(n1156) );
  DFFR_X1 \regfile/rx_13/data_out_reg[6]  ( .D(n3771), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][6] ), .QN(n937) );
  DFFR_X1 \regfile/rx_13/data_out_reg[5]  ( .D(n3729), .CK(CLK), .RN(n7753), 
        .Q(\regfile/reg_out[13][5] ), .QN(n893) );
  DFFR_X1 \regfile/rx_13/data_out_reg[4]  ( .D(n4251), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[13][4] ), .QN(n1310) );
  DFFR_X1 \regfile/rx_13/data_out_reg[3]  ( .D(n4252), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][3] ), .QN(n1311) );
  DFFR_X1 \regfile/rx_13/data_out_reg[2]  ( .D(n4255), .CK(CLK), .RN(n7750), 
        .Q(\regfile/reg_out[13][2] ), .QN(n1314) );
  DFFR_X1 \regfile/rx_14/data_out_reg[15]  ( .D(n3500), .CK(CLK), .RN(n7807), 
        .QN(n636) );
  DFFR_X1 \regfile/rx_14/data_out_reg[9]  ( .D(n3856), .CK(CLK), .RN(n6550), 
        .QN(n1016) );
  DFFR_X1 \regfile/rx_14/data_out_reg[8]  ( .D(n4026), .CK(CLK), .RN(n7748), 
        .QN(n1151) );
  DFFR_X1 \regfile/rx_13/data_out_reg[15]  ( .D(n3499), .CK(CLK), .RN(n7821), 
        .Q(\regfile/reg_out[13][15] ), .QN(n635) );
  DFFR_X1 \regfile/rx_13/data_out_reg[9]  ( .D(n3855), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[13][9] ), .QN(n1015) );
  DFFR_X1 \regfile/rx_13/data_out_reg[8]  ( .D(n4250), .CK(CLK), .RN(n7838), 
        .Q(\regfile/reg_out[13][8] ), .QN(n1309) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[25]  ( .D(n4401), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [25]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[24]  ( .D(n4400), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [24]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[23]  ( .D(n4399), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [23]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[22]  ( .D(n4398), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [22]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[21]  ( .D(n4397), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [21]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[20]  ( .D(n4396), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [20]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[19]  ( .D(n4394), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [19]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[18]  ( .D(n4392), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [18]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[17]  ( .D(n4391), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [17]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[16]  ( .D(n4389), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [16]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[15]  ( .D(n4388), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [15]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[14]  ( .D(n4387), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [14]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[13]  ( .D(n4386), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [13]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[12]  ( .D(n4385), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [12]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[11]  ( .D(n4384), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [11]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[10]  ( .D(n4383), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [10]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[9]  ( .D(n4382), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [9]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[8]  ( .D(n4381), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [8]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[7]  ( .D(n4380), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [7]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[6]  ( .D(n4379), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [6]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[5]  ( .D(n4378), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [5]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[2]  ( .D(n4369), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [2]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[1]  ( .D(n4365), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [1]) );
  DFFR_X1 \Mcontrol/ir_fd/data_out_reg[0]  ( .D(n4361), .CK(CLK), .RN(
        \Mcontrol/int_reset ), .Q(\Mcontrol/d_sampled_finstr [0]) );
  DFFR_X1 \regfile/rx_30/data_out_reg[23]  ( .D(n3924), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[30][23] ), .QN(n1103) );
  DFFR_X1 \regfile/rx_30/data_out_reg[30]  ( .D(n3918), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][30] ), .QN(n1097) );
  DFFR_X1 \regfile/rx_30/data_out_reg[29]  ( .D(n3920), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[30][29] ), .QN(n1099) );
  DFFR_X1 \regfile/rx_30/data_out_reg[28]  ( .D(n3921), .CK(CLK), .RN(n7851), 
        .Q(\regfile/reg_out[30][28] ), .QN(n1100) );
  DFFR_X1 \regfile/rx_30/data_out_reg[27]  ( .D(n3922), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][27] ), .QN(n1101) );
  DFFR_X1 \regfile/rx_30/data_out_reg[31]  ( .D(n3917), .CK(CLK), .RN(n7761), 
        .Q(\regfile/reg_out[30][31] ), .QN(n1096) );
  DFFR_X1 \regfile/rx_30/data_out_reg[26]  ( .D(n3923), .CK(CLK), .RN(n7742), 
        .Q(\regfile/reg_out[30][26] ), .QN(n1102) );
  DFFR_X1 \regfile/rx_30/data_out_reg[25]  ( .D(n3169), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][25] ), .QN(n296) );
  DFFR_X1 \regfile/rx_30/data_out_reg[24]  ( .D(n3203), .CK(CLK), .RN(n7735), 
        .Q(\regfile/reg_out[30][24] ), .QN(n350) );
  DFFR_X1 \regfile/rx_30/data_out_reg[22]  ( .D(n3242), .CK(CLK), .RN(n7738), 
        .Q(\regfile/reg_out[30][22] ), .QN(n394) );
  DFFR_X1 \regfile/rx_30/data_out_reg[21]  ( .D(n3281), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][21] ), .QN(n430) );
  DFFR_X1 \regfile/rx_30/data_out_reg[20]  ( .D(n3320), .CK(CLK), .RN(n7731), 
        .Q(\regfile/reg_out[30][20] ), .QN(n465) );
  DFFR_X1 \regfile/rx_30/data_out_reg[19]  ( .D(n3359), .CK(CLK), .RN(n7843), 
        .Q(\regfile/reg_out[30][19] ), .QN(n500) );
  DFFR_X1 \regfile/rx_30/data_out_reg[18]  ( .D(n3398), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][18] ), .QN(n535) );
  DFFR_X1 \regfile/rx_30/data_out_reg[17]  ( .D(n3437), .CK(CLK), .RN(n7723), 
        .Q(\regfile/reg_out[30][17] ), .QN(n570) );
  DFFR_X1 \regfile/rx_30/data_out_reg[16]  ( .D(n3476), .CK(CLK), .RN(n7839), 
        .Q(\regfile/reg_out[30][16] ), .QN(n605) );
  DFFR_X1 \regfile/rx_30/data_out_reg[7]  ( .D(n3832), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][7] ), .QN(n987) );
  DFFR_X1 \regfile/rx_30/data_out_reg[1]  ( .D(n3925), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[30][1] ), .QN(n1104) );
  DFFR_X1 \regfile/rx_30/data_out_reg[0]  ( .D(n3927), .CK(CLK), .RN(n7840), 
        .Q(\regfile/reg_out[30][0] ), .QN(n1106) );
  DFFR_X1 \regfile/rx_30/data_out_reg[14]  ( .D(n3926), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][14] ), .QN(n1105) );
  DFFR_X1 \regfile/rx_30/data_out_reg[13]  ( .D(n3676), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[30][13] ), .QN(n809) );
  DFFR_X1 \regfile/rx_30/data_out_reg[12]  ( .D(n3637), .CK(CLK), .RN(n7841), 
        .Q(\regfile/reg_out[30][12] ), .QN(n771) );
  DFFR_X1 \regfile/rx_30/data_out_reg[11]  ( .D(n3598), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][11] ), .QN(n733) );
  DFFR_X1 \regfile/rx_30/data_out_reg[10]  ( .D(n3559), .CK(CLK), .RN(n7824), 
        .Q(\regfile/reg_out[30][10] ), .QN(n695) );
  DFFR_X1 \regfile/rx_30/data_out_reg[6]  ( .D(n3790), .CK(CLK), .RN(n7836), 
        .Q(\regfile/reg_out[30][6] ), .QN(n948) );
  DFFR_X1 \regfile/rx_30/data_out_reg[5]  ( .D(n3748), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][5] ), .QN(n904) );
  DFFR_X1 \regfile/rx_30/data_out_reg[4]  ( .D(n3915), .CK(CLK), .RN(n7850), 
        .Q(\regfile/reg_out[30][4] ), .QN(n1094) );
  DFFR_X1 \regfile/rx_30/data_out_reg[3]  ( .D(n3916), .CK(CLK), .RN(n7837), 
        .Q(\regfile/reg_out[30][3] ), .QN(n1095) );
  DFFR_X1 \regfile/rx_30/data_out_reg[2]  ( .D(n3919), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][2] ), .QN(n1098) );
  DFFR_X1 \regfile/rx_30/data_out_reg[15]  ( .D(n3518), .CK(CLK), .RN(n7849), 
        .Q(\regfile/reg_out[30][15] ), .QN(n646) );
  DFFR_X1 \regfile/rx_30/data_out_reg[9]  ( .D(n3874), .CK(CLK), .RN(n7838), 
        .Q(\regfile/reg_out[30][9] ), .QN(n1026) );
  DFFR_X1 \regfile/rx_30/data_out_reg[8]  ( .D(n3914), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[30][8] ), .QN(n1093) );
  DFFR_X1 \regfile/rx_7/data_out_reg[31]  ( .D(n4295), .CK(CLK), .RN(n7848), 
        .QN(n1354) );
  DFFR_X1 \regfile/rx_7/data_out_reg[30]  ( .D(n4296), .CK(CLK), .RN(n7833), 
        .QN(n1355) );
  DFFR_X1 \regfile/rx_7/data_out_reg[29]  ( .D(n4298), .CK(CLK), .RN(n6550), 
        .QN(n1357) );
  DFFR_X1 \regfile/rx_7/data_out_reg[28]  ( .D(n4299), .CK(CLK), .RN(n7847), 
        .QN(n1358) );
  DFFR_X1 \regfile/rx_7/data_out_reg[27]  ( .D(n4300), .CK(CLK), .RN(n7834), 
        .QN(n1359) );
  DFFR_X1 \regfile/rx_7/data_out_reg[26]  ( .D(n4301), .CK(CLK), .RN(n6550), 
        .QN(n1360) );
  DFFR_X1 \regfile/rx_7/data_out_reg[25]  ( .D(n3175), .CK(CLK), .RN(n7846), 
        .QN(n312) );
  DFFR_X1 \regfile/rx_7/data_out_reg[24]  ( .D(n3209), .CK(CLK), .RN(n7835), 
        .QN(n354) );
  DFFR_X1 \regfile/rx_7/data_out_reg[23]  ( .D(n4302), .CK(CLK), .RN(n6550), 
        .QN(n1361) );
  DFFR_X1 \regfile/rx_7/data_out_reg[22]  ( .D(n3248), .CK(CLK), .RN(n7738), 
        .QN(n398) );
  DFFR_X1 \regfile/rx_7/data_out_reg[21]  ( .D(n3287), .CK(CLK), .RN(n7830), 
        .QN(n434) );
  DFFR_X1 \regfile/rx_7/data_out_reg[20]  ( .D(n3326), .CK(CLK), .RN(n6550), 
        .QN(n469) );
  DFFR_X1 \regfile/rx_7/data_out_reg[19]  ( .D(n3365), .CK(CLK), .RN(n7742), 
        .QN(n504) );
  DFFR_X1 \regfile/rx_7/data_out_reg[18]  ( .D(n3404), .CK(CLK), .RN(n7831), 
        .QN(n539) );
  DFFR_X1 \regfile/rx_7/data_out_reg[17]  ( .D(n3443), .CK(CLK), .RN(n6550), 
        .QN(n574) );
  DFFR_X1 \regfile/rx_7/data_out_reg[16]  ( .D(n3482), .CK(CLK), .RN(n7823), 
        .QN(n609) );
  DFFR_X1 \regfile/rx_7/data_out_reg[6]  ( .D(n3796), .CK(CLK), .RN(n7832), 
        .QN(n952) );
  DFFR_X1 \regfile/rx_7/data_out_reg[5]  ( .D(n3754), .CK(CLK), .RN(n6550), 
        .QN(n908) );
  DFFR_X1 \regfile/rx_7/data_out_reg[4]  ( .D(n4293), .CK(CLK), .RN(n7852), 
        .QN(n1352) );
  DFFR_X1 \regfile/rx_7/data_out_reg[3]  ( .D(n4294), .CK(CLK), .RN(n7827), 
        .QN(n1353) );
  DFFR_X1 \regfile/rx_7/data_out_reg[2]  ( .D(n4297), .CK(CLK), .RN(n6550), 
        .QN(n1356) );
  DFFR_X1 \regfile/rx_7/data_out_reg[15]  ( .D(n3524), .CK(CLK), .RN(n7825), 
        .QN(n650) );
  DFFR_X1 \regfile/rx_7/data_out_reg[14]  ( .D(n4304), .CK(CLK), .RN(n7828), 
        .QN(n1363) );
  DFFR_X1 \regfile/rx_7/data_out_reg[13]  ( .D(n3682), .CK(CLK), .RN(n6550), 
        .QN(n813) );
  DFFR_X1 \regfile/rx_7/data_out_reg[12]  ( .D(n3643), .CK(CLK), .RN(n7851), 
        .QN(n775) );
  DFFR_X1 \regfile/rx_7/data_out_reg[11]  ( .D(n3604), .CK(CLK), .RN(n7829), 
        .QN(n737) );
  DFFR_X1 \regfile/rx_7/data_out_reg[10]  ( .D(n3565), .CK(CLK), .RN(n6550), 
        .QN(n699) );
  DFFR_X1 \regfile/rx_7/data_out_reg[9]  ( .D(n3880), .CK(CLK), .RN(n7743), 
        .QN(n1030) );
  DFFR_X1 \regfile/rx_7/data_out_reg[8]  ( .D(n4292), .CK(CLK), .RN(n7826), 
        .QN(n1351) );
  DFFR_X1 \regfile/rx_7/data_out_reg[7]  ( .D(n3838), .CK(CLK), .RN(n6550), 
        .QN(n991) );
  DFFR_X1 \regfile/rx_7/data_out_reg[1]  ( .D(n4303), .CK(CLK), .RN(n7826), 
        .QN(n1362) );
  DFFR_X1 \regfile/rx_7/data_out_reg[0]  ( .D(n4305), .CK(CLK), .RN(n7842), 
        .QN(n1364) );
  DFFR_X1 \regfile/rx_16/data_out_reg[23]  ( .D(n4022), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][23] ), .QN(n1147) );
  DFFR_X1 \regfile/rx_16/data_out_reg[30]  ( .D(n4016), .CK(CLK), .RN(n7829), 
        .Q(\regfile/reg_out[16][30] ), .QN(n1141) );
  DFFR_X1 \regfile/rx_16/data_out_reg[29]  ( .D(n4018), .CK(CLK), .RN(n7845), 
        .Q(\regfile/reg_out[16][29] ), .QN(n1143) );
  DFFR_X1 \regfile/rx_16/data_out_reg[28]  ( .D(n4019), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][28] ), .QN(n1144) );
  DFFR_X1 \regfile/rx_16/data_out_reg[27]  ( .D(n4020), .CK(CLK), .RN(n7828), 
        .Q(\regfile/reg_out[16][27] ), .QN(n1145) );
  DFFR_X1 \regfile/rx_16/data_out_reg[31]  ( .D(n4015), .CK(CLK), .RN(n7846), 
        .Q(\regfile/reg_out[16][31] ), .QN(n1140) );
  DFFR_X1 \regfile/rx_16/data_out_reg[26]  ( .D(n4021), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][26] ), .QN(n1146) );
  DFFR_X1 \regfile/rx_16/data_out_reg[25]  ( .D(n3153), .CK(CLK), .RN(n7827), 
        .Q(\regfile/reg_out[16][25] ), .QN(n256) );
  DFFR_X1 \regfile/rx_16/data_out_reg[24]  ( .D(n3187), .CK(CLK), .RN(n7847), 
        .Q(\regfile/reg_out[16][24] ), .QN(n342) );
  DFFR_X1 \regfile/rx_16/data_out_reg[22]  ( .D(n3226), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][22] ), .QN(n386) );
  DFFR_X1 \regfile/rx_16/data_out_reg[21]  ( .D(n3265), .CK(CLK), .RN(n7832), 
        .Q(\regfile/reg_out[16][21] ), .QN(n422) );
  DFFR_X1 \regfile/rx_16/data_out_reg[20]  ( .D(n3304), .CK(CLK), .RN(n7848), 
        .Q(\regfile/reg_out[16][20] ), .QN(n457) );
  DFFR_X1 \regfile/rx_16/data_out_reg[19]  ( .D(n3343), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][19] ), .QN(n492) );
  DFFR_X1 \regfile/rx_16/data_out_reg[18]  ( .D(n3382), .CK(CLK), .RN(n7831), 
        .Q(\regfile/reg_out[16][18] ), .QN(n527) );
  DFFR_X1 \regfile/rx_16/data_out_reg[17]  ( .D(n3421), .CK(CLK), .RN(n7849), 
        .Q(\regfile/reg_out[16][17] ), .QN(n562) );
  DFFR_X1 \regfile/rx_16/data_out_reg[16]  ( .D(n3460), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][16] ), .QN(n597) );
  DFFR_X1 \regfile/rx_16/data_out_reg[7]  ( .D(n3816), .CK(CLK), .RN(n7830), 
        .Q(\regfile/reg_out[16][7] ), .QN(n979) );
  DFFR_X1 \regfile/rx_16/data_out_reg[1]  ( .D(n4023), .CK(CLK), .RN(n7850), 
        .Q(\regfile/reg_out[16][1] ), .QN(n1148) );
  DFFR_X1 \regfile/rx_16/data_out_reg[0]  ( .D(n4025), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][0] ), .QN(n1150) );
  DFFR_X1 \regfile/rx_16/data_out_reg[14]  ( .D(n4024), .CK(CLK), .RN(n7835), 
        .Q(\regfile/reg_out[16][14] ), .QN(n1149) );
  DFFR_X1 \regfile/rx_16/data_out_reg[13]  ( .D(n3660), .CK(CLK), .RN(n7823), 
        .Q(\regfile/reg_out[16][13] ), .QN(n801) );
  DFFR_X1 \regfile/rx_16/data_out_reg[12]  ( .D(n3621), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][12] ), .QN(n763) );
  DFFR_X1 \regfile/rx_16/data_out_reg[11]  ( .D(n3582), .CK(CLK), .RN(n7834), 
        .Q(\regfile/reg_out[16][11] ), .QN(n725) );
  DFFR_X1 \regfile/rx_16/data_out_reg[10]  ( .D(n3543), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[16][10] ), .QN(n687) );
  DFFR_X1 \regfile/rx_16/data_out_reg[6]  ( .D(n3774), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][6] ), .QN(n940) );
  DFFR_X1 \regfile/rx_16/data_out_reg[5]  ( .D(n3732), .CK(CLK), .RN(n7833), 
        .Q(\regfile/reg_out[16][5] ), .QN(n896) );
  DFFR_X1 \regfile/rx_16/data_out_reg[4]  ( .D(n4013), .CK(CLK), .RN(n7723), 
        .Q(\regfile/reg_out[16][4] ), .QN(n1138) );
  DFFR_X1 \regfile/rx_16/data_out_reg[3]  ( .D(n4014), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[16][3] ), .QN(n1139) );
  DFFR_X1 \regfile/rx_16/data_out_reg[2]  ( .D(n4017), .CK(CLK), .RN(n7838), 
        .Q(\regfile/reg_out[16][2] ), .QN(n1142) );
  DFFR_X1 \regfile/rx_16/data_out_reg[15]  ( .D(n3502), .CK(CLK), .RN(n7735), 
        .Q(\regfile/reg_out[16][15] ), .QN(n638) );
  DFFR_X1 \regfile/rx_16/data_out_reg[9]  ( .D(n3858), .CK(CLK), .RN(n7837), 
        .Q(\regfile/reg_out[16][9] ), .QN(n1018) );
  DFFR_X1 \regfile/rx_16/data_out_reg[8]  ( .D(n4012), .CK(CLK), .RN(n7836), 
        .Q(\regfile/reg_out[16][8] ), .QN(n1137) );
  DFFR_X1 \regfile/rx_17/data_out_reg[23]  ( .D(n4232), .CK(CLK), .RN(n7761), 
        .Q(\regfile/reg_out[17][23] ), .QN(n1291) );
  DFFR_X1 \regfile/rx_17/data_out_reg[30]  ( .D(n4226), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][30] ), .QN(n1285) );
  DFFR_X1 \regfile/rx_17/data_out_reg[29]  ( .D(n4228), .CK(CLK), .RN(n7841), 
        .Q(\regfile/reg_out[17][29] ), .QN(n1287) );
  DFFR_X1 \regfile/rx_17/data_out_reg[28]  ( .D(n4229), .CK(CLK), .RN(n7837), 
        .Q(\regfile/reg_out[17][28] ), .QN(n1288) );
  DFFR_X1 \regfile/rx_17/data_out_reg[27]  ( .D(n4230), .CK(CLK), .RN(n7823), 
        .Q(\regfile/reg_out[17][27] ), .QN(n1289) );
  DFFR_X1 \regfile/rx_17/data_out_reg[31]  ( .D(n4225), .CK(CLK), .RN(n7790), 
        .Q(\regfile/reg_out[17][31] ), .QN(n1284) );
  DFFR_X1 \regfile/rx_17/data_out_reg[26]  ( .D(n4231), .CK(CLK), .RN(n7840), 
        .Q(\regfile/reg_out[17][26] ), .QN(n1290) );
  DFFR_X1 \regfile/rx_17/data_out_reg[25]  ( .D(n3154), .CK(CLK), .RN(n7787), 
        .Q(\regfile/reg_out[17][25] ), .QN(n259) );
  DFFR_X1 \regfile/rx_17/data_out_reg[24]  ( .D(n3188), .CK(CLK), .RN(n7851), 
        .Q(\regfile/reg_out[17][24] ), .QN(n343) );
  DFFR_X1 \regfile/rx_17/data_out_reg[22]  ( .D(n3227), .CK(CLK), .RN(n7839), 
        .Q(\regfile/reg_out[17][22] ), .QN(n387) );
  DFFR_X1 \regfile/rx_17/data_out_reg[21]  ( .D(n3266), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][21] ), .QN(n423) );
  DFFR_X1 \regfile/rx_17/data_out_reg[20]  ( .D(n3305), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][20] ), .QN(n458) );
  DFFR_X1 \regfile/rx_17/data_out_reg[19]  ( .D(n3344), .CK(CLK), .RN(n7843), 
        .Q(\regfile/reg_out[17][19] ), .QN(n493) );
  DFFR_X1 \regfile/rx_17/data_out_reg[18]  ( .D(n3383), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][18] ), .QN(n528) );
  DFFR_X1 \regfile/rx_17/data_out_reg[17]  ( .D(n3422), .CK(CLK), .RN(n7842), 
        .Q(\regfile/reg_out[17][17] ), .QN(n563) );
  DFFR_X1 \regfile/rx_17/data_out_reg[16]  ( .D(n3461), .CK(CLK), .RN(n7823), 
        .Q(\regfile/reg_out[17][16] ), .QN(n598) );
  DFFR_X1 \regfile/rx_17/data_out_reg[7]  ( .D(n3817), .CK(CLK), .RN(n7793), 
        .Q(\regfile/reg_out[17][7] ), .QN(n980) );
  DFFR_X1 \regfile/rx_17/data_out_reg[1]  ( .D(n4233), .CK(CLK), .RN(n7815), 
        .Q(\regfile/reg_out[17][1] ), .QN(n1292) );
  DFFR_X1 \regfile/rx_17/data_out_reg[0]  ( .D(n4235), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[17][0] ), .QN(n1294) );
  DFFR_X1 \regfile/rx_17/data_out_reg[14]  ( .D(n4234), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][14] ), .QN(n1293) );
  DFFR_X1 \regfile/rx_17/data_out_reg[13]  ( .D(n3661), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[17][13] ), .QN(n802) );
  DFFR_X1 \regfile/rx_17/data_out_reg[12]  ( .D(n3622), .CK(CLK), .RN(n7809), 
        .Q(\regfile/reg_out[17][12] ), .QN(n764) );
  DFFR_X1 \regfile/rx_17/data_out_reg[11]  ( .D(n3583), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][11] ), .QN(n726) );
  DFFR_X1 \regfile/rx_17/data_out_reg[10]  ( .D(n3544), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[17][10] ), .QN(n688) );
  DFFR_X1 \regfile/rx_17/data_out_reg[6]  ( .D(n3775), .CK(CLK), .RN(n7812), 
        .Q(\regfile/reg_out[17][6] ), .QN(n941) );
  DFFR_X1 \regfile/rx_17/data_out_reg[5]  ( .D(n3733), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][5] ), .QN(n897) );
  DFFR_X1 \regfile/rx_17/data_out_reg[4]  ( .D(n4223), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[17][4] ), .QN(n1282) );
  DFFR_X1 \regfile/rx_17/data_out_reg[3]  ( .D(n4224), .CK(CLK), .RN(n7824), 
        .Q(\regfile/reg_out[17][3] ), .QN(n1283) );
  DFFR_X1 \regfile/rx_17/data_out_reg[2]  ( .D(n4227), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][2] ), .QN(n1286) );
  DFFR_X1 \regfile/rx_17/data_out_reg[15]  ( .D(n3503), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[17][15] ), .QN(n639) );
  DFFR_X1 \regfile/rx_17/data_out_reg[9]  ( .D(n3859), .CK(CLK), .RN(n7844), 
        .Q(\regfile/reg_out[17][9] ), .QN(n1019) );
  DFFR_X1 \regfile/rx_17/data_out_reg[8]  ( .D(n4222), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[17][8] ), .QN(n1281) );
  DFFR_X1 \regfile/rx_12/data_out_reg[31]  ( .D(n4043), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[12][31] ), .QN(n1168) );
  DFFR_X1 \regfile/rx_12/data_out_reg[30]  ( .D(n4044), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[12][30] ), .QN(n1169) );
  DFFR_X1 \regfile/rx_12/data_out_reg[29]  ( .D(n4046), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][29] ), .QN(n1171) );
  DFFR_X1 \regfile/rx_12/data_out_reg[28]  ( .D(n4047), .CK(CLK), .RN(n7810), 
        .Q(\regfile/reg_out[12][28] ), .QN(n1172) );
  DFFR_X1 \regfile/rx_12/data_out_reg[27]  ( .D(n4048), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[12][27] ), .QN(n1173) );
  DFFR_X1 \regfile/rx_12/data_out_reg[26]  ( .D(n4049), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][26] ), .QN(n1174) );
  DFFR_X1 \regfile/rx_12/data_out_reg[25]  ( .D(n3149), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[12][25] ), .QN(n244) );
  DFFR_X1 \regfile/rx_12/data_out_reg[24]  ( .D(n3183), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[12][24] ), .QN(n338) );
  DFFR_X1 \regfile/rx_12/data_out_reg[23]  ( .D(n4050), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][23] ), .QN(n1175) );
  DFFR_X1 \regfile/rx_12/data_out_reg[22]  ( .D(n3222), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[12][22] ), .QN(n382) );
  DFFR_X1 \regfile/rx_12/data_out_reg[21]  ( .D(n3261), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[12][21] ), .QN(n418) );
  DFFR_X1 \regfile/rx_12/data_out_reg[20]  ( .D(n3300), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][20] ), .QN(n453) );
  DFFR_X1 \regfile/rx_12/data_out_reg[19]  ( .D(n3339), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[12][19] ), .QN(n488) );
  DFFR_X1 \regfile/rx_12/data_out_reg[18]  ( .D(n3378), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[12][18] ), .QN(n523) );
  DFFR_X1 \regfile/rx_12/data_out_reg[17]  ( .D(n3417), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][17] ), .QN(n558) );
  DFFR_X1 \regfile/rx_12/data_out_reg[16]  ( .D(n3456), .CK(CLK), .RN(n7816), 
        .Q(\regfile/reg_out[12][16] ), .QN(n593) );
  DFFR_X1 \regfile/rx_12/data_out_reg[6]  ( .D(n3770), .CK(CLK), .RN(n7721), 
        .Q(\regfile/reg_out[12][6] ), .QN(n936) );
  DFFR_X1 \regfile/rx_12/data_out_reg[5]  ( .D(n3728), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][5] ), .QN(n892) );
  DFFR_X1 \regfile/rx_12/data_out_reg[4]  ( .D(n4041), .CK(CLK), .RN(n7814), 
        .Q(\regfile/reg_out[12][4] ), .QN(n1166) );
  DFFR_X1 \regfile/rx_12/data_out_reg[3]  ( .D(n4042), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[12][3] ), .QN(n1167) );
  DFFR_X1 \regfile/rx_12/data_out_reg[2]  ( .D(n4045), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][2] ), .QN(n1170) );
  DFFR_X1 \regfile/rx_12/data_out_reg[15]  ( .D(n3498), .CK(CLK), .RN(n7789), 
        .Q(\regfile/reg_out[12][15] ), .QN(n634) );
  DFFR_X1 \regfile/rx_12/data_out_reg[14]  ( .D(n4052), .CK(CLK), .RN(n7746), 
        .Q(\regfile/reg_out[12][14] ), .QN(n1177) );
  DFFR_X1 \regfile/rx_12/data_out_reg[13]  ( .D(n3656), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][13] ), .QN(n797) );
  DFFR_X1 \regfile/rx_12/data_out_reg[12]  ( .D(n3617), .CK(CLK), .RN(n7788), 
        .Q(\regfile/reg_out[12][12] ), .QN(n759) );
  DFFR_X1 \regfile/rx_12/data_out_reg[11]  ( .D(n3578), .CK(CLK), .RN(n7747), 
        .Q(\regfile/reg_out[12][11] ), .QN(n721) );
  DFFR_X1 \regfile/rx_12/data_out_reg[10]  ( .D(n3539), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][10] ), .QN(n683) );
  DFFR_X1 \regfile/rx_12/data_out_reg[9]  ( .D(n3854), .CK(CLK), .RN(n7787), 
        .Q(\regfile/reg_out[12][9] ), .QN(n1014) );
  DFFR_X1 \regfile/rx_12/data_out_reg[8]  ( .D(n4040), .CK(CLK), .RN(n7737), 
        .Q(\regfile/reg_out[12][8] ), .QN(n1165) );
  DFFR_X1 \regfile/rx_12/data_out_reg[7]  ( .D(n3812), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[12][7] ), .QN(n975) );
  DFFR_X1 \regfile/rx_12/data_out_reg[1]  ( .D(n4051), .CK(CLK), .RN(n7786), 
        .Q(\regfile/reg_out[12][1] ), .QN(n1176) );
  DFFR_X1 \regfile/rx_12/data_out_reg[0]  ( .D(n4053), .CK(CLK), .RN(n7740), 
        .Q(\regfile/reg_out[12][0] ), .QN(n1178) );
  DFFR_X1 \regfile/rx_9/data_out_reg[31]  ( .D(n4281), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][31] ), .QN(n1340) );
  DFFR_X1 \regfile/rx_9/data_out_reg[30]  ( .D(n4282), .CK(CLK), .RN(n7785), 
        .Q(\regfile/reg_out[9][30] ), .QN(n1341) );
  DFFR_X1 \regfile/rx_9/data_out_reg[29]  ( .D(n4284), .CK(CLK), .RN(n7732), 
        .Q(\regfile/reg_out[9][29] ), .QN(n1343) );
  DFFR_X1 \regfile/rx_9/data_out_reg[28]  ( .D(n4285), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][28] ), .QN(n1344) );
  DFFR_X1 \regfile/rx_9/data_out_reg[27]  ( .D(n4286), .CK(CLK), .RN(n7784), 
        .Q(\regfile/reg_out[9][27] ), .QN(n1345) );
  DFFR_X1 \regfile/rx_9/data_out_reg[26]  ( .D(n4287), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[9][26] ), .QN(n1346) );
  DFFR_X1 \regfile/rx_9/data_out_reg[25]  ( .D(n3177), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][25] ), .QN(n318) );
  DFFR_X1 \regfile/rx_9/data_out_reg[24]  ( .D(n3211), .CK(CLK), .RN(n7795), 
        .Q(\regfile/reg_out[9][24] ), .QN(n356) );
  DFFR_X1 \regfile/rx_9/data_out_reg[23]  ( .D(n4288), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[9][23] ), .QN(n1347) );
  DFFR_X1 \regfile/rx_9/data_out_reg[22]  ( .D(n3250), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][22] ), .QN(n400) );
  DFFR_X1 \regfile/rx_9/data_out_reg[21]  ( .D(n3289), .CK(CLK), .RN(n7794), 
        .Q(\regfile/reg_out[9][21] ), .QN(n436) );
  DFFR_X1 \regfile/rx_9/data_out_reg[20]  ( .D(n3328), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[9][20] ), .QN(n471) );
  DFFR_X1 \regfile/rx_9/data_out_reg[19]  ( .D(n3367), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][19] ), .QN(n506) );
  DFFR_X1 \regfile/rx_9/data_out_reg[18]  ( .D(n3406), .CK(CLK), .RN(n7792), 
        .Q(\regfile/reg_out[9][18] ), .QN(n541) );
  DFFR_X1 \regfile/rx_9/data_out_reg[17]  ( .D(n3445), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[9][17] ), .QN(n576) );
  DFFR_X1 \regfile/rx_9/data_out_reg[16]  ( .D(n3484), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][16] ), .QN(n611) );
  DFFR_X1 \regfile/rx_9/data_out_reg[6]  ( .D(n3798), .CK(CLK), .RN(n7790), 
        .Q(\regfile/reg_out[9][6] ), .QN(n954) );
  DFFR_X1 \regfile/rx_9/data_out_reg[5]  ( .D(n3756), .CK(CLK), .RN(n7783), 
        .Q(\regfile/reg_out[9][5] ), .QN(n910) );
  DFFR_X1 \regfile/rx_9/data_out_reg[4]  ( .D(n4279), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][4] ), .QN(n1338) );
  DFFR_X1 \regfile/rx_9/data_out_reg[3]  ( .D(n4280), .CK(CLK), .RN(n7801), 
        .Q(\regfile/reg_out[9][3] ), .QN(n1339) );
  DFFR_X1 \regfile/rx_9/data_out_reg[2]  ( .D(n4283), .CK(CLK), .RN(n7772), 
        .Q(\regfile/reg_out[9][2] ), .QN(n1342) );
  DFFR_X1 \regfile/rx_9/data_out_reg[15]  ( .D(n3526), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][15] ), .QN(n652) );
  DFFR_X1 \regfile/rx_9/data_out_reg[14]  ( .D(n4290), .CK(CLK), .RN(n7799), 
        .Q(\regfile/reg_out[9][14] ), .QN(n1349) );
  DFFR_X1 \regfile/rx_9/data_out_reg[13]  ( .D(n3684), .CK(CLK), .RN(n7766), 
        .Q(\regfile/reg_out[9][13] ), .QN(n815) );
  DFFR_X1 \regfile/rx_9/data_out_reg[12]  ( .D(n3645), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][12] ), .QN(n777) );
  DFFR_X1 \regfile/rx_9/data_out_reg[11]  ( .D(n3606), .CK(CLK), .RN(n7798), 
        .Q(\regfile/reg_out[9][11] ), .QN(n739) );
  DFFR_X1 \regfile/rx_9/data_out_reg[10]  ( .D(n3567), .CK(CLK), .RN(n7767), 
        .Q(\regfile/reg_out[9][10] ), .QN(n701) );
  DFFR_X1 \regfile/rx_9/data_out_reg[9]  ( .D(n3882), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][9] ), .QN(n1032) );
  DFFR_X1 \regfile/rx_9/data_out_reg[8]  ( .D(n4278), .CK(CLK), .RN(n7796), 
        .Q(\regfile/reg_out[9][8] ), .QN(n1337) );
  DFFR_X1 \regfile/rx_9/data_out_reg[7]  ( .D(n3840), .CK(CLK), .RN(n7768), 
        .Q(\regfile/reg_out[9][7] ), .QN(n993) );
  DFFR_X1 \regfile/rx_9/data_out_reg[1]  ( .D(n4289), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[9][1] ), .QN(n1348) );
  DFFR_X1 \regfile/rx_9/data_out_reg[0]  ( .D(n4291), .CK(CLK), .RN(n7771), 
        .Q(\regfile/reg_out[9][0] ), .QN(n1350) );
  DFFR_X1 \regfile/rx_8/data_out_reg[31]  ( .D(n4071), .CK(CLK), .RN(n7769), 
        .QN(n1196) );
  DFFR_X1 \regfile/rx_8/data_out_reg[30]  ( .D(n4072), .CK(CLK), .RN(n6550), 
        .QN(n1197) );
  DFFR_X1 \regfile/rx_8/data_out_reg[29]  ( .D(n4074), .CK(CLK), .RN(n7769), 
        .QN(n1199) );
  DFFR_X1 \regfile/rx_8/data_out_reg[28]  ( .D(n4075), .CK(CLK), .RN(n7771), 
        .QN(n1200) );
  DFFR_X1 \regfile/rx_8/data_out_reg[27]  ( .D(n4076), .CK(CLK), .RN(n6550), 
        .QN(n1201) );
  DFFR_X1 \regfile/rx_8/data_out_reg[26]  ( .D(n4077), .CK(CLK), .RN(n7768), 
        .QN(n1202) );
  DFFR_X1 \regfile/rx_8/data_out_reg[25]  ( .D(n3176), .CK(CLK), .RN(n7796), 
        .QN(n315) );
  DFFR_X1 \regfile/rx_8/data_out_reg[24]  ( .D(n3210), .CK(CLK), .RN(n6550), 
        .QN(n355) );
  DFFR_X1 \regfile/rx_8/data_out_reg[23]  ( .D(n4078), .CK(CLK), .RN(n7767), 
        .QN(n1203) );
  DFFR_X1 \regfile/rx_8/data_out_reg[22]  ( .D(n3249), .CK(CLK), .RN(n7801), 
        .QN(n399) );
  DFFR_X1 \regfile/rx_8/data_out_reg[21]  ( .D(n3288), .CK(CLK), .RN(n6550), 
        .QN(n435) );
  DFFR_X1 \regfile/rx_8/data_out_reg[20]  ( .D(n3327), .CK(CLK), .RN(n7766), 
        .QN(n470) );
  DFFR_X1 \regfile/rx_8/data_out_reg[19]  ( .D(n3366), .CK(CLK), .RN(n7790), 
        .QN(n505) );
  DFFR_X1 \regfile/rx_8/data_out_reg[18]  ( .D(n3405), .CK(CLK), .RN(n6550), 
        .QN(n540) );
  DFFR_X1 \regfile/rx_8/data_out_reg[17]  ( .D(n3444), .CK(CLK), .RN(n7777), 
        .QN(n575) );
  DFFR_X1 \regfile/rx_8/data_out_reg[16]  ( .D(n3483), .CK(CLK), .RN(n7794), 
        .QN(n610) );
  DFFR_X1 \regfile/rx_8/data_out_reg[6]  ( .D(n3797), .CK(CLK), .RN(n6550), 
        .QN(n953) );
  DFFR_X1 \regfile/rx_8/data_out_reg[5]  ( .D(n3755), .CK(CLK), .RN(n7775), 
        .QN(n909) );
  DFFR_X1 \regfile/rx_8/data_out_reg[4]  ( .D(n4069), .CK(CLK), .RN(n7784), 
        .QN(n1194) );
  DFFR_X1 \regfile/rx_8/data_out_reg[3]  ( .D(n4070), .CK(CLK), .RN(n6550), 
        .QN(n1195) );
  DFFR_X1 \regfile/rx_8/data_out_reg[2]  ( .D(n4073), .CK(CLK), .RN(n7774), 
        .QN(n1198) );
  DFFR_X1 \regfile/rx_8/data_out_reg[15]  ( .D(n3525), .CK(CLK), .RN(n7785), 
        .QN(n651) );
  DFFR_X1 \regfile/rx_8/data_out_reg[14]  ( .D(n4080), .CK(CLK), .RN(n6550), 
        .QN(n1205) );
  DFFR_X1 \regfile/rx_8/data_out_reg[13]  ( .D(n3683), .CK(CLK), .RN(n7772), 
        .QN(n814) );
  DFFR_X1 \regfile/rx_8/data_out_reg[12]  ( .D(n3644), .CK(CLK), .RN(n7786), 
        .QN(n776) );
  DFFR_X1 \regfile/rx_8/data_out_reg[11]  ( .D(n3605), .CK(CLK), .RN(n6550), 
        .QN(n738) );
  DFFR_X1 \regfile/rx_8/data_out_reg[10]  ( .D(n3566), .CK(CLK), .RN(n7783), 
        .QN(n700) );
  DFFR_X1 \regfile/rx_8/data_out_reg[9]  ( .D(n3881), .CK(CLK), .RN(n7787), 
        .QN(n1031) );
  DFFR_X1 \regfile/rx_8/data_out_reg[8]  ( .D(n4068), .CK(CLK), .RN(n6550), 
        .QN(n1193) );
  DFFR_X1 \regfile/rx_8/data_out_reg[7]  ( .D(n3839), .CK(CLK), .RN(n7781), 
        .QN(n992) );
  DFFR_X1 \regfile/rx_8/data_out_reg[1]  ( .D(n4079), .CK(CLK), .RN(n7788), 
        .QN(n1204) );
  DFFR_X1 \regfile/rx_8/data_out_reg[0]  ( .D(n4081), .CK(CLK), .RN(n6550), 
        .QN(n1206) );
  DFFR_X1 \regfile/rx_27/data_out_reg[23]  ( .D(n4162), .CK(CLK), .RN(n7780), 
        .Q(\regfile/reg_out[27][23] ), .QN(n1263) );
  DFFR_X1 \regfile/rx_27/data_out_reg[30]  ( .D(n4156), .CK(CLK), .RN(n7789), 
        .Q(\regfile/reg_out[27][30] ), .QN(n1257) );
  DFFR_X1 \regfile/rx_27/data_out_reg[29]  ( .D(n4158), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][29] ), .QN(n1259) );
  DFFR_X1 \regfile/rx_27/data_out_reg[28]  ( .D(n4159), .CK(CLK), .RN(n7778), 
        .Q(\regfile/reg_out[27][28] ), .QN(n1260) );
  DFFR_X1 \regfile/rx_27/data_out_reg[27]  ( .D(n4160), .CK(CLK), .RN(n7814), 
        .Q(\regfile/reg_out[27][27] ), .QN(n1261) );
  DFFR_X1 \regfile/rx_27/data_out_reg[31]  ( .D(n4155), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][31] ), .QN(n1256) );
  DFFR_X1 \regfile/rx_27/data_out_reg[26]  ( .D(n4161), .CK(CLK), .RN(n7749), 
        .Q(\regfile/reg_out[27][26] ), .QN(n1262) );
  DFFR_X1 \regfile/rx_27/data_out_reg[25]  ( .D(n3165), .CK(CLK), .RN(n7818), 
        .Q(\regfile/reg_out[27][25] ), .QN(n286) );
  DFFR_X1 \regfile/rx_27/data_out_reg[24]  ( .D(n3199), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][24] ), .QN(n348) );
  DFFR_X1 \regfile/rx_27/data_out_reg[22]  ( .D(n3238), .CK(CLK), .RN(n7759), 
        .Q(\regfile/reg_out[27][22] ), .QN(n392) );
  DFFR_X1 \regfile/rx_27/data_out_reg[21]  ( .D(n3277), .CK(CLK), .RN(n7819), 
        .Q(\regfile/reg_out[27][21] ), .QN(n428) );
  DFFR_X1 \regfile/rx_27/data_out_reg[20]  ( .D(n3316), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][20] ), .QN(n463) );
  DFFR_X1 \regfile/rx_27/data_out_reg[19]  ( .D(n3355), .CK(CLK), .RN(n7757), 
        .Q(\regfile/reg_out[27][19] ), .QN(n498) );
  DFFR_X1 \regfile/rx_27/data_out_reg[18]  ( .D(n3394), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[27][18] ), .QN(n533) );
  DFFR_X1 \regfile/rx_27/data_out_reg[17]  ( .D(n3433), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][17] ), .QN(n568) );
  DFFR_X1 \regfile/rx_27/data_out_reg[16]  ( .D(n3472), .CK(CLK), .RN(n7756), 
        .Q(\regfile/reg_out[27][16] ), .QN(n603) );
  DFFR_X1 \regfile/rx_27/data_out_reg[7]  ( .D(n3828), .CK(CLK), .RN(n7811), 
        .Q(\regfile/reg_out[27][7] ), .QN(n985) );
  DFFR_X1 \regfile/rx_27/data_out_reg[1]  ( .D(n4163), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][1] ), .QN(n1264) );
  DFFR_X1 \regfile/rx_27/data_out_reg[0]  ( .D(n4165), .CK(CLK), .RN(n7765), 
        .Q(\regfile/reg_out[27][0] ), .QN(n1266) );
  DFFR_X1 \regfile/rx_27/data_out_reg[14]  ( .D(n4164), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[27][14] ), .QN(n1265) );
  DFFR_X1 \regfile/rx_27/data_out_reg[13]  ( .D(n3672), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][13] ), .QN(n807) );
  DFFR_X1 \regfile/rx_27/data_out_reg[12]  ( .D(n3633), .CK(CLK), .RN(n7764), 
        .Q(\regfile/reg_out[27][12] ), .QN(n769) );
  DFFR_X1 \regfile/rx_27/data_out_reg[11]  ( .D(n3594), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[27][11] ), .QN(n731) );
  DFFR_X1 \regfile/rx_27/data_out_reg[10]  ( .D(n3555), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][10] ), .QN(n693) );
  DFFR_X1 \regfile/rx_27/data_out_reg[6]  ( .D(n3786), .CK(CLK), .RN(n7762), 
        .Q(\regfile/reg_out[27][6] ), .QN(n946) );
  DFFR_X1 \regfile/rx_27/data_out_reg[5]  ( .D(n3744), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[27][5] ), .QN(n902) );
  DFFR_X1 \regfile/rx_27/data_out_reg[4]  ( .D(n4153), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][4] ), .QN(n1254) );
  DFFR_X1 \regfile/rx_27/data_out_reg[3]  ( .D(n4154), .CK(CLK), .RN(n7760), 
        .Q(\regfile/reg_out[27][3] ), .QN(n1255) );
  DFFR_X1 \regfile/rx_27/data_out_reg[2]  ( .D(n4157), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[27][2] ), .QN(n1258) );
  DFFR_X1 \regfile/rx_27/data_out_reg[15]  ( .D(n3514), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[27][15] ), .QN(n644) );
  DFFR_X1 \regfile/rx_27/data_out_reg[9]  ( .D(n3870), .CK(CLK), .RN(n7734), 
        .Q(\regfile/reg_out[27][9] ), .QN(n1024) );
  DFFR_X1 \regfile/rx_27/data_out_reg[8]  ( .D(n4152), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[27][8] ), .QN(n1253) );
  DFFR_X1 \regfile/rx_6/data_out_reg[23]  ( .D(n4092), .CK(CLK), .RN(n6550), 
        .QN(n1217) );
  DFFR_X1 \regfile/rx_6/data_out_reg[30]  ( .D(n4086), .CK(CLK), .RN(n7733), 
        .QN(n1211) );
  DFFR_X1 \regfile/rx_6/data_out_reg[29]  ( .D(n4088), .CK(CLK), .RN(n7743), 
        .QN(n1213) );
  DFFR_X1 \regfile/rx_6/data_out_reg[28]  ( .D(n4089), .CK(CLK), .RN(n6550), 
        .QN(n1214) );
  DFFR_X1 \regfile/rx_6/data_out_reg[27]  ( .D(n4090), .CK(CLK), .RN(n7732), 
        .QN(n1215) );
  DFFR_X1 \regfile/rx_6/data_out_reg[31]  ( .D(n4085), .CK(CLK), .RN(n7851), 
        .QN(n1210) );
  DFFR_X1 \regfile/rx_6/data_out_reg[26]  ( .D(n4091), .CK(CLK), .RN(n6550), 
        .QN(n1216) );
  DFFR_X1 \regfile/rx_6/data_out_reg[25]  ( .D(n3174), .CK(CLK), .RN(n7730), 
        .QN(n309) );
  DFFR_X1 \regfile/rx_6/data_out_reg[24]  ( .D(n3208), .CK(CLK), .RN(n7742), 
        .QN(n353) );
  DFFR_X1 \regfile/rx_6/data_out_reg[22]  ( .D(n3247), .CK(CLK), .RN(n6550), 
        .QN(n397) );
  DFFR_X1 \regfile/rx_6/data_out_reg[21]  ( .D(n3286), .CK(CLK), .RN(n7740), 
        .QN(n433) );
  DFFR_X1 \regfile/rx_6/data_out_reg[20]  ( .D(n3325), .CK(CLK), .RN(n7845), 
        .QN(n468) );
  DFFR_X1 \regfile/rx_6/data_out_reg[19]  ( .D(n3364), .CK(CLK), .RN(n6550), 
        .QN(n503) );
  DFFR_X1 \regfile/rx_6/data_out_reg[18]  ( .D(n3403), .CK(CLK), .RN(n7739), 
        .QN(n538) );
  DFFR_X1 \regfile/rx_6/data_out_reg[17]  ( .D(n3442), .CK(CLK), .RN(n7846), 
        .QN(n573) );
  DFFR_X1 \regfile/rx_6/data_out_reg[16]  ( .D(n3481), .CK(CLK), .RN(n6550), 
        .QN(n608) );
  DFFR_X1 \regfile/rx_6/data_out_reg[7]  ( .D(n3837), .CK(CLK), .RN(n7737), 
        .QN(n990) );
  DFFR_X1 \regfile/rx_6/data_out_reg[1]  ( .D(n4093), .CK(CLK), .RN(n7847), 
        .QN(n1218) );
  DFFR_X1 \regfile/rx_6/data_out_reg[0]  ( .D(n4095), .CK(CLK), .RN(n6550), 
        .QN(n1220) );
  DFFR_X1 \regfile/rx_6/data_out_reg[14]  ( .D(n4094), .CK(CLK), .RN(n7736), 
        .QN(n1219) );
  DFFR_X1 \regfile/rx_6/data_out_reg[13]  ( .D(n3681), .CK(CLK), .RN(n7848), 
        .QN(n812) );
  DFFR_X1 \regfile/rx_6/data_out_reg[12]  ( .D(n3642), .CK(CLK), .RN(n6550), 
        .QN(n774) );
  DFFR_X1 \regfile/rx_6/data_out_reg[11]  ( .D(n3603), .CK(CLK), .RN(n7747), 
        .QN(n736) );
  DFFR_X1 \regfile/rx_6/data_out_reg[10]  ( .D(n3564), .CK(CLK), .RN(n7849), 
        .QN(n698) );
  DFFR_X1 \regfile/rx_6/data_out_reg[6]  ( .D(n3795), .CK(CLK), .RN(n6550), 
        .QN(n951) );
  DFFR_X1 \regfile/rx_6/data_out_reg[5]  ( .D(n3753), .CK(CLK), .RN(n7746), 
        .QN(n907) );
  DFFR_X1 \regfile/rx_6/data_out_reg[4]  ( .D(n4083), .CK(CLK), .RN(n7850), 
        .QN(n1208) );
  DFFR_X1 \regfile/rx_6/data_out_reg[3]  ( .D(n4084), .CK(CLK), .RN(n6550), 
        .QN(n1209) );
  DFFR_X1 \regfile/rx_6/data_out_reg[2]  ( .D(n4087), .CK(CLK), .RN(n7722), 
        .QN(n1212) );
  DFFR_X1 \regfile/rx_6/data_out_reg[15]  ( .D(n3523), .CK(CLK), .RN(n7823), 
        .QN(n649) );
  DFFR_X1 \regfile/rx_6/data_out_reg[9]  ( .D(n3879), .CK(CLK), .RN(n6550), 
        .QN(n1029) );
  DFFR_X1 \regfile/rx_6/data_out_reg[8]  ( .D(n4082), .CK(CLK), .RN(n7721), 
        .QN(n1207) );
  DFFR_X1 \regfile/rx_23/data_out_reg[31]  ( .D(n4183), .CK(CLK), .RN(n7843), 
        .Q(\regfile/reg_out[23][31] ), .QN(n1270) );
  DFFR_X1 \regfile/rx_23/data_out_reg[30]  ( .D(n4184), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][30] ), .QN(n1271) );
  DFFR_X1 \regfile/rx_23/data_out_reg[29]  ( .D(n4186), .CK(CLK), .RN(n7719), 
        .Q(\regfile/reg_out[23][29] ), .QN(n1273) );
  DFFR_X1 \regfile/rx_23/data_out_reg[28]  ( .D(n4187), .CK(CLK), .RN(n7839), 
        .Q(\regfile/reg_out[23][28] ), .QN(n1274) );
  DFFR_X1 \regfile/rx_23/data_out_reg[27]  ( .D(n4188), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][27] ), .QN(n1275) );
  DFFR_X1 \regfile/rx_23/data_out_reg[26]  ( .D(n4189), .CK(CLK), .RN(n7718), 
        .Q(\regfile/reg_out[23][26] ), .QN(n1276) );
  DFFR_X1 \regfile/rx_23/data_out_reg[25]  ( .D(n3161), .CK(CLK), .RN(n7840), 
        .Q(\regfile/reg_out[23][25] ), .QN(n276) );
  DFFR_X1 \regfile/rx_23/data_out_reg[24]  ( .D(n3195), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][24] ), .QN(n346) );
  DFFR_X1 \regfile/rx_23/data_out_reg[23]  ( .D(n4190), .CK(CLK), .RN(n7728), 
        .Q(\regfile/reg_out[23][23] ), .QN(n1277) );
  DFFR_X1 \regfile/rx_23/data_out_reg[22]  ( .D(n3234), .CK(CLK), .RN(n7841), 
        .Q(\regfile/reg_out[23][22] ), .QN(n390) );
  DFFR_X1 \regfile/rx_23/data_out_reg[21]  ( .D(n3273), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][21] ), .QN(n426) );
  DFFR_X1 \regfile/rx_23/data_out_reg[20]  ( .D(n3312), .CK(CLK), .RN(n7727), 
        .Q(\regfile/reg_out[23][20] ), .QN(n461) );
  DFFR_X1 \regfile/rx_23/data_out_reg[19]  ( .D(n3351), .CK(CLK), .RN(n7794), 
        .Q(\regfile/reg_out[23][19] ), .QN(n496) );
  DFFR_X1 \regfile/rx_23/data_out_reg[18]  ( .D(n3390), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][18] ), .QN(n531) );
  DFFR_X1 \regfile/rx_23/data_out_reg[17]  ( .D(n3429), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][17] ), .QN(n566) );
  DFFR_X1 \regfile/rx_23/data_out_reg[16]  ( .D(n3468), .CK(CLK), .RN(n7850), 
        .Q(\regfile/reg_out[23][16] ), .QN(n601) );
  DFFR_X1 \regfile/rx_23/data_out_reg[6]  ( .D(n3782), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][6] ), .QN(n944) );
  DFFR_X1 \regfile/rx_23/data_out_reg[5]  ( .D(n3740), .CK(CLK), .RN(n7726), 
        .Q(\regfile/reg_out[23][5] ), .QN(n900) );
  DFFR_X1 \regfile/rx_23/data_out_reg[4]  ( .D(n4181), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][4] ), .QN(n1268) );
  DFFR_X1 \regfile/rx_23/data_out_reg[3]  ( .D(n4182), .CK(CLK), .RN(n7725), 
        .Q(\regfile/reg_out[23][3] ), .QN(n1269) );
  DFFR_X1 \regfile/rx_23/data_out_reg[2]  ( .D(n4185), .CK(CLK), .RN(n7724), 
        .Q(\regfile/reg_out[23][2] ), .QN(n1272) );
  DFFR_X1 \regfile/rx_23/data_out_reg[15]  ( .D(n3510), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][15] ), .QN(n642) );
  DFFR_X1 \regfile/rx_23/data_out_reg[14]  ( .D(n4192), .CK(CLK), .RN(n7791), 
        .Q(\regfile/reg_out[23][14] ), .QN(n1279) );
  DFFR_X1 \regfile/rx_23/data_out_reg[13]  ( .D(n3668), .CK(CLK), .RN(n7716), 
        .Q(\regfile/reg_out[23][13] ), .QN(n805) );
  DFFR_X1 \regfile/rx_23/data_out_reg[12]  ( .D(n3629), .CK(CLK), .RN(n7833), 
        .Q(\regfile/reg_out[23][12] ), .QN(n767) );
  DFFR_X1 \regfile/rx_23/data_out_reg[11]  ( .D(n3590), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][11] ), .QN(n729) );
  DFFR_X1 \regfile/rx_23/data_out_reg[10]  ( .D(n3551), .CK(CLK), .RN(n7821), 
        .Q(\regfile/reg_out[23][10] ), .QN(n691) );
  DFFR_X1 \regfile/rx_23/data_out_reg[9]  ( .D(n3866), .CK(CLK), .RN(n7834), 
        .Q(\regfile/reg_out[23][9] ), .QN(n1022) );
  DFFR_X1 \regfile/rx_23/data_out_reg[8]  ( .D(n4180), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][8] ), .QN(n1267) );
  DFFR_X1 \regfile/rx_23/data_out_reg[7]  ( .D(n3824), .CK(CLK), .RN(n7845), 
        .Q(\regfile/reg_out[23][7] ), .QN(n983) );
  DFFR_X1 \regfile/rx_23/data_out_reg[1]  ( .D(n4191), .CK(CLK), .RN(n7835), 
        .Q(\regfile/reg_out[23][1] ), .QN(n1278) );
  DFFR_X1 \regfile/rx_23/data_out_reg[0]  ( .D(n4193), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[23][0] ), .QN(n1280) );
  DFFR_X1 \regfile/rx_26/data_out_reg[23]  ( .D(n3952), .CK(CLK), .RN(n7844), 
        .Q(\regfile/reg_out[26][23] ), .QN(n1119) );
  DFFR_X1 \regfile/rx_26/data_out_reg[30]  ( .D(n3946), .CK(CLK), .RN(n7830), 
        .Q(\regfile/reg_out[26][30] ), .QN(n1113) );
  DFFR_X1 \regfile/rx_26/data_out_reg[29]  ( .D(n3948), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][29] ), .QN(n1115) );
  DFFR_X1 \regfile/rx_26/data_out_reg[28]  ( .D(n3949), .CK(CLK), .RN(n7744), 
        .Q(\regfile/reg_out[26][28] ), .QN(n1116) );
  DFFR_X1 \regfile/rx_26/data_out_reg[27]  ( .D(n3950), .CK(CLK), .RN(n7831), 
        .Q(\regfile/reg_out[26][27] ), .QN(n1117) );
  DFFR_X1 \regfile/rx_26/data_out_reg[31]  ( .D(n3945), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][31] ), .QN(n1112) );
  DFFR_X1 \regfile/rx_26/data_out_reg[26]  ( .D(n3951), .CK(CLK), .RN(n7822), 
        .Q(\regfile/reg_out[26][26] ), .QN(n1118) );
  DFFR_X1 \regfile/rx_26/data_out_reg[25]  ( .D(n3164), .CK(CLK), .RN(n7832), 
        .Q(\regfile/reg_out[26][25] ), .QN(n283) );
  DFFR_X1 \regfile/rx_26/data_out_reg[24]  ( .D(n3198), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][24] ), .QN(n347) );
  DFFR_X1 \regfile/rx_26/data_out_reg[22]  ( .D(n3237), .CK(CLK), .RN(n7824), 
        .Q(\regfile/reg_out[26][22] ), .QN(n391) );
  DFFR_X1 \regfile/rx_26/data_out_reg[21]  ( .D(n3276), .CK(CLK), .RN(n7827), 
        .Q(\regfile/reg_out[26][21] ), .QN(n427) );
  DFFR_X1 \regfile/rx_26/data_out_reg[20]  ( .D(n3315), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][20] ), .QN(n462) );
  DFFR_X1 \regfile/rx_26/data_out_reg[19]  ( .D(n3354), .CK(CLK), .RN(n7850), 
        .Q(\regfile/reg_out[26][19] ), .QN(n497) );
  DFFR_X1 \regfile/rx_26/data_out_reg[18]  ( .D(n3393), .CK(CLK), .RN(n7828), 
        .Q(\regfile/reg_out[26][18] ), .QN(n532) );
  DFFR_X1 \regfile/rx_26/data_out_reg[17]  ( .D(n3432), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][17] ), .QN(n567) );
  DFFR_X1 \regfile/rx_26/data_out_reg[16]  ( .D(n3471), .CK(CLK), .RN(n7849), 
        .Q(\regfile/reg_out[26][16] ), .QN(n602) );
  DFFR_X1 \regfile/rx_26/data_out_reg[7]  ( .D(n3827), .CK(CLK), .RN(n7829), 
        .Q(\regfile/reg_out[26][7] ), .QN(n984) );
  DFFR_X1 \regfile/rx_26/data_out_reg[1]  ( .D(n3953), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][1] ), .QN(n1120) );
  DFFR_X1 \regfile/rx_26/data_out_reg[0]  ( .D(n3955), .CK(CLK), .RN(n7848), 
        .Q(\regfile/reg_out[26][0] ), .QN(n1122) );
  DFFR_X1 \regfile/rx_26/data_out_reg[14]  ( .D(n3954), .CK(CLK), .RN(n7826), 
        .Q(\regfile/reg_out[26][14] ), .QN(n1121) );
  DFFR_X1 \regfile/rx_26/data_out_reg[13]  ( .D(n3671), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][13] ), .QN(n806) );
  DFFR_X1 \regfile/rx_26/data_out_reg[12]  ( .D(n3632), .CK(CLK), .RN(n7847), 
        .Q(\regfile/reg_out[26][12] ), .QN(n768) );
  DFFR_X1 \regfile/rx_26/data_out_reg[11]  ( .D(n3593), .CK(CLK), .RN(n7842), 
        .Q(\regfile/reg_out[26][11] ), .QN(n730) );
  DFFR_X1 \regfile/rx_26/data_out_reg[10]  ( .D(n3554), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][10] ), .QN(n692) );
  DFFR_X1 \regfile/rx_26/data_out_reg[6]  ( .D(n3785), .CK(CLK), .RN(n7846), 
        .Q(\regfile/reg_out[26][6] ), .QN(n945) );
  DFFR_X1 \regfile/rx_26/data_out_reg[5]  ( .D(n3743), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[26][5] ), .QN(n901) );
  DFFR_X1 \regfile/rx_26/data_out_reg[4]  ( .D(n3943), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][4] ), .QN(n1110) );
  DFFR_X1 \regfile/rx_26/data_out_reg[3]  ( .D(n3944), .CK(CLK), .RN(n7806), 
        .Q(\regfile/reg_out[26][3] ), .QN(n1111) );
  DFFR_X1 \regfile/rx_26/data_out_reg[2]  ( .D(n3947), .CK(CLK), .RN(n7761), 
        .Q(\regfile/reg_out[26][2] ), .QN(n1114) );
  DFFR_X1 \regfile/rx_26/data_out_reg[15]  ( .D(n3513), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[26][15] ), .QN(n643) );
  DFFR_X1 \regfile/rx_26/data_out_reg[9]  ( .D(n3869), .CK(CLK), .RN(n7803), 
        .Q(\regfile/reg_out[26][9] ), .QN(n1023) );
  DFFR_X1 \regfile/rx_26/data_out_reg[8]  ( .D(n3942), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[26][8] ), .QN(n1109) );
  DFFR_X1 \regfile/rx_15/data_out_reg[31]  ( .D(n4239), .CK(CLK), .RN(n6550), 
        .QN(n1298) );
  DFFR_X1 \regfile/rx_15/data_out_reg[30]  ( .D(n4240), .CK(CLK), .RN(n7812), 
        .QN(n1299) );
  DFFR_X1 \regfile/rx_15/data_out_reg[29]  ( .D(n4242), .CK(CLK), .RN(n7758), 
        .QN(n1301) );
  DFFR_X1 \regfile/rx_15/data_out_reg[28]  ( .D(n4243), .CK(CLK), .RN(n6550), 
        .QN(n1302) );
  DFFR_X1 \regfile/rx_15/data_out_reg[27]  ( .D(n4244), .CK(CLK), .RN(n7809), 
        .QN(n1303) );
  DFFR_X1 \regfile/rx_15/data_out_reg[26]  ( .D(n4245), .CK(CLK), .RN(n7776), 
        .QN(n1304) );
  DFFR_X1 \regfile/rx_15/data_out_reg[25]  ( .D(n3152), .CK(CLK), .RN(n6550), 
        .QN(n253) );
  DFFR_X1 \regfile/rx_15/data_out_reg[24]  ( .D(n3186), .CK(CLK), .RN(n7817), 
        .QN(n341) );
  DFFR_X1 \regfile/rx_15/data_out_reg[23]  ( .D(n4246), .CK(CLK), .RN(n7791), 
        .QN(n1305) );
  DFFR_X1 \regfile/rx_15/data_out_reg[22]  ( .D(n3225), .CK(CLK), .RN(n6550), 
        .QN(n385) );
  DFFR_X1 \regfile/rx_15/data_out_reg[21]  ( .D(n3264), .CK(CLK), .RN(n7815), 
        .QN(n421) );
  DFFR_X1 \regfile/rx_15/data_out_reg[20]  ( .D(n3303), .CK(CLK), .RN(n7815), 
        .QN(n456) );
  DFFR_X1 \regfile/rx_15/data_out_reg[19]  ( .D(n3342), .CK(CLK), .RN(n6550), 
        .QN(n491) );
  DFFR_X1 \regfile/rx_15/data_out_reg[18]  ( .D(n3381), .CK(CLK), .RN(n7793), 
        .QN(n526) );
  DFFR_X1 \regfile/rx_15/data_out_reg[17]  ( .D(n3420), .CK(CLK), .RN(n7809), 
        .QN(n561) );
  DFFR_X1 \regfile/rx_15/data_out_reg[16]  ( .D(n3459), .CK(CLK), .RN(n6550), 
        .QN(n596) );
  DFFR_X1 \regfile/rx_15/data_out_reg[6]  ( .D(n3773), .CK(CLK), .RN(n7791), 
        .QN(n939) );
  DFFR_X1 \regfile/rx_15/data_out_reg[5]  ( .D(n3731), .CK(CLK), .RN(n7812), 
        .QN(n895) );
  DFFR_X1 \regfile/rx_15/data_out_reg[4]  ( .D(n4237), .CK(CLK), .RN(n6550), 
        .QN(n1296) );
  DFFR_X1 \regfile/rx_15/data_out_reg[3]  ( .D(n4238), .CK(CLK), .RN(n7800), 
        .QN(n1297) );
  DFFR_X1 \regfile/rx_15/data_out_reg[2]  ( .D(n4241), .CK(CLK), .RN(n7824), 
        .QN(n1300) );
  DFFR_X1 \regfile/rx_15/data_out_reg[15]  ( .D(n3501), .CK(CLK), .RN(n6550), 
        .QN(n637) );
  DFFR_X1 \regfile/rx_15/data_out_reg[14]  ( .D(n4248), .CK(CLK), .RN(n7797), 
        .QN(n1307) );
  DFFR_X1 \regfile/rx_15/data_out_reg[13]  ( .D(n3659), .CK(CLK), .RN(n7844), 
        .QN(n800) );
  DFFR_X1 \regfile/rx_15/data_out_reg[12]  ( .D(n3620), .CK(CLK), .RN(n6550), 
        .QN(n762) );
  DFFR_X1 \regfile/rx_15/data_out_reg[11]  ( .D(n3581), .CK(CLK), .RN(n7770), 
        .QN(n724) );
  DFFR_X1 \regfile/rx_15/data_out_reg[10]  ( .D(n3542), .CK(CLK), .RN(n7727), 
        .QN(n686) );
  DFFR_X1 \regfile/rx_15/data_out_reg[9]  ( .D(n3857), .CK(CLK), .RN(n6550), 
        .QN(n1017) );
  DFFR_X1 \regfile/rx_15/data_out_reg[8]  ( .D(n4236), .CK(CLK), .RN(n7776), 
        .QN(n1295) );
  DFFR_X1 \regfile/rx_15/data_out_reg[7]  ( .D(n3815), .CK(CLK), .RN(n7728), 
        .QN(n978) );
  DFFR_X1 \regfile/rx_15/data_out_reg[1]  ( .D(n4247), .CK(CLK), .RN(n6550), 
        .QN(n1306) );
  DFFR_X1 \regfile/rx_15/data_out_reg[0]  ( .D(n4249), .CK(CLK), .RN(n6550), 
        .QN(n1308) );
  DFFR_X1 \regfile/rx_11/data_out_reg[31]  ( .D(n4267), .CK(CLK), .RN(n7721), 
        .QN(n1326) );
  DFFR_X1 \regfile/rx_11/data_out_reg[30]  ( .D(n4268), .CK(CLK), .RN(n6550), 
        .QN(n1327) );
  DFFR_X1 \regfile/rx_11/data_out_reg[29]  ( .D(n4270), .CK(CLK), .RN(n7782), 
        .QN(n1329) );
  DFFR_X1 \regfile/rx_11/data_out_reg[28]  ( .D(n4271), .CK(CLK), .RN(n7746), 
        .QN(n1330) );
  DFFR_X1 \regfile/rx_11/data_out_reg[27]  ( .D(n4272), .CK(CLK), .RN(n6550), 
        .QN(n1331) );
  DFFR_X1 \regfile/rx_11/data_out_reg[26]  ( .D(n4273), .CK(CLK), .RN(n7779), 
        .QN(n1332) );
  DFFR_X1 \regfile/rx_11/data_out_reg[25]  ( .D(n3148), .CK(CLK), .RN(n7747), 
        .QN(n241) );
  DFFR_X1 \regfile/rx_11/data_out_reg[24]  ( .D(n3182), .CK(CLK), .RN(n6550), 
        .QN(n337) );
  DFFR_X1 \regfile/rx_11/data_out_reg[23]  ( .D(n4274), .CK(CLK), .RN(n7753), 
        .QN(n1333) );
  DFFR_X1 \regfile/rx_11/data_out_reg[22]  ( .D(n3221), .CK(CLK), .RN(n7732), 
        .QN(n381) );
  DFFR_X1 \regfile/rx_11/data_out_reg[21]  ( .D(n3260), .CK(CLK), .RN(n6550), 
        .QN(n417) );
  DFFR_X1 \regfile/rx_11/data_out_reg[20]  ( .D(n3299), .CK(CLK), .RN(n7750), 
        .QN(n452) );
  DFFR_X1 \regfile/rx_11/data_out_reg[19]  ( .D(n3338), .CK(CLK), .RN(n7760), 
        .QN(n487) );
  DFFR_X1 \regfile/rx_11/data_out_reg[18]  ( .D(n3377), .CK(CLK), .RN(n6550), 
        .QN(n522) );
  DFFR_X1 \regfile/rx_11/data_out_reg[17]  ( .D(n3416), .CK(CLK), .RN(n7748), 
        .QN(n557) );
  DFFR_X1 \regfile/rx_11/data_out_reg[16]  ( .D(n3455), .CK(CLK), .RN(n7783), 
        .QN(n592) );
  DFFR_X1 \regfile/rx_11/data_out_reg[6]  ( .D(n3769), .CK(CLK), .RN(n6550), 
        .QN(n935) );
  DFFR_X1 \regfile/rx_11/data_out_reg[5]  ( .D(n3727), .CK(CLK), .RN(n7758), 
        .QN(n891) );
  DFFR_X1 \regfile/rx_11/data_out_reg[4]  ( .D(n4265), .CK(CLK), .RN(n7767), 
        .QN(n1324) );
  DFFR_X1 \regfile/rx_11/data_out_reg[3]  ( .D(n4266), .CK(CLK), .RN(n6550), 
        .QN(n1325) );
  DFFR_X1 \regfile/rx_11/data_out_reg[2]  ( .D(n4269), .CK(CLK), .RN(n7763), 
        .QN(n1328) );
  DFFR_X1 \regfile/rx_11/data_out_reg[15]  ( .D(n3497), .CK(CLK), .RN(n7758), 
        .QN(n633) );
  DFFR_X1 \regfile/rx_11/data_out_reg[14]  ( .D(n4276), .CK(CLK), .RN(n7761), 
        .QN(n1335) );
  DFFR_X1 \regfile/rx_11/data_out_reg[13]  ( .D(n3655), .CK(CLK), .RN(n7735), 
        .QN(n796) );
  DFFR_X1 \regfile/rx_11/data_out_reg[12]  ( .D(n3616), .CK(CLK), .RN(n7844), 
        .QN(n758) );
  DFFR_X1 \regfile/rx_11/data_out_reg[11]  ( .D(n3577), .CK(CLK), .RN(n6550), 
        .QN(n720) );
  DFFR_X1 \regfile/rx_11/data_out_reg[10]  ( .D(n3538), .CK(CLK), .RN(n7731), 
        .QN(n682) );
  DFFR_X1 \regfile/rx_11/data_out_reg[9]  ( .D(n3853), .CK(CLK), .RN(n7786), 
        .QN(n1013) );
  DFFR_X1 \regfile/rx_11/data_out_reg[8]  ( .D(n4264), .CK(CLK), .RN(n7810), 
        .QN(n1323) );
  DFFR_X1 \regfile/rx_11/data_out_reg[7]  ( .D(n3811), .CK(CLK), .RN(n6550), 
        .QN(n974) );
  DFFR_X1 \regfile/rx_11/data_out_reg[1]  ( .D(n4275), .CK(CLK), .RN(n7785), 
        .QN(n1334) );
  DFFR_X1 \regfile/rx_11/data_out_reg[0]  ( .D(n4277), .CK(CLK), .RN(n7811), 
        .QN(n1336) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[1]  ( .D(n3714), .CK(CLK), .RN(
        n6550), .Q(\Mcontrol/f_currpc[1] ), .QN(n869) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[0]  ( .D(n3888), .CK(CLK), .RN(
        n7784), .Q(\Mcontrol/f_currpc[0] ), .QN(n1042) );
  DFFR_X1 \regfile/rx_31/data_out_reg[23]  ( .D(n4134), .CK(CLK), .RN(n7813), 
        .Q(\regfile/reg_out[31][23] ), .QN(n1247) );
  DFFR_X1 \regfile/rx_31/data_out_reg[30]  ( .D(n4128), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][30] ), .QN(n1241) );
  DFFR_X1 \regfile/rx_31/data_out_reg[29]  ( .D(n4130), .CK(CLK), .RN(n7794), 
        .Q(\regfile/reg_out[31][29] ), .QN(n1243) );
  DFFR_X1 \regfile/rx_31/data_out_reg[28]  ( .D(n4131), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[31][28] ), .QN(n1244) );
  DFFR_X1 \regfile/rx_31/data_out_reg[27]  ( .D(n4132), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][27] ), .QN(n1245) );
  DFFR_X1 \regfile/rx_31/data_out_reg[31]  ( .D(n4127), .CK(CLK), .RN(n7783), 
        .Q(\regfile/reg_out[31][31] ), .QN(n1240) );
  DFFR_X1 \regfile/rx_31/data_out_reg[26]  ( .D(n4133), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[31][26] ), .QN(n1246) );
  DFFR_X1 \regfile/rx_31/data_out_reg[25]  ( .D(n3170), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][25] ), .QN(n299) );
  DFFR_X1 \regfile/rx_31/data_out_reg[24]  ( .D(n3204), .CK(CLK), .RN(n7844), 
        .Q(\regfile/reg_out[31][24] ), .QN(n351) );
  DFFR_X1 \regfile/rx_31/data_out_reg[22]  ( .D(n3243), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[31][22] ), .QN(n395) );
  DFFR_X1 \regfile/rx_31/data_out_reg[21]  ( .D(n3282), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][21] ), .QN(n431) );
  DFFR_X1 \regfile/rx_31/data_out_reg[20]  ( .D(n3321), .CK(CLK), .RN(n7758), 
        .Q(\regfile/reg_out[31][20] ), .QN(n466) );
  DFFR_X1 \regfile/rx_31/data_out_reg[19]  ( .D(n3360), .CK(CLK), .RN(n7807), 
        .Q(\regfile/reg_out[31][19] ), .QN(n501) );
  DFFR_X1 \regfile/rx_31/data_out_reg[18]  ( .D(n3399), .CK(CLK), .RN(n7797), 
        .Q(\regfile/reg_out[31][18] ), .QN(n536) );
  DFFR_X1 \regfile/rx_31/data_out_reg[17]  ( .D(n3438), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][17] ), .QN(n571) );
  DFFR_X1 \regfile/rx_31/data_out_reg[16]  ( .D(n3477), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][16] ), .QN(n606) );
  DFFR_X1 \regfile/rx_31/data_out_reg[7]  ( .D(n3833), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][7] ), .QN(n988) );
  DFFR_X1 \regfile/rx_31/data_out_reg[1]  ( .D(n4135), .CK(CLK), .RN(n7763), 
        .Q(\regfile/reg_out[31][1] ), .QN(n1248) );
  DFFR_X1 \regfile/rx_31/data_out_reg[0]  ( .D(n4137), .CK(CLK), .RN(n7844), 
        .Q(\regfile/reg_out[31][0] ), .QN(n1250) );
  DFFR_X1 \regfile/rx_31/data_out_reg[14]  ( .D(n4136), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][14] ), .QN(n1249) );
  DFFR_X1 \regfile/rx_31/data_out_reg[13]  ( .D(n3677), .CK(CLK), .RN(n7849), 
        .Q(\regfile/reg_out[31][13] ), .QN(n810) );
  DFFR_X1 \regfile/rx_31/data_out_reg[12]  ( .D(n3638), .CK(CLK), .RN(n7743), 
        .Q(\regfile/reg_out[31][12] ), .QN(n772) );
  DFFR_X1 \regfile/rx_31/data_out_reg[11]  ( .D(n3599), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][11] ), .QN(n734) );
  DFFR_X1 \regfile/rx_31/data_out_reg[10]  ( .D(n3560), .CK(CLK), .RN(n7848), 
        .Q(\regfile/reg_out[31][10] ), .QN(n696) );
  DFFR_X1 \regfile/rx_31/data_out_reg[6]  ( .D(n3791), .CK(CLK), .RN(n7845), 
        .Q(\regfile/reg_out[31][6] ), .QN(n949) );
  DFFR_X1 \regfile/rx_31/data_out_reg[5]  ( .D(n3749), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][5] ), .QN(n905) );
  DFFR_X1 \regfile/rx_31/data_out_reg[4]  ( .D(n4125), .CK(CLK), .RN(n7847), 
        .Q(\regfile/reg_out[31][4] ), .QN(n1238) );
  DFFR_X1 \regfile/rx_31/data_out_reg[3]  ( .D(n4126), .CK(CLK), .RN(n7851), 
        .Q(\regfile/reg_out[31][3] ), .QN(n1239) );
  DFFR_X1 \regfile/rx_31/data_out_reg[2]  ( .D(n4129), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][2] ), .QN(n1242) );
  DFFR_X1 \regfile/rx_31/data_out_reg[15]  ( .D(n3519), .CK(CLK), .RN(n7846), 
        .Q(\regfile/reg_out[31][15] ), .QN(n647) );
  DFFR_X1 \regfile/rx_31/data_out_reg[9]  ( .D(n3875), .CK(CLK), .RN(n7823), 
        .Q(\regfile/reg_out[31][9] ), .QN(n1027) );
  DFFR_X1 \regfile/rx_31/data_out_reg[8]  ( .D(n4124), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[31][8] ), .QN(n1237) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[18]  ( .D(n3373), .CK(CLK), 
        .RN(n7845), .Q(\Mcontrol/f_currpc[18] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[21]  ( .D(n6969), .CK(CLK), 
        .RN(n7742), .Q(\Mcontrol/f_currpc[21] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[17]  ( .D(n3412), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/f_currpc[17] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[15]  ( .D(n3490), .CK(CLK), 
        .RN(n7851), .Q(\Mcontrol/f_currpc[15] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[14]  ( .D(n3532), .CK(CLK), 
        .RN(n7738), .Q(\Mcontrol/f_currpc[14] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[13]  ( .D(n3651), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/f_currpc[13] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[12]  ( .D(n3612), .CK(CLK), 
        .RN(n7807), .Q(\Mcontrol/f_currpc[12] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[16]  ( .D(n3451), .CK(CLK), 
        .RN(n7825), .Q(\Mcontrol/f_currpc[16] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[19]  ( .D(n3334), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/f_currpc[19] ) );
  DFFR_X1 \regfile/rx_3/data_out_reg[15]  ( .D(n3520), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[3][15] ), .QN(n648) );
  DFFR_X1 \regfile/rx_3/data_out_reg[23]  ( .D(n4330), .CK(CLK), .RN(n7852), 
        .Q(\regfile/reg_out[3][23] ), .QN(n1375) );
  DFFR_X1 \regfile/rx_3/data_out_reg[30]  ( .D(n4324), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][30] ), .QN(n1369) );
  DFFR_X1 \regfile/rx_3/data_out_reg[29]  ( .D(n4326), .CK(CLK), .RN(n7808), 
        .Q(\regfile/reg_out[3][29] ), .QN(n1371) );
  DFFR_X1 \regfile/rx_3/data_out_reg[28]  ( .D(n4327), .CK(CLK), .RN(n7820), 
        .Q(\regfile/reg_out[3][28] ), .QN(n1372) );
  DFFR_X1 \regfile/rx_3/data_out_reg[27]  ( .D(n4328), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][27] ), .QN(n1373) );
  DFFR_X1 \regfile/rx_3/data_out_reg[31]  ( .D(n4323), .CK(CLK), .RN(n7789), 
        .Q(\regfile/reg_out[3][31] ), .QN(n1368) );
  DFFR_X1 \regfile/rx_3/data_out_reg[26]  ( .D(n4329), .CK(CLK), .RN(n7717), 
        .Q(\regfile/reg_out[3][26] ), .QN(n1374) );
  DFFR_X1 \regfile/rx_3/data_out_reg[25]  ( .D(n3171), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][25] ), .QN(n302) );
  DFFR_X1 \regfile/rx_3/data_out_reg[24]  ( .D(n3205), .CK(CLK), .RN(n7788), 
        .Q(\regfile/reg_out[3][24] ), .QN(n352) );
  DFFR_X1 \regfile/rx_3/data_out_reg[22]  ( .D(n3244), .CK(CLK), .RN(n7729), 
        .Q(\regfile/reg_out[3][22] ), .QN(n396) );
  DFFR_X1 \regfile/rx_3/data_out_reg[21]  ( .D(n3283), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][21] ), .QN(n432) );
  DFFR_X1 \regfile/rx_3/data_out_reg[20]  ( .D(n3322), .CK(CLK), .RN(n7787), 
        .Q(\regfile/reg_out[3][20] ), .QN(n467) );
  DFFR_X1 \regfile/rx_3/data_out_reg[19]  ( .D(n3361), .CK(CLK), .RN(n7723), 
        .Q(\regfile/reg_out[3][19] ), .QN(n502) );
  DFFR_X1 \regfile/rx_3/data_out_reg[18]  ( .D(n3400), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][18] ), .QN(n537) );
  DFFR_X1 \regfile/rx_3/data_out_reg[17]  ( .D(n3439), .CK(CLK), .RN(n7786), 
        .Q(\regfile/reg_out[3][17] ), .QN(n572) );
  DFFR_X1 \regfile/rx_3/data_out_reg[16]  ( .D(n3478), .CK(CLK), .RN(n7745), 
        .Q(\regfile/reg_out[3][16] ), .QN(n607) );
  DFFR_X1 \regfile/rx_3/data_out_reg[7]  ( .D(n3834), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][7] ), .QN(n989) );
  DFFR_X1 \regfile/rx_3/data_out_reg[1]  ( .D(n4331), .CK(CLK), .RN(n7785), 
        .Q(\regfile/reg_out[3][1] ), .QN(n1376) );
  DFFR_X1 \regfile/rx_3/data_out_reg[0]  ( .D(n4333), .CK(CLK), .RN(n7741), 
        .Q(\regfile/reg_out[3][0] ), .QN(n1378) );
  DFFR_X1 \regfile/rx_3/data_out_reg[14]  ( .D(n4332), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][14] ), .QN(n1377) );
  DFFR_X1 \regfile/rx_3/data_out_reg[13]  ( .D(n3678), .CK(CLK), .RN(n7784), 
        .Q(\regfile/reg_out[3][13] ), .QN(n811) );
  DFFR_X1 \regfile/rx_3/data_out_reg[12]  ( .D(n3639), .CK(CLK), .RN(n7802), 
        .Q(\regfile/reg_out[3][12] ), .QN(n773) );
  DFFR_X1 \regfile/rx_3/data_out_reg[11]  ( .D(n3600), .CK(CLK), .RN(n7851), 
        .Q(\regfile/reg_out[3][11] ), .QN(n735) );
  DFFR_X1 \regfile/rx_3/data_out_reg[10]  ( .D(n3561), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][10] ), .QN(n697) );
  DFFR_X1 \regfile/rx_3/data_out_reg[6]  ( .D(n3792), .CK(CLK), .RN(n7804), 
        .Q(\regfile/reg_out[3][6] ), .QN(n950) );
  DFFR_X1 \regfile/rx_3/data_out_reg[5]  ( .D(n3750), .CK(CLK), .RN(n7758), 
        .Q(\regfile/reg_out[3][5] ), .QN(n906) );
  DFFR_X1 \regfile/rx_3/data_out_reg[4]  ( .D(n4321), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][4] ), .QN(n1366) );
  DFFR_X1 \regfile/rx_3/data_out_reg[3]  ( .D(n4322), .CK(CLK), .RN(n7852), 
        .Q(\regfile/reg_out[3][3] ), .QN(n1367) );
  DFFR_X1 \regfile/rx_3/data_out_reg[2]  ( .D(n4325), .CK(CLK), .RN(n7776), 
        .Q(\regfile/reg_out[3][2] ), .QN(n1370) );
  DFFR_X1 \regfile/rx_3/data_out_reg[9]  ( .D(n3876), .CK(CLK), .RN(n6550), 
        .Q(\regfile/reg_out[3][9] ), .QN(n1028) );
  DFFR_X1 \regfile/rx_3/data_out_reg[8]  ( .D(n4320), .CK(CLK), .RN(n7805), 
        .Q(\regfile/reg_out[3][8] ), .QN(n1365) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[23]  ( .D(n7565), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/f_currpc[23] ) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[15]  ( .D(n3486), .CK(CLK), .RN(
        n7761), .Q(epc[15]), .QN(n615) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[14]  ( .D(n3528), .CK(CLK), .RN(
        n6550), .Q(epc[14]), .QN(n662) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[13]  ( .D(n3647), .CK(CLK), .RN(
        n7808), .Q(epc[13]), .QN(n783) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[12]  ( .D(n3608), .CK(CLK), .RN(
        n7787), .Q(epc[12]), .QN(n745) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[11]  ( .D(n3569), .CK(CLK), .RN(
        n6550), .Q(epc[11]), .QN(n707) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[10]  ( .D(n3535), .CK(CLK), .RN(
        n6550), .Q(epc[10]), .QN(n677) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[9]  ( .D(n3842), .CK(CLK), .RN(
        n7807), .Q(epc[9]), .QN(n999) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[8]  ( .D(n3686), .CK(CLK), .RN(
        n7836), .Q(epc[8]), .QN(n821) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[7]  ( .D(n3800), .CK(CLK), .RN(
        n6550), .Q(epc[7]), .QN(n960) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[6]  ( .D(n3758), .CK(CLK), .RN(
        n7758), .Q(epc[6]), .QN(n921) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[5]  ( .D(n3715), .CK(CLK), .RN(
        n7810), .Q(epc[5]), .QN(n873) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[4]  ( .D(n3692), .CK(CLK), .RN(
        n7750), .Q(epc[4]), .QN(n832) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[3]  ( .D(n3698), .CK(CLK), .RN(
        n7790), .Q(epc[3]), .QN(n843) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[2]  ( .D(n3704), .CK(CLK), .RN(
        n6550), .Q(epc[2]), .QN(n854) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[1]  ( .D(n3710), .CK(CLK), .RN(
        n7821), .Q(epc[1]), .QN(n865) );
  DFFR_X1 \Scc_coproc/EPC_REG/data_out_reg[0]  ( .D(n3889), .CK(CLK), .RN(
        n7811), .Q(epc[0]), .QN(n1045) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[22]  ( .D(n6988), .CK(CLK), 
        .RN(n6550), .Q(\Mcontrol/f_currpc[22] ) );
  DFFR_X1 \Mcontrol/Program_counter/out_pc_reg[20]  ( .D(n3295), .CK(CLK), 
        .RN(n7773), .Q(\Mcontrol/f_currpc[20] ) );
  DFFS_X2 \Mcontrol/ir_xm/out_mem_command_reg[MR]  ( .D(n4411), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .Q(\m_mem_command[MR] ), .QN(n5745) );
  DFFS_X2 \Mcontrol/ir_xm/out_serve_exception_reg  ( .D(n4425), .CK(CLK), .SN(
        \Mcontrol/int_reset ), .QN(n6102) );
  CLKBUF_X1 U5456 ( .A(n6550), .Z(n7852) );
  CLKBUF_X1 U5457 ( .A(n7852), .Z(n7851) );
  CLKBUF_X1 U5458 ( .A(n7845), .Z(n7844) );
  INV_X1 U5459 ( .A(n6102), .ZN(net59736) );
  INV_X1 U5460 ( .A(n6102), .ZN(n6940) );
  OR3_X2 U5461 ( .A1(n6102), .A2(n6932), .A3(net59612), .ZN(n1557) );
  CLKBUF_X1 U5462 ( .A(D_DATA_INBUS[6]), .Z(n6514) );
  INV_X1 U5463 ( .A(n5856), .ZN(n6515) );
  CLKBUF_X1 U5464 ( .A(D_DATA_INBUS[5]), .Z(n6516) );
  AOI222_X1 U5465 ( .A1(n6102), .A2(n6516), .B1(
        \Mcontrol/Nextpc_decoding/Bta [5]), .B2(n1560), .C1(jar_in[5]), .C2(
        net57184), .ZN(n2576) );
  INV_X1 U5466 ( .A(n5831), .ZN(n6517) );
  CLKBUF_X1 U5467 ( .A(D_DATA_INBUS[4]), .Z(n6518) );
  INV_X1 U5468 ( .A(n5821), .ZN(n6519) );
  CLKBUF_X1 U5469 ( .A(D_DATA_INBUS[3]), .Z(n6520) );
  INV_X1 U5470 ( .A(n5811), .ZN(n6521) );
  CLKBUF_X1 U5471 ( .A(D_DATA_INBUS[2]), .Z(n6522) );
  INV_X1 U5472 ( .A(n5799), .ZN(n6523) );
  CLKBUF_X1 U5473 ( .A(D_DATA_INBUS[21]), .Z(n6524) );
  NAND2_X1 U5474 ( .A1(n6102), .A2(n6524), .ZN(n7373) );
  CLKBUF_X1 U5475 ( .A(D_DATA_INBUS[22]), .Z(n6525) );
  NAND2_X1 U5476 ( .A1(n6525), .A2(n6102), .ZN(n6936) );
  CLKBUF_X1 U5477 ( .A(D_DATA_INBUS[20]), .Z(n6526) );
  NAND2_X1 U5478 ( .A1(n6102), .A2(n6526), .ZN(n7346) );
  CLKBUF_X1 U5479 ( .A(D_DATA_INBUS[24]), .Z(n6527) );
  CLKBUF_X1 U5480 ( .A(D_DATA_INBUS[19]), .Z(n6528) );
  CLKBUF_X1 U5481 ( .A(D_DATA_INBUS[25]), .Z(n6529) );
  CLKBUF_X1 U5482 ( .A(D_DATA_INBUS[18]), .Z(n6530) );
  AND2_X1 U5483 ( .A1(n6102), .A2(n6530), .ZN(n7243) );
  CLKBUF_X1 U5484 ( .A(D_DATA_INBUS[26]), .Z(n6531) );
  CLKBUF_X1 U5485 ( .A(D_DATA_INBUS[17]), .Z(n6532) );
  CLKBUF_X1 U5486 ( .A(D_DATA_INBUS[27]), .Z(n6533) );
  CLKBUF_X1 U5487 ( .A(D_DATA_INBUS[16]), .Z(n6534) );
  CLKBUF_X1 U5488 ( .A(D_DATA_INBUS[28]), .Z(n6535) );
  CLKBUF_X1 U5489 ( .A(D_DATA_INBUS[9]), .Z(n6536) );
  CLKBUF_X1 U5490 ( .A(D_DATA_INBUS[29]), .Z(n6537) );
  CLKBUF_X1 U5491 ( .A(D_DATA_INBUS[8]), .Z(n6538) );
  CLKBUF_X1 U5492 ( .A(D_DATA_INBUS[30]), .Z(n6539) );
  CLKBUF_X1 U5493 ( .A(D_DATA_INBUS[7]), .Z(n6540) );
  CLKBUF_X1 U5494 ( .A(D_DATA_INBUS[31]), .Z(n6541) );
  CLKBUF_X1 U5495 ( .A(D_DATA_INBUS[1]), .Z(n6542) );
  CLKBUF_X1 U5496 ( .A(D_NREADY), .Z(n6543) );
  AND2_X1 U5497 ( .A1(\Mcontrol/N34 ), .A2(n6543), .ZN(I_BUSY) );
  INV_X1 U5498 ( .A(n6543), .ZN(n7215) );
  CLKBUF_X1 U5499 ( .A(D_DATA_INBUS[23]), .Z(n6544) );
  NAND2_X1 U5500 ( .A1(n6102), .A2(n6544), .ZN(n7012) );
  CLKBUF_X1 U5501 ( .A(I_NREADY), .Z(n6545) );
  NAND3_X1 U5502 ( .A1(n6545), .A2(n6543), .A3(\Mcontrol/N25 ), .ZN(n1655) );
  INV_X1 U5503 ( .A(n6545), .ZN(n7214) );
  CLKBUF_X1 U5504 ( .A(D_DATA_INBUS[15]), .Z(n6546) );
  CLKBUF_X1 U5505 ( .A(reboot), .Z(n6547) );
  CLKBUF_X1 U5506 ( .A(freeze), .Z(D_BUSY) );
  NAND2_X2 U5507 ( .A1(n6543), .A2(D_BUSY), .ZN(n220) );
  AND2_X1 U5508 ( .A1(\Mcontrol/stall_decode ), .A2(D_BUSY), .ZN(
        \Mcontrol/N25 ) );
  AND2_X1 U5509 ( .A1(\Mcontrol/stall_decode ), .A2(D_BUSY), .ZN(
        \Mcontrol/N34 ) );
  INV_X2 U5510 ( .A(reset), .ZN(n6549) );
  INV_X16 U5511 ( .A(n6549), .ZN(n6550) );
  INV_X1 U5512 ( .A(n621), .ZN(n6551) );
  INV_X1 U5513 ( .A(n7488), .ZN(n7161) );
  INV_X1 U5514 ( .A(n7488), .ZN(n7147) );
  OR2_X1 U5515 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(
        \Mcontrol/Nextpc_decoding/N323 ), .ZN(\Mcontrol/Nextpc_decoding/N324 )
         );
  OR2_X1 U5516 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(
        \Mcontrol/Nextpc_decoding/N311 ), .ZN(\Mcontrol/Nextpc_decoding/N312 )
         );
  OR2_X1 U5517 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(
        \Mcontrol/Nextpc_decoding/N299 ), .ZN(\Mcontrol/Nextpc_decoding/N300 )
         );
  OR2_X1 U5518 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(
        \Mcontrol/Nextpc_decoding/N287 ), .ZN(\Mcontrol/Nextpc_decoding/N288 )
         );
  INV_X1 U5519 ( .A(\Mcontrol/d_jump_type[0] ), .ZN(n6929) );
  OR2_X1 U5520 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(
        \Mcontrol/Nextpc_decoding/N169 ), .ZN(\Mcontrol/Nextpc_decoding/N170 )
         );
  INV_X1 U5521 ( .A(\Mcontrol/d_jump_type[0] ), .ZN(
        \Mcontrol/Nextpc_decoding/N173 ) );
  OR2_X1 U5522 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(\Mcontrol/st_logic/N62 ), 
        .ZN(\Mcontrol/st_logic/N63 ) );
  OR2_X1 U5523 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(\Mcontrol/st_logic/N100 ), 
        .ZN(\Mcontrol/st_logic/N101 ) );
  OR2_X1 U5524 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(\Mcontrol/st_logic/N87 ), 
        .ZN(\Mcontrol/st_logic/N88 ) );
  OR2_X1 U5525 ( .A1(\Mcontrol/d_jump_type[0] ), .A2(\Mcontrol/st_logic/N75 ), 
        .ZN(\Mcontrol/st_logic/N76 ) );
  INV_X1 U5526 ( .A(\Mcontrol/d_jump_type[0] ), .ZN(\Mcontrol/st_logic/N65 )
         );
  INV_X1 U5527 ( .A(net55890), .ZN(net57331) );
  INV_X1 U5528 ( .A(net55890), .ZN(net57757) );
  INV_X1 U5529 ( .A(net55890), .ZN(net57465) );
  INV_X1 U5530 ( .A(net55890), .ZN(net57255) );
  OR3_X1 U5531 ( .A1(\regfile/N391 ), .A2(net55890), .A3(n1108), .ZN(n7407) );
  AOI221_X1 U5532 ( .B1(\d_chk/N7 ), .B2(n6447), .C1(n7131), .C2(n6474), .A(
        \d_chk/N10 ), .ZN(n6494) );
  NOR2_X2 U5533 ( .A1(n5505), .A2(n4508), .ZN(n6447) );
  INV_X2 U5534 ( .A(n1661), .ZN(n192) );
  INV_X2 U5535 ( .A(n1658), .ZN(n197) );
  OR3_X1 U5536 ( .A1(\Mpath/the_shift/N115 ), .A2(\Mpath/the_shift/N118 ), 
        .A3(n1914), .ZN(n6552) );
  INV_X2 U5537 ( .A(n6552), .ZN(n6553) );
  AND2_X2 U5538 ( .A1(n1676), .A2(n184), .ZN(n195) );
  AND2_X4 U5539 ( .A1(n6503), .A2(\Mpath/the_shift/N107 ), .ZN(n1703) );
  NAND2_X2 U5540 ( .A1(n184), .A2(n183), .ZN(n53) );
  NAND2_X2 U5541 ( .A1(n183), .A2(n185), .ZN(n51) );
  INV_X2 U5542 ( .A(n5769), .ZN(n1926) );
  NAND3_X2 U5543 ( .A1(n1675), .A2(n322), .A3(\Mpath/N197 ), .ZN(n323) );
  CLKBUF_X1 U5544 ( .A(n232), .Z(n6554) );
  AND2_X2 U5545 ( .A1(n182), .A2(n183), .ZN(n55) );
  NAND3_X1 U5546 ( .A1(net55862), .A2(\Mcontrol/st_logic/N47 ), .A3(
        byp_controlA[2]), .ZN(n6555) );
  INV_X2 U5547 ( .A(n6555), .ZN(n6556) );
  OR3_X1 U5548 ( .A1(\regfile/N286 ), .A2(net55894), .A3(n1251), .ZN(n6557) );
  INV_X1 U5549 ( .A(n6557), .ZN(n6558) );
  INV_X1 U5550 ( .A(n6557), .ZN(n6559) );
  INV_X1 U5551 ( .A(n6558), .ZN(n303) );
  INV_X2 U5552 ( .A(n624), .ZN(n119) );
  INV_X2 U5553 ( .A(n671), .ZN(n123) );
  INV_X2 U5554 ( .A(n588), .ZN(n115) );
  INV_X2 U5555 ( .A(n792), .ZN(n127) );
  INV_X2 U5556 ( .A(n553), .ZN(n111) );
  INV_X2 U5557 ( .A(n754), .ZN(n131) );
  INV_X2 U5558 ( .A(n518), .ZN(n107) );
  INV_X2 U5559 ( .A(n716), .ZN(n135) );
  INV_X2 U5560 ( .A(n483), .ZN(n103) );
  INV_X2 U5561 ( .A(n675), .ZN(n139) );
  INV_X2 U5562 ( .A(n448), .ZN(n99) );
  INV_X2 U5563 ( .A(n1008), .ZN(n143) );
  INV_X2 U5564 ( .A(n413), .ZN(n95) );
  INV_X2 U5565 ( .A(n830), .ZN(n147) );
  INV_X2 U5566 ( .A(n377), .ZN(n91) );
  INV_X2 U5567 ( .A(n969), .ZN(n151) );
  INV_X2 U5568 ( .A(n1404), .ZN(n87) );
  INV_X2 U5569 ( .A(n930), .ZN(n155) );
  INV_X2 U5570 ( .A(n328), .ZN(n83) );
  INV_X2 U5571 ( .A(n882), .ZN(n159) );
  INV_X2 U5572 ( .A(n230), .ZN(n79) );
  INV_X2 U5573 ( .A(n841), .ZN(n163) );
  INV_X2 U5574 ( .A(n222), .ZN(n75) );
  INV_X2 U5575 ( .A(n216), .ZN(n71) );
  INV_X2 U5576 ( .A(n852), .ZN(n167) );
  INV_X2 U5577 ( .A(n863), .ZN(n171) );
  INV_X2 U5578 ( .A(n207), .ZN(n67) );
  INV_X2 U5579 ( .A(n202), .ZN(n63) );
  INV_X2 U5580 ( .A(n1406), .ZN(n175) );
  INV_X2 U5581 ( .A(n1668), .ZN(n179) );
  INV_X2 U5582 ( .A(n196), .ZN(n59) );
  NAND2_X2 U5583 ( .A1(net55840), .A2(n187), .ZN(n57) );
  INV_X2 U5584 ( .A(n1390), .ZN(n52) );
  OR2_X2 U5585 ( .A1(exe_outsel[0]), .A2(\Mpath/N193 ), .ZN(n322) );
  OR2_X1 U5586 ( .A1(\Mpath/N187 ), .A2(exe_outsel[2]), .ZN(\Mpath/N193 ) );
  NOR2_X4 U5587 ( .A1(n2877), .A2(n2878), .ZN(n1563) );
  AOI222_X1 U5588 ( .A1(\Mcontrol/Nextpc_decoding/Bta [0]), .A2(n1560), .B1(
        epc[0]), .B2(n1562), .C1(n1563), .C2(net56595), .ZN(n1566) );
  INV_X1 U5589 ( .A(n1563), .ZN(n6941) );
  NOR2_X4 U5590 ( .A1(n1051), .A2(n1049), .ZN(n361) );
  CLKBUF_X2 U5591 ( .A(n235), .Z(n6560) );
  AND2_X4 U5592 ( .A1(n7822), .A2(n6547), .ZN(\Mcontrol/int_reset ) );
  INV_X1 U5593 ( .A(n7078), .ZN(n6890) );
  INV_X1 U5594 ( .A(n6890), .ZN(n6891) );
  INV_X1 U5595 ( .A(n5765), .ZN(n6892) );
  INV_X1 U5596 ( .A(n2523), .ZN(n6893) );
  NOR4_X2 U5597 ( .A1(n2515), .A2(n2516), .A3(n2517), .A4(n2518), .ZN(n2514)
         );
  NAND2_X1 U5598 ( .A1(n6910), .A2(n6911), .ZN(
        \Mcontrol/Operation_decoding32/N1963 ) );
  CLKBUF_X1 U5599 ( .A(n7886), .Z(I_ADDR_OUTBUS[2]) );
  INV_X1 U5600 ( .A(n267), .ZN(n6895) );
  INV_X1 U5601 ( .A(n267), .ZN(n6896) );
  INV_X1 U5602 ( .A(n267), .ZN(n6897) );
  INV_X4 U5603 ( .A(n265), .ZN(n6898) );
  NOR3_X1 U5604 ( .A1(\regfile/N273 ), .A2(net55894), .A3(n1252), .ZN(n265) );
  INV_X1 U5605 ( .A(n265), .ZN(n267) );
  NOR2_X2 U5606 ( .A1(\Mcontrol/Operation_decoding32/N2003 ), .A2(n7221), .ZN(
        n7273) );
  OAI22_X1 U5607 ( .A1(\Mcontrol/Nextpc_decoding/N31 ), .A2(n6404), .B1(n6405), 
        .B2(\Mcontrol/Nextpc_decoding/N313 ), .ZN(n6401) );
  NOR4_X2 U5608 ( .A1(n2619), .A2(n2620), .A3(n2621), .A4(n2622), .ZN(n2618)
         );
  AND2_X1 U5609 ( .A1(n6899), .A2(\Mcontrol/st_logic/N88 ), .ZN(n7188) );
  NOR2_X1 U5610 ( .A1(\Mcontrol/st_logic/N77 ), .A2(\Mcontrol/st_logic/N83 ), 
        .ZN(n6899) );
  AND2_X4 U5611 ( .A1(n6037), .A2(n6034), .ZN(n6033) );
  NOR2_X1 U5612 ( .A1(n7595), .A2(n7594), .ZN(\Mcontrol/Nextpc_decoding/N36 )
         );
  OR2_X1 U5613 ( .A1(\Mcontrol/st_logic/N65 ), .A2(\Mcontrol/st_logic/N107 ), 
        .ZN(\Mcontrol/st_logic/N108 ) );
  OR2_X1 U5614 ( .A1(\Mcontrol/st_logic/N65 ), .A2(\Mcontrol/st_logic/N69 ), 
        .ZN(\Mcontrol/st_logic/N70 ) );
  OR2_X1 U5615 ( .A1(\Mcontrol/st_logic/N65 ), .A2(\Mcontrol/st_logic/N94 ), 
        .ZN(\Mcontrol/st_logic/N95 ) );
  OAI21_X2 U5616 ( .B1(n6069), .B2(n7309), .A(n7585), .ZN(n2502) );
  INV_X1 U5617 ( .A(n7602), .ZN(n6900) );
  NAND2_X1 U5618 ( .A1(n6901), .A2(n6902), .ZN(n7237) );
  AND2_X1 U5619 ( .A1(n7555), .A2(n7554), .ZN(n6901) );
  NOR2_X2 U5620 ( .A1(n6981), .A2(n6900), .ZN(n6902) );
  NOR2_X2 U5621 ( .A1(branch_rega[18]), .A2(\Mcontrol/Nextpc_decoding/N198 ), 
        .ZN(n7554) );
  AND3_X4 U5622 ( .A1(rs2_addr[1]), .A2(rs2_addr[0]), .A3(n6017), .ZN(n5752)
         );
  NAND2_X1 U5623 ( .A1(n7101), .A2(n7103), .ZN(n6903) );
  NAND2_X1 U5624 ( .A1(n7102), .A2(n6904), .ZN(n6969) );
  INV_X1 U5625 ( .A(n6903), .ZN(n6904) );
  NAND2_X1 U5626 ( .A1(n7704), .A2(n7264), .ZN(n7265) );
  NOR4_X1 U5627 ( .A1(n2798), .A2(n2799), .A3(n2800), .A4(n2801), .ZN(n2797)
         );
  NOR2_X1 U5628 ( .A1(n7280), .A2(n6989), .ZN(n6496) );
  BUF_X1 U5629 ( .A(\Mpath/the_alu/diff[31] ), .Z(n7658) );
  NOR2_X1 U5630 ( .A1(n7656), .A2(branch_rega[26]), .ZN(n7480) );
  OR2_X1 U5631 ( .A1(\Mcontrol/Nextpc_decoding/N221 ), .A2(branch_rega[28]), 
        .ZN(n7281) );
  INV_X2 U5632 ( .A(n7213), .ZN(n2477) );
  INV_X2 U5633 ( .A(n5754), .ZN(n6905) );
  INV_X4 U5634 ( .A(n6905), .ZN(n6906) );
  NAND2_X4 U5635 ( .A1(n1379), .A2(n1221), .ZN(n1252) );
  NAND2_X2 U5636 ( .A1(\Mcontrol/Operation_decoding32/N2084 ), .A2(net57388), 
        .ZN(net57268) );
  NAND2_X2 U5637 ( .A1(net56922), .A2(n7399), .ZN(net57388) );
  OR2_X1 U5638 ( .A1(rs2_addr[3]), .A2(rs2_addr[4]), .ZN(\regfile/N265 ) );
  OAI222_X4 U5639 ( .A1(n5623), .A2(n5526), .B1(n7486), .B2(n2510), .C1(n5621), 
        .C2(n5522), .ZN(branch_rega[9]) );
  OR2_X2 U5640 ( .A1(n7475), .A2(branch_rega[10]), .ZN(n7474) );
  NAND2_X1 U5641 ( .A1(n6431), .A2(n7327), .ZN(n5653) );
  NAND2_X2 U5642 ( .A1(n7705), .A2(\Mcontrol/Operation_decoding32/N1871 ), 
        .ZN(n7675) );
  INV_X2 U5643 ( .A(n7516), .ZN(n7519) );
  NOR2_X1 U5644 ( .A1(n7032), .A2(n7234), .ZN(n7452) );
  NOR4_X2 U5645 ( .A1(n2532), .A2(n2533), .A3(n2534), .A4(n2535), .ZN(n2531)
         );
  INV_X1 U5646 ( .A(n7256), .ZN(n6907) );
  NAND2_X1 U5647 ( .A1(n6908), .A2(n6909), .ZN(
        \Mcontrol/Operation_decoding32/N1944 ) );
  AND2_X1 U5648 ( .A1(n7455), .A2(n7431), .ZN(n6908) );
  NOR2_X1 U5649 ( .A1(\Mcontrol/d_instr [27]), .A2(n6907), .ZN(n6909) );
  NOR2_X1 U5650 ( .A1(n7063), .A2(n7066), .ZN(n6910) );
  AND2_X1 U5651 ( .A1(n7079), .A2(n7569), .ZN(n6911) );
  NOR2_X1 U5652 ( .A1(n7341), .A2(n7339), .ZN(n6912) );
  NOR2_X1 U5653 ( .A1(n7340), .A2(n6913), .ZN(n2715) );
  INV_X1 U5654 ( .A(n6912), .ZN(n6913) );
  INV_X2 U5655 ( .A(branch_rega[4]), .ZN(n7651) );
  INV_X2 U5656 ( .A(branch_rega[4]), .ZN(n7674) );
  OR2_X2 U5657 ( .A1(branch_rega[29]), .A2(\Mcontrol/Nextpc_decoding/N252 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N188 ) );
  NAND2_X1 U5658 ( .A1(rd_addr[1]), .A2(n1222), .ZN(n1107) );
  NAND2_X4 U5659 ( .A1(n1379), .A2(rd_addr[1]), .ZN(n1251) );
  INV_X4 U5660 ( .A(n7688), .ZN(n5646) );
  NOR2_X1 U5661 ( .A1(n7208), .A2(n7183), .ZN(n7213) );
  INV_X1 U5662 ( .A(\d_chk/N12 ), .ZN(\d_chk/N7 ) );
  AND2_X4 U5663 ( .A1(n6028), .A2(n6037), .ZN(n1937) );
  AND2_X4 U5664 ( .A1(n6030), .A2(n6020), .ZN(n6028) );
  OR2_X2 U5665 ( .A1(n2880), .A2(net57323), .ZN(n2509) );
  NOR2_X4 U5666 ( .A1(net57268), .A2(n7548), .ZN(n1434) );
  INV_X1 U5667 ( .A(branch_rega[5]), .ZN(n7660) );
  INV_X1 U5668 ( .A(n6974), .ZN(n6914) );
  NOR2_X1 U5669 ( .A1(n6915), .A2(n6973), .ZN(n7595) );
  NAND2_X1 U5670 ( .A1(n7179), .A2(n6914), .ZN(n6915) );
  OR2_X2 U5671 ( .A1(branch_rega[29]), .A2(\Mcontrol/Nextpc_decoding/N252 ), 
        .ZN(\Mcontrol/Nextpc_decoding/N253 ) );
  OAI21_X1 U5672 ( .B1(n2461), .B2(\Mcontrol/Operation_decoding32/N1901 ), .A(
        n2462), .ZN(break_code[0]) );
  CLKBUF_X1 U5673 ( .A(break_code[0]), .Z(net56595) );
  NAND2_X1 U5674 ( .A1(n6080), .A2(n6922), .ZN(n2462) );
  INV_X1 U5675 ( .A(n6921), .ZN(n6922) );
  NAND2_X1 U5676 ( .A1(net57253), .A2(\Mcontrol/d_instr[6] ), .ZN(n6921) );
  INV_X2 U5677 ( .A(n6120), .ZN(\Mcontrol/d_instr[6] ) );
  AND2_X2 U5678 ( .A1(n6916), .A2(n6917), .ZN(n2461) );
  OR2_X1 U5679 ( .A1(n2461), .A2(n5519), .ZN(n2458) );
  NAND2_X1 U5680 ( .A1(n5521), .A2(net57268), .ZN(n6917) );
  INV_X1 U5681 ( .A(n6918), .ZN(n5521) );
  INV_X1 U5682 ( .A(net57386), .ZN(n6918) );
  NAND2_X1 U5683 ( .A1(n6079), .A2(n1482), .ZN(n6916) );
  NOR2_X1 U5684 ( .A1(n6924), .A2(n6919), .ZN(n1482) );
  INV_X1 U5685 ( .A(net57386), .ZN(n6919) );
  INV_X1 U5686 ( .A(n6919), .ZN(net58547) );
  NAND2_X1 U5687 ( .A1(n6925), .A2(net57388), .ZN(n6924) );
  INV_X1 U5688 ( .A(n6923), .ZN(n6925) );
  CLKBUF_X1 U5689 ( .A(n6925), .Z(net57954) );
  NOR2_X1 U5690 ( .A1(net58300), .A2(net57313), .ZN(n6923) );
  AOI21_X2 U5691 ( .B1(n6101), .B2(n6920), .A(net56668), .ZN(n6100) );
  NOR2_X1 U5692 ( .A1(net56765), .A2(net58543), .ZN(n6920) );
  INV_X2 U5693 ( .A(\Mcontrol/Nextpc_decoding/N298 ), .ZN(n6928) );
  INV_X1 U5694 ( .A(\Mcontrol/d_jump_type[1] ), .ZN(n6939) );
  INV_X1 U5695 ( .A(n6939), .ZN(n6953) );
  CLKBUF_X1 U5696 ( .A(branch_rega[22]), .Z(n6952) );
  CLKBUF_X1 U5697 ( .A(net55921), .Z(n6951) );
  BUF_X1 U5698 ( .A(n1560), .Z(net58826) );
  OR2_X2 U5699 ( .A1(branch_rega[9]), .A2(branch_rega[8]), .ZN(n7556) );
  INV_X4 U5700 ( .A(n7675), .ZN(rs1_addr[0]) );
  INV_X8 U5701 ( .A(n7120), .ZN(n282) );
  OAI211_X1 U5702 ( .C1(n2627), .C2(n1557), .A(n2628), .B(n2629), .ZN(n7886)
         );
  INV_X4 U5703 ( .A(branch_rega[2]), .ZN(n7685) );
  CLKBUF_X1 U5704 ( .A(n7009), .Z(n6954) );
  INV_X2 U5705 ( .A(\Mpath/out_regB[8] ), .ZN(n7613) );
  NOR2_X1 U5706 ( .A1(\Mcontrol/Operation_decoding32/N1923 ), .A2(n6955), .ZN(
        n7541) );
  OR2_X2 U5707 ( .A1(n7145), .A2(n6956), .ZN(n6955) );
  INV_X1 U5708 ( .A(n7256), .ZN(n6956) );
  NOR2_X2 U5709 ( .A1(\Mcontrol/Operation_decoding32/N1924 ), .A2(n7302), .ZN(
        \Mcontrol/Operation_decoding32/N1928 ) );
  OR2_X2 U5710 ( .A1(n7098), .A2(n7425), .ZN(
        \Mcontrol/Operation_decoding32/N1916 ) );
  AND2_X4 U5711 ( .A1(n7325), .A2(n7659), .ZN(rs1_addr[4]) );
  INV_X1 U5712 ( .A(\Mcontrol/d_instr [26]), .ZN(net56678) );
  INV_X2 U5713 ( .A(\Mcontrol/d_instr [26]), .ZN(
        \Mcontrol/Operation_decoding32/N1922 ) );
  INV_X2 U5714 ( .A(\Mcontrol/d_instr [26]), .ZN(net56922) );
  INV_X2 U5715 ( .A(\Mcontrol/d_instr [26]), .ZN(net58533) );
  NAND2_X1 U5716 ( .A1(\Mpath/the_alu/N465 ), .A2(\Mpath/the_alu/N448 ), .ZN(
        n6497) );
  NAND2_X1 U5717 ( .A1(n7560), .A2(n7561), .ZN(n6957) );
  NAND2_X1 U5718 ( .A1(net56784), .A2(n6958), .ZN(n6988) );
  INV_X1 U5719 ( .A(n6957), .ZN(n6958) );
  NOR2_X2 U5720 ( .A1(n7032), .A2(n7149), .ZN(n7300) );
  NAND3_X4 U5721 ( .A1(n6018), .A2(rs2_addr[4]), .A3(n6030), .ZN(n5760) );
  AND2_X4 U5722 ( .A1(rs1_addr[1]), .A2(n7687), .ZN(n6414) );
  INV_X4 U5723 ( .A(rs1_addr[0]), .ZN(n7687) );
  INV_X1 U5724 ( .A(n1474), .ZN(n6959) );
  INV_X1 U5725 ( .A(n6959), .ZN(n6960) );
  OR2_X1 U5726 ( .A1(n2507), .A2(n2577), .ZN(n6961) );
  OR2_X1 U5727 ( .A1(n5515), .A2(n2509), .ZN(n6962) );
  NAND2_X1 U5728 ( .A1(n6961), .A2(n6962), .ZN(break_code[5]) );
  NAND2_X1 U5729 ( .A1(n6954), .A2(n7010), .ZN(net56216) );
  NAND3_X4 U5730 ( .A1(rs2_addr[1]), .A2(n6032), .A3(n6037), .ZN(n5777) );
  INV_X4 U5731 ( .A(net55921), .ZN(net57184) );
  NAND3_X4 U5732 ( .A1(n6030), .A2(rs2_addr[1]), .A3(n6037), .ZN(n5779) );
  NOR2_X2 U5733 ( .A1(n6034), .A2(rs2_addr[2]), .ZN(n6030) );
  NAND2_X1 U5734 ( .A1(n371), .A2(\Mcontrol/f_currpc[20] ), .ZN(n6963) );
  NAND2_X1 U5735 ( .A1(n7872), .A2(n372), .ZN(n6964) );
  INV_X1 U5736 ( .A(n373), .ZN(n6965) );
  AND3_X2 U5737 ( .A1(n6964), .A2(n6963), .A3(n6965), .ZN(n444) );
  INV_X1 U5738 ( .A(\regfile/N358 ), .ZN(n6966) );
  INV_X1 U5739 ( .A(n6966), .ZN(n6967) );
  INV_X1 U5740 ( .A(n1573), .ZN(n6968) );
  AND2_X2 U5741 ( .A1(\Mcontrol/m_sampled_xrd[4] ), .A2(n5503), .ZN(
        \regfile/N358 ) );
  OAI211_X1 U5742 ( .C1(\Mpath/the_alu/N81 ), .C2(n1695), .A(n2439), .B(n2440), 
        .ZN(daddr_out[1]) );
  INV_X1 U5743 ( .A(\regfile/N358 ), .ZN(n7195) );
  CLKBUF_X1 U5744 ( .A(\Mcontrol/Operation_decoding32/N1939 ), .Z(n6970) );
  NAND2_X1 U5745 ( .A1(n7009), .A2(n7010), .ZN(n7002) );
  NAND2_X1 U5746 ( .A1(\Mcontrol/Nextpc_decoding/Bta [23]), .A2(net58826), 
        .ZN(n7009) );
  INV_X2 U5747 ( .A(rs2_addr[0]), .ZN(n6019) );
  NOR2_X4 U5748 ( .A1(n6019), .A2(rs2_addr[4]), .ZN(n6037) );
  NOR2_X2 U5749 ( .A1(n6026), .A2(n6019), .ZN(n6029) );
  AND2_X2 U5750 ( .A1(n6025), .A2(n6019), .ZN(n6024) );
  AND3_X2 U5751 ( .A1(rs2_addr[4]), .A2(n6019), .A3(n6028), .ZN(n5763) );
  AND2_X4 U5752 ( .A1(n6028), .A2(n6029), .ZN(n5762) );
  CLKBUF_X1 U5753 ( .A(n7585), .Z(n6971) );
  OR2_X2 U5754 ( .A1(daddr_out[0]), .A2(daddr_out[1]), .ZN(\d_chk/N12 ) );
  INV_X8 U5755 ( .A(n7406), .ZN(n270) );
  INV_X8 U5756 ( .A(n7407), .ZN(n268) );
  NOR2_X1 U5757 ( .A1(n7200), .A2(n2451), .ZN(n2450) );
  OR2_X2 U5758 ( .A1(rd_addr[3]), .A2(\regfile/N358 ), .ZN(\regfile/N272 ) );
  AOI22_X1 U5759 ( .A1(n2441), .A2(\Mpath/the_alu/N82 ), .B1(n2442), .B2(n2443), .ZN(n2439) );
  INV_X1 U5760 ( .A(n7080), .ZN(n6972) );
  NAND2_X1 U5761 ( .A1(n7288), .A2(n7289), .ZN(n6973) );
  NAND2_X1 U5762 ( .A1(n7082), .A2(n6972), .ZN(n6974) );
  NAND2_X1 U5763 ( .A1(n1434), .A2(n7420), .ZN(n2792) );
  INV_X1 U5764 ( .A(n1673), .ZN(n6992) );
  INV_X1 U5765 ( .A(net58101), .ZN(n1500) );
  INV_X1 U5766 ( .A(net58101), .ZN(n6995) );
  INV_X1 U5767 ( .A(\Mcontrol/st_logic/branchlw_stall ), .ZN(
        \Mcontrol/st_logic/N13 ) );
  NAND2_X1 U5768 ( .A1(n7002), .A2(n372), .ZN(net56316) );
  NOR2_X4 U5769 ( .A1(n6034), .A2(n6022), .ZN(n6032) );
  NAND3_X4 U5770 ( .A1(n6018), .A2(rs2_addr[2]), .A3(n6021), .ZN(n5755) );
  OAI222_X2 U5771 ( .A1(n5564), .A2(n5523), .B1(n5565), .B2(n5525), .C1(n5566), 
        .C2(n5527), .ZN(branch_regb[26]) );
  INV_X4 U5772 ( .A(n5750), .ZN(n1936) );
  AOI21_X1 U5773 ( .B1(\Mcontrol/Nextpc_decoding/N36 ), .B2(
        \Mcontrol/Nextpc_decoding/N289 ), .A(\Mcontrol/Nextpc_decoding/N295 ), 
        .ZN(n6411) );
  INV_X2 U5774 ( .A(rs2_addr[2]), .ZN(n6022) );
  AND2_X2 U5775 ( .A1(n6976), .A2(n6975), .ZN(n5503) );
  INV_X32 U5776 ( .A(m_we), .ZN(n6975) );
  NAND2_X1 U5777 ( .A1(n7108), .A2(\Mcontrol/N17 ), .ZN(n6976) );
  INV_X1 U5778 ( .A(branch_rega[23]), .ZN(n7005) );
  OR2_X2 U5779 ( .A1(branch_rega[23]), .A2(branch_rega[24]), .ZN(n7635) );
  AND2_X2 U5780 ( .A1(n2447), .A2(\Mpath/the_alu/N473 ), .ZN(n7293) );
  NAND2_X1 U5781 ( .A1(\Mpath/the_alu/N474 ), .A2(n2447), .ZN(n1692) );
  NAND2_X1 U5782 ( .A1(n5503), .A2(\Mcontrol/m_sampled_xrd[0] ), .ZN(n1222) );
  NAND3_X4 U5783 ( .A1(n2311), .A2(n2312), .A3(n6028), .ZN(n1934) );
  CLKBUF_X1 U5784 ( .A(daddr_out[0]), .Z(n6977) );
  NAND2_X1 U5785 ( .A1(n6979), .A2(n7651), .ZN(n6978) );
  AND2_X1 U5786 ( .A1(n7624), .A2(n7136), .ZN(n6979) );
  INV_X1 U5787 ( .A(n6978), .ZN(n6980) );
  NAND2_X1 U5788 ( .A1(n7320), .A2(n6980), .ZN(n6981) );
  AND2_X1 U5789 ( .A1(\Mpath/the_alu/sum[31] ), .A2(n7634), .ZN(n7294) );
  NOR2_X1 U5790 ( .A1(n7281), .A2(n6982), .ZN(n7563) );
  NAND2_X1 U5791 ( .A1(n6983), .A2(n7046), .ZN(n6982) );
  NOR2_X1 U5792 ( .A1(n7282), .A2(n7472), .ZN(n6983) );
  NOR2_X2 U5793 ( .A1(n7468), .A2(n6984), .ZN(n7676) );
  NAND2_X2 U5794 ( .A1(n6985), .A2(n7644), .ZN(n6984) );
  NOR2_X1 U5795 ( .A1(n7265), .A2(n7153), .ZN(n6985) );
  AND2_X1 U5796 ( .A1(n6406), .A2(n6407), .ZN(n6986) );
  NOR2_X1 U5797 ( .A1(n6986), .A2(n6408), .ZN(n6405) );
  OAI222_X4 U5798 ( .A1(n5546), .A2(n5621), .B1(n5506), .B2(n7485), .C1(n5548), 
        .C2(n5623), .ZN(n7086) );
  AND4_X2 U5799 ( .A1(n2095), .A2(n2096), .A3(n2097), .A4(n2098), .ZN(n6987)
         );
  INV_X4 U5800 ( .A(n6987), .ZN(n93) );
  NOR2_X2 U5801 ( .A1(n7457), .A2(n7137), .ZN(n7696) );
  AND3_X4 U5802 ( .A1(n6029), .A2(rs2_addr[3]), .A3(n6025), .ZN(n5767) );
  AND2_X1 U5803 ( .A1(\Mpath/the_alu/diff[0] ), .A2(n1698), .ZN(n7200) );
  INV_X8 U5804 ( .A(n7362), .ZN(n255) );
  OR3_X4 U5805 ( .A1(\regfile/N367 ), .A2(net55892), .A3(n1108), .ZN(n7362) );
  AOI222_X1 U5806 ( .A1(n6102), .A2(n6538), .B1(
        \Mcontrol/Nextpc_decoding/Bta [8]), .B2(n1560), .C1(net57184), .C2(
        jar_in[8]), .ZN(n2525) );
  OAI222_X1 U5807 ( .A1(n5558), .A2(n5523), .B1(n5559), .B2(n5525), .C1(n5560), 
        .C2(n5527), .ZN(branch_regb[28]) );
  NOR2_X2 U5808 ( .A1(n6020), .A2(rs2_addr[0]), .ZN(n6018) );
  NAND2_X4 U5809 ( .A1(n6035), .A2(n6030), .ZN(n5778) );
  AND2_X4 U5810 ( .A1(n6018), .A2(n6026), .ZN(n6035) );
  INV_X2 U5811 ( .A(\Mcontrol/Operation_decoding32/N1898 ), .ZN(
        \Mcontrol/Operation_decoding32/N1899 ) );
  AND3_X4 U5812 ( .A1(n6024), .A2(n2312), .A3(rs2_addr[3]), .ZN(n1932) );
  NAND2_X1 U5813 ( .A1(\Mpath/the_alu/N1 ), .A2(n7171), .ZN(n6989) );
  OR2_X2 U5814 ( .A1(n7669), .A2(n7668), .ZN(n7672) );
  OR2_X1 U5815 ( .A1(\Mcontrol/Nextpc_decoding/N252 ), .A2(branch_rega[29]), 
        .ZN(\Mcontrol/Nextpc_decoding/N221 ) );
  INV_X8 U5816 ( .A(n5749), .ZN(n1938) );
  NAND3_X2 U5817 ( .A1(rs2_addr[0]), .A2(n6020), .A3(n6017), .ZN(n5749) );
  INV_X1 U5818 ( .A(n7690), .ZN(n7691) );
  AND2_X2 U5819 ( .A1(\Mcontrol/d_sampled_finstr [5]), .A2(n7278), .ZN(n7623)
         );
  AOI21_X2 U5820 ( .B1(\Scc_coproc/N580 ), .B2(\Scc_coproc/interrupt_active ), 
        .A(n5740), .ZN(\Scc_coproc/N553 ) );
  OR2_X2 U5821 ( .A1(rd_addr[2]), .A2(\regfile/N272 ), .ZN(\regfile/N273 ) );
  CLKBUF_X1 U5822 ( .A(net57942), .Z(net56319) );
  CLKBUF_X1 U5823 ( .A(net57184), .Z(net59543) );
  CLKBUF_X1 U5824 ( .A(n6951), .Z(net59767) );
  INV_X1 U5825 ( .A(n7041), .ZN(n7513) );
  BUF_X4 U5826 ( .A(n1935), .Z(n7017) );
  CLKBUF_X1 U5827 ( .A(n7878), .Z(I_ADDR_OUTBUS[13]) );
  CLKBUF_X1 U5828 ( .A(n7879), .Z(I_ADDR_OUTBUS[12]) );
  CLKBUF_X1 U5829 ( .A(n7877), .Z(I_ADDR_OUTBUS[14]) );
  CLKBUF_X1 U5830 ( .A(n7876), .Z(I_ADDR_OUTBUS[15]) );
  CLKBUF_X1 U5831 ( .A(n7885), .Z(I_ADDR_OUTBUS[3]) );
  INV_X1 U5832 ( .A(n5776), .ZN(n7023) );
  INV_X1 U5833 ( .A(n7023), .ZN(n7024) );
  INV_X4 U5834 ( .A(n7023), .ZN(n7025) );
  BUF_X4 U5835 ( .A(n5764), .Z(n7026) );
  AND3_X2 U5836 ( .A1(n7027), .A2(net55850), .A3(n7428), .ZN(n258) );
  NOR2_X1 U5837 ( .A1(rd_addr[2]), .A2(\regfile/N372 ), .ZN(n7027) );
  CLKBUF_X2 U5838 ( .A(n220), .Z(net55896) );
  INV_X2 U5839 ( .A(n1252), .ZN(n7428) );
  NOR2_X1 U5840 ( .A1(\Mcontrol/Operation_decoding32/N2087 ), .A2(n7028), .ZN(
        n7399) );
  OR2_X2 U5841 ( .A1(n7134), .A2(n7029), .ZN(n7028) );
  INV_X1 U5842 ( .A(n7072), .ZN(n7029) );
  OR2_X2 U5843 ( .A1(n7066), .A2(n7160), .ZN(
        \Mcontrol/Operation_decoding32/N1924 ) );
  NAND3_X4 U5844 ( .A1(n7190), .A2(n7191), .A3(\Mcontrol/N34 ), .ZN(n7030) );
  INV_X1 U5845 ( .A(n7215), .ZN(n7191) );
  AND3_X2 U5846 ( .A1(n7031), .A2(net58625), .A3(n7366), .ZN(n308) );
  INV_X32 U5847 ( .A(net55894), .ZN(net58625) );
  NOR2_X1 U5848 ( .A1(\regfile/N290 ), .A2(\regfile/N304 ), .ZN(n7031) );
  INV_X1 U5849 ( .A(n1107), .ZN(n7366) );
  OR2_X2 U5850 ( .A1(n7463), .A2(n7039), .ZN(n7032) );
  CLKBUF_X1 U5851 ( .A(n7535), .Z(n7033) );
  OR2_X1 U5852 ( .A1(n7652), .A2(n7065), .ZN(n7060) );
  AND2_X2 U5853 ( .A1(\Mcontrol/d_sampled_finstr [27]), .A2(n7278), .ZN(
        \Mcontrol/d_instr [27]) );
  CLKBUF_X1 U5854 ( .A(n7425), .Z(n7034) );
  NAND2_X1 U5855 ( .A1(n7099), .A2(n7307), .ZN(
        \Mcontrol/Operation_decoding32/N2070 ) );
  NOR2_X1 U5856 ( .A1(net58300), .A2(net57313), .ZN(n7035) );
  OR2_X1 U5857 ( .A1(n7124), .A2(n6956), .ZN(net58300) );
  OR2_X2 U5858 ( .A1(\Mcontrol/Operation_decoding32/N1990 ), .A2(
        \Mcontrol/d_instr [28]), .ZN(n7566) );
  CLKBUF_X1 U5859 ( .A(n7303), .Z(n7036) );
  INV_X1 U5860 ( .A(branch_rega[1]), .ZN(n7467) );
  NOR2_X2 U5861 ( .A1(\Mcontrol/Operation_decoding32/N2045 ), .A2(n7408), .ZN(
        n7087) );
  INV_X1 U5862 ( .A(n7175), .ZN(n7037) );
  BUF_X1 U5863 ( .A(n7673), .Z(n7055) );
  INV_X1 U5864 ( .A(n7034), .ZN(n7038) );
  INV_X1 U5865 ( .A(n7251), .ZN(n7039) );
  INV_X1 U5866 ( .A(n7251), .ZN(n7253) );
  NOR4_X1 U5867 ( .A1(n2671), .A2(n2672), .A3(n2673), .A4(n2674), .ZN(n2670)
         );
  AOI221_X1 U5868 ( .B1(n371), .B2(\Mcontrol/f_currpc[3] ), .C1(n372), .C2(
        n7885), .A(n373), .ZN(n848) );
  AND2_X1 U5869 ( .A1(\Mcontrol/Operation_decoding32/N2066 ), .A2(n7570), .ZN(
        n7040) );
  NAND2_X1 U5870 ( .A1(\Mcontrol/d_sampled_finstr [27]), .A2(n7278), .ZN(n7041) );
  NAND2_X2 U5871 ( .A1(\Mcontrol/Operation_decoding32/N2037 ), .A2(n7225), 
        .ZN(n6093) );
  CLKBUF_X1 U5872 ( .A(n6101), .Z(net58594) );
  NOR2_X2 U5873 ( .A1(n7253), .A2(n7599), .ZN(n7143) );
  CLKBUF_X1 U5874 ( .A(n7252), .Z(n7042) );
  OR2_X4 U5875 ( .A1(n3086), .A2(n7055), .ZN(n7043) );
  OAI221_X4 U5876 ( .B1(net55834), .B2(\Mcontrol/st_logic/N26 ), .C1(n5518), 
        .C2(net55918), .A(n1456), .ZN(n4368) );
  OAI221_X4 U5877 ( .B1(n2500), .B2(n2737), .C1(n5518), .C2(n2718), .A(n2719), 
        .ZN(break_code[18]) );
  INV_X1 U5878 ( .A(n7053), .ZN(n7522) );
  INV_X1 U5879 ( .A(n7053), .ZN(n7569) );
  OR2_X2 U5880 ( .A1(n7144), .A2(\Mcontrol/d_instr [26]), .ZN(n7225) );
  CLKBUF_X2 U5881 ( .A(\Mcontrol/Operation_decoding32/N2041 ), .Z(n7144) );
  AND2_X4 U5882 ( .A1(n7167), .A2(n7168), .ZN(
        \Mcontrol/Operation_decoding32/N89 ) );
  INV_X2 U5883 ( .A(n7055), .ZN(n7207) );
  OR2_X2 U5884 ( .A1(\Mcontrol/Operation_decoding32/N1996 ), .A2(n7536), .ZN(
        n7044) );
  NOR2_X2 U5885 ( .A1(n7060), .A2(n7045), .ZN(n7390) );
  OR2_X1 U5886 ( .A1(n7536), .A2(n7099), .ZN(n7045) );
  NOR2_X1 U5887 ( .A1(net57843), .A2(branch_rega[23]), .ZN(n7046) );
  CLKBUF_X1 U5888 ( .A(n7504), .Z(n7047) );
  NOR2_X1 U5889 ( .A1(n7032), .A2(n7048), .ZN(n7419) );
  NAND2_X1 U5890 ( .A1(n7050), .A2(n7099), .ZN(n7048) );
  AND2_X1 U5891 ( .A1(\Mcontrol/Operation_decoding32/N1963 ), .A2(
        \Mcontrol/Operation_decoding32/N1969 ), .ZN(n7049) );
  BUF_X2 U5892 ( .A(n7065), .Z(n7098) );
  NAND3_X4 U5893 ( .A1(rs2_addr[1]), .A2(n6029), .A3(n6030), .ZN(n5759) );
  INV_X1 U5894 ( .A(n7222), .ZN(n7050) );
  OR2_X1 U5895 ( .A1(n7252), .A2(n7462), .ZN(n7051) );
  INV_X2 U5896 ( .A(n7513), .ZN(n7052) );
  NAND2_X1 U5897 ( .A1(\Mcontrol/d_sampled_finstr [26]), .A2(n7278), .ZN(n7053) );
  AND2_X2 U5898 ( .A1(n7143), .A2(n7455), .ZN(n7307) );
  NAND2_X1 U5899 ( .A1(n7152), .A2(n7252), .ZN(n7054) );
  AOI221_X1 U5900 ( .B1(n1417), .B2(n2497), .C1(n6970), .C2(n2501), .A(n7441), 
        .ZN(n2499) );
  NAND2_X2 U5901 ( .A1(n7546), .A2(n7522), .ZN(n7568) );
  NAND2_X1 U5902 ( .A1(n1846), .A2(n7585), .ZN(n2494) );
  NAND2_X1 U5903 ( .A1(net56765), .A2(n7056), .ZN(n7524) );
  NOR2_X1 U5904 ( .A1(\Mcontrol/Operation_decoding32/N2021 ), .A2(n7299), .ZN(
        n7056) );
  NOR2_X1 U5905 ( .A1(n7057), .A2(net57236), .ZN(net57253) );
  NAND2_X1 U5906 ( .A1(\Mcontrol/Operation_decoding32/N2084 ), .A2(net58547), 
        .ZN(n7057) );
  INV_X2 U5907 ( .A(net57388), .ZN(net57236) );
  INV_X1 U5908 ( .A(\Mcontrol/Operation_decoding32/N2017 ), .ZN(net58542) );
  INV_X1 U5909 ( .A(net58542), .ZN(net58543) );
  OR2_X1 U5910 ( .A1(net56678), .A2(n7125), .ZN(n7058) );
  NOR2_X1 U5911 ( .A1(n7088), .A2(n7125), .ZN(n7059) );
  OR2_X1 U5912 ( .A1(n7053), .A2(n7299), .ZN(n7126) );
  AND2_X1 U5913 ( .A1(n6066), .A2(n7438), .ZN(n7061) );
  INV_X1 U5914 ( .A(n7647), .ZN(n7062) );
  OR2_X2 U5915 ( .A1(n7673), .A2(n7653), .ZN(n7647) );
  INV_X1 U5916 ( .A(n1509), .ZN(n7063) );
  INV_X2 U5917 ( .A(n7254), .ZN(n7536) );
  OR2_X2 U5918 ( .A1(\Mcontrol/Operation_decoding32/N2056 ), .A2(n7536), .ZN(
        \Mcontrol/Operation_decoding32/N2045 ) );
  CLKBUF_X1 U5919 ( .A(\Mcontrol/Operation_decoding32/N1951 ), .Z(n7064) );
  INV_X1 U5920 ( .A(n7246), .ZN(n7065) );
  INV_X1 U5921 ( .A(n7246), .ZN(n7251) );
  NAND2_X1 U5922 ( .A1(\Mcontrol/Operation_decoding32/N1921 ), .A2(net56922), 
        .ZN(n7515) );
  NOR2_X2 U5923 ( .A1(\Mcontrol/Operation_decoding32/N1917 ), .A2(n6907), .ZN(
        n7167) );
  OR2_X2 U5924 ( .A1(n7146), .A2(\Mcontrol/Operation_decoding32/N1916 ), .ZN(
        \Mcontrol/Operation_decoding32/N1917 ) );
  OR2_X2 U5925 ( .A1(n7463), .A2(n7039), .ZN(n7066) );
  AND2_X1 U5926 ( .A1(n7536), .A2(n7062), .ZN(n7067) );
  NAND2_X1 U5927 ( .A1(n7067), .A2(n7068), .ZN(
        \Mcontrol/Operation_decoding32/N1955 ) );
  AND2_X1 U5928 ( .A1(n7069), .A2(n7098), .ZN(n7068) );
  INV_X1 U5929 ( .A(\Mcontrol/d_instr [28]), .ZN(n7069) );
  NAND2_X1 U5930 ( .A1(n7152), .A2(n7039), .ZN(
        \Mcontrol/Operation_decoding32/N1990 ) );
  NOR2_X1 U5931 ( .A1(\Mcontrol/Operation_decoding32/N2087 ), .A2(n7070), .ZN(
        n7400) );
  NAND2_X1 U5932 ( .A1(n7221), .A2(n7041), .ZN(n7070) );
  OR2_X2 U5933 ( .A1(n7536), .A2(n7051), .ZN(
        \Mcontrol/Operation_decoding32/N2087 ) );
  CLKBUF_X2 U5934 ( .A(net57253), .Z(net56996) );
  INV_X2 U5935 ( .A(n7415), .ZN(\Mcontrol/Operation_decoding32/N2037 ) );
  OR2_X2 U5936 ( .A1(n7569), .A2(\Mcontrol/Operation_decoding32/N2035 ), .ZN(
        n7415) );
  CLKBUF_X1 U5937 ( .A(n7049), .Z(n7071) );
  INV_X4 U5938 ( .A(n1107), .ZN(n7291) );
  INV_X4 U5939 ( .A(n1107), .ZN(n7316) );
  INV_X2 U5940 ( .A(n1107), .ZN(n7417) );
  INV_X2 U5941 ( .A(n1107), .ZN(n7364) );
  OR3_X1 U5942 ( .A1(\regfile/N427 ), .A2(net55888), .A3(n1107), .ZN(n7120) );
  INV_X1 U5943 ( .A(n7041), .ZN(n7072) );
  INV_X1 U5944 ( .A(n311), .ZN(n7073) );
  INV_X8 U5945 ( .A(n7073), .ZN(n7074) );
  NOR3_X1 U5946 ( .A1(\regfile/N311 ), .A2(net55896), .A3(n1251), .ZN(n311) );
  INV_X2 U5947 ( .A(n303), .ZN(n7075) );
  INV_X4 U5948 ( .A(n7075), .ZN(n7076) );
  OR2_X2 U5949 ( .A1(n7060), .A2(n7222), .ZN(n7088) );
  NOR2_X1 U5950 ( .A1(n7077), .A2(\Mcontrol/Operation_decoding32/N2056 ), .ZN(
        n7435) );
  NAND2_X1 U5951 ( .A1(\Mcontrol/d_instr [28]), .A2(n7455), .ZN(n7077) );
  CLKBUF_X1 U5952 ( .A(n7043), .Z(n7078) );
  AND2_X2 U5953 ( .A1(n6066), .A2(n7438), .ZN(n6103) );
  AND2_X1 U5954 ( .A1(n7528), .A2(n7043), .ZN(n7079) );
  NAND2_X1 U5955 ( .A1(n7649), .A2(n7674), .ZN(n7080) );
  INV_X1 U5956 ( .A(n7597), .ZN(n7081) );
  NOR2_X1 U5957 ( .A1(n7257), .A2(n7081), .ZN(n7082) );
  OAI211_X1 U5958 ( .C1(n1556), .C2(n1557), .A(n1558), .B(n1559), .ZN(n7083)
         );
  NOR2_X1 U5959 ( .A1(n7478), .A2(n7477), .ZN(n7084) );
  NOR2_X1 U5960 ( .A1(n7479), .A2(n7085), .ZN(n1559) );
  INV_X1 U5961 ( .A(n7084), .ZN(n7085) );
  OAI211_X1 U5962 ( .C1(n1556), .C2(n1557), .A(n1558), .B(n1559), .ZN(n871) );
  AND2_X1 U5963 ( .A1(n6102), .A2(n6542), .ZN(n7477) );
  AND2_X1 U5964 ( .A1(jar_in[1]), .A2(n1561), .ZN(n7479) );
  INV_X2 U5965 ( .A(n6435), .ZN(n5546) );
  OR2_X2 U5966 ( .A1(n7256), .A2(n7043), .ZN(n7408) );
  NOR2_X1 U5967 ( .A1(n7408), .A2(\Mcontrol/Operation_decoding32/N2045 ), .ZN(
        n7546) );
  AND2_X1 U5968 ( .A1(n7351), .A2(n7623), .ZN(
        \Mcontrol/Operation_decoding32/N1883 ) );
  OR2_X2 U5969 ( .A1(n7351), .A2(n7623), .ZN(
        \Mcontrol/Operation_decoding32/N1908 ) );
  INV_X1 U5970 ( .A(n7246), .ZN(n7263) );
  OR2_X4 U5971 ( .A1(n7100), .A2(n3087), .ZN(n7256) );
  INV_X1 U5972 ( .A(\Mcontrol/d_instr [28]), .ZN(n7221) );
  OR2_X1 U5973 ( .A1(n7398), .A2(\Mcontrol/Operation_decoding32/N2070 ), .ZN(
        n7570) );
  OR2_X2 U5974 ( .A1(n7584), .A2(n7235), .ZN(n7397) );
  NAND2_X2 U5975 ( .A1(n7090), .A2(n7091), .ZN(n7089) );
  NOR2_X1 U5976 ( .A1(branch_rega[13]), .A2(n7495), .ZN(n7090) );
  NOR2_X1 U5977 ( .A1(branch_rega[15]), .A2(branch_rega[14]), .ZN(n7091) );
  NAND2_X2 U5978 ( .A1(n7448), .A2(net58533), .ZN(n7535) );
  NAND2_X2 U5979 ( .A1(\Mcontrol/Operation_decoding32/N1951 ), .A2(
        \Mcontrol/Operation_decoding32/N1957 ), .ZN(n6068) );
  NAND2_X1 U5980 ( .A1(n7087), .A2(n7522), .ZN(n7092) );
  OR2_X1 U5981 ( .A1(rd_addr[2]), .A2(\regfile/N420 ), .ZN(\regfile/N421 ) );
  OR2_X1 U5982 ( .A1(rd_addr[2]), .A2(\regfile/N323 ), .ZN(\regfile/N324 ) );
  OR2_X1 U5983 ( .A1(rd_addr[2]), .A2(\regfile/N317 ), .ZN(\regfile/N318 ) );
  OR2_X1 U5984 ( .A1(rd_addr[2]), .A2(\regfile/N414 ), .ZN(\regfile/N415 ) );
  OR2_X1 U5985 ( .A1(rd_addr[2]), .A2(\regfile/N432 ), .ZN(\regfile/N433 ) );
  OR2_X1 U5986 ( .A1(rd_addr[2]), .A2(\regfile/N378 ), .ZN(\regfile/N379 ) );
  OR2_X1 U5987 ( .A1(rd_addr[2]), .A2(\regfile/N335 ), .ZN(\regfile/N336 ) );
  OR2_X1 U5988 ( .A1(rd_addr[2]), .A2(\regfile/N384 ), .ZN(\regfile/N385 ) );
  OR2_X1 U5989 ( .A1(rd_addr[2]), .A2(\regfile/N426 ), .ZN(\regfile/N427 ) );
  OR2_X1 U5990 ( .A1(rd_addr[2]), .A2(\regfile/N366 ), .ZN(\regfile/N367 ) );
  OR2_X1 U5991 ( .A1(rd_addr[2]), .A2(\regfile/N285 ), .ZN(\regfile/N286 ) );
  INV_X2 U5992 ( .A(rd_addr[2]), .ZN(\regfile/N290 ) );
  AND2_X2 U5993 ( .A1(n6413), .A2(n6414), .ZN(n5628) );
  NOR4_X1 U5994 ( .A1(n2654), .A2(n2655), .A3(n2656), .A4(n2657), .ZN(n2653)
         );
  INV_X1 U5995 ( .A(branch_rega[21]), .ZN(n7443) );
  OR2_X1 U5996 ( .A1(branch_rega[21]), .A2(branch_rega[20]), .ZN(n7588) );
  INV_X1 U5997 ( .A(n7623), .ZN(n5515) );
  NAND2_X1 U5998 ( .A1(n7568), .A2(\Mcontrol/Operation_decoding32/N2054 ), 
        .ZN(n7093) );
  OR2_X2 U5999 ( .A1(n7520), .A2(n7521), .ZN(
        \Mcontrol/Operation_decoding32/N2054 ) );
  INV_X1 U6000 ( .A(n7632), .ZN(n7633) );
  INV_X2 U6001 ( .A(n7110), .ZN(serve_exception) );
  INV_X4 U6002 ( .A(n7107), .ZN(n7110) );
  NOR2_X4 U6003 ( .A1(n1049), .A2(n1050), .ZN(n362) );
  AND2_X4 U6004 ( .A1(rs1_addr[4]), .A2(n7686), .ZN(n6417) );
  OAI211_X2 U6005 ( .C1(n2523), .C2(n1557), .A(n2524), .B(n2525), .ZN(
        I_ADDR_OUTBUS[8]) );
  AND2_X1 U6006 ( .A1(\Mcontrol/d_sampled_finstr [27]), .A2(n7278), .ZN(n7526)
         );
  INV_X1 U6007 ( .A(n7697), .ZN(n7698) );
  OR2_X2 U6008 ( .A1(n7204), .A2(n7205), .ZN(n7357) );
  AND3_X2 U6009 ( .A1(n6025), .A2(rs2_addr[0]), .A3(n6021), .ZN(n5757) );
  NAND3_X2 U6010 ( .A1(rs2_addr[2]), .A2(n6034), .A3(n6035), .ZN(n5772) );
  OR2_X2 U6011 ( .A1(\Mcontrol/Operation_decoding32/N2070 ), .A2(n7398), .ZN(
        n7379) );
  OR2_X2 U6012 ( .A1(net57366), .A2(\Mcontrol/Operation_decoding32/N1944 ), 
        .ZN(n7585) );
  NAND2_X1 U6013 ( .A1(n5637), .A2(\regfile/reg_out[25][12] ), .ZN(n7094) );
  NAND2_X1 U6014 ( .A1(n5638), .A2(\regfile/reg_out[24][12] ), .ZN(n7095) );
  AND2_X2 U6015 ( .A1(n7094), .A2(n7095), .ZN(n6361) );
  CLKBUF_X1 U6016 ( .A(n5638), .Z(n7096) );
  NAND2_X1 U6017 ( .A1(n7508), .A2(n7097), .ZN(n7301) );
  NOR2_X1 U6018 ( .A1(n7401), .A2(\Mcontrol/d_instr [26]), .ZN(n7097) );
  OR2_X2 U6019 ( .A1(n7599), .A2(n7065), .ZN(
        \Mcontrol/Operation_decoding32/N1996 ) );
  CLKBUF_X1 U6020 ( .A(n7256), .Z(n7099) );
  AND2_X2 U6021 ( .A1(n6417), .A2(n7173), .ZN(n6413) );
  OAI22_X2 U6022 ( .A1(n5656), .A2(n5657), .B1(n5658), .B2(n5659), .ZN(n5655)
         );
  OAI211_X2 U6023 ( .C1(n2574), .C2(n1557), .A(n2575), .B(n2576), .ZN(
        I_ADDR_OUTBUS[5]) );
  AOI221_X1 U6024 ( .B1(n1561), .B2(jar_in[0]), .C1(n1564), .C2(n6102), .A(
        n1565), .ZN(n1043) );
  INV_X1 U6025 ( .A(n6073), .ZN(n7100) );
  INV_X1 U6026 ( .A(n6073), .ZN(n7277) );
  OAI222_X4 U6027 ( .A1(n7454), .A2(n6051), .B1(n7279), .B2(n5517), .C1(n5515), 
        .C2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n6156) );
  AND2_X2 U6028 ( .A1(n6021), .A2(n6022), .ZN(n6017) );
  AND3_X2 U6029 ( .A1(n6020), .A2(n6022), .A3(n6033), .ZN(n1931) );
  AND2_X1 U6030 ( .A1(n7573), .A2(n7572), .ZN(n7203) );
  NAND2_X1 U6031 ( .A1(n371), .A2(\Mcontrol/f_currpc[21] ), .ZN(n7101) );
  NAND2_X1 U6032 ( .A1(n7871), .A2(n372), .ZN(n7102) );
  INV_X1 U6033 ( .A(n373), .ZN(n7103) );
  INV_X1 U6034 ( .A(n7392), .ZN(n7394) );
  INV_X1 U6035 ( .A(n1905), .ZN(n5658) );
  AOI22_X2 U6036 ( .A1(n7503), .A2(\regfile/reg_out[21][12] ), .B1(n7611), 
        .B2(\regfile/reg_out[20][12] ), .ZN(n6360) );
  INV_X2 U6037 ( .A(n5651), .ZN(n7516) );
  NOR4_X2 U6038 ( .A1(n2343), .A2(n2344), .A3(n2345), .A4(n2346), .ZN(n2342)
         );
  NOR4_X2 U6039 ( .A1(n2866), .A2(n2867), .A3(n2868), .A4(n2869), .ZN(n2865)
         );
  INV_X2 U6040 ( .A(branch_rega[12]), .ZN(n7644) );
  INV_X2 U6041 ( .A(\Mpath/out_regB[13] ), .ZN(n7104) );
  INV_X1 U6042 ( .A(n7104), .ZN(n7105) );
  INV_X2 U6043 ( .A(n7104), .ZN(n7106) );
  INV_X2 U6044 ( .A(\Scc_coproc/N553 ), .ZN(n7107) );
  INV_X1 U6045 ( .A(n7107), .ZN(n7108) );
  INV_X1 U6046 ( .A(n7107), .ZN(n7109) );
  INV_X1 U6047 ( .A(n306), .ZN(n7111) );
  INV_X8 U6048 ( .A(n7111), .ZN(n7112) );
  NOR3_X2 U6049 ( .A1(\regfile/N299 ), .A2(net55894), .A3(n1252), .ZN(n306) );
  OR3_X4 U6050 ( .A1(\regfile/N293 ), .A2(net55892), .A3(n1108), .ZN(n7113) );
  INV_X4 U6051 ( .A(n7113), .ZN(n304) );
  OAI21_X2 U6052 ( .B1(\Mpath/the_alu/N465 ), .B2(n6496), .A(n6497), .ZN(
        \exc[ALU_OFLOW1] ) );
  INV_X1 U6053 ( .A(branch_rega[6]), .ZN(n7444) );
  INV_X1 U6054 ( .A(branch_rega[6]), .ZN(n7597) );
  INV_X1 U6055 ( .A(n261), .ZN(n7114) );
  INV_X4 U6056 ( .A(n7114), .ZN(n7115) );
  NOR3_X1 U6057 ( .A1(\regfile/N379 ), .A2(net55892), .A3(n1107), .ZN(n261) );
  INV_X2 U6058 ( .A(n260), .ZN(n7116) );
  INV_X4 U6059 ( .A(n7116), .ZN(n7117) );
  INV_X2 U6060 ( .A(n258), .ZN(n260) );
  INV_X2 U6061 ( .A(n285), .ZN(n7118) );
  INV_X8 U6062 ( .A(n7118), .ZN(n7119) );
  NOR3_X1 U6063 ( .A1(\regfile/N433 ), .A2(net55894), .A3(n1251), .ZN(n285) );
  INV_X1 U6064 ( .A(n280), .ZN(n7121) );
  INV_X8 U6065 ( .A(n7121), .ZN(n7122) );
  NOR3_X2 U6066 ( .A1(\regfile/N421 ), .A2(net55888), .A3(n1252), .ZN(n280) );
  INV_X1 U6067 ( .A(branch_rega[5]), .ZN(n7649) );
  AND2_X2 U6068 ( .A1(\Scc_coproc/x_exc_word[4] ), .A2(
        \Scc_coproc/x_exc_word[5] ), .ZN(\Scc_coproc/N576 ) );
  BUF_X4 U6069 ( .A(\Mpath/out_regB[2] ), .Z(n7711) );
  INV_X4 U6070 ( .A(branch_rega[14]), .ZN(n7704) );
  OR2_X1 U6071 ( .A1(branch_rega[14]), .A2(branch_rega[13]), .ZN(n7697) );
  OAI222_X1 U6072 ( .A1(n5534), .A2(n5523), .B1(n5535), .B2(n5525), .C1(n5536), 
        .C2(n5527), .ZN(branch_regb[6]) );
  NAND2_X4 U6073 ( .A1(\BYP_BRANCH_MUXB/N4 ), .A2(\Mcontrol/st_logic/N42 ), 
        .ZN(n5523) );
  INV_X4 U6074 ( .A(\BYP_BRANCH_MUXB/N39 ), .ZN(\BYP_BRANCH_MUXB/N4 ) );
  NAND2_X1 U6075 ( .A1(n7132), .A2(n7133), .ZN(n7123) );
  AND2_X2 U6076 ( .A1(\Mcontrol/d_instr [28]), .A2(n7098), .ZN(n7133) );
  OR2_X2 U6077 ( .A1(\Mcontrol/Operation_decoding32/N2062 ), .A2(n7536), .ZN(
        n7124) );
  AND2_X2 U6078 ( .A1(n7535), .A2(n7379), .ZN(n7543) );
  NAND2_X2 U6079 ( .A1(n1817), .A2(n1818), .ZN(n6155) );
  BUF_X8 U6080 ( .A(\Mpath/out_regB[2] ), .Z(n7709) );
  NAND2_X1 U6081 ( .A1(\Mcontrol/d_instr [27]), .A2(n7256), .ZN(n7125) );
  AND2_X1 U6082 ( .A1(n7203), .A2(n7127), .ZN(n7288) );
  NOR2_X1 U6083 ( .A1(n7496), .A2(branch_rega[19]), .ZN(n7127) );
  OR2_X2 U6084 ( .A1(n7044), .A2(n7523), .ZN(
        \Mcontrol/Operation_decoding32/N2005 ) );
  OR2_X2 U6085 ( .A1(\Mcontrol/Operation_decoding32/N2064 ), .A2(n7515), .ZN(
        \Mcontrol/Operation_decoding32/N2066 ) );
  INV_X1 U6086 ( .A(n7538), .ZN(n7128) );
  NAND2_X1 U6087 ( .A1(n7537), .A2(n7129), .ZN(
        \Mcontrol/Operation_decoding32/N2030 ) );
  NOR2_X1 U6088 ( .A1(net58533), .A2(n7128), .ZN(n7129) );
  NOR2_X1 U6089 ( .A1(n7160), .A2(n7054), .ZN(n7537) );
  OAI222_X1 U6090 ( .A1(n5623), .A2(n5608), .B1(n7487), .B2(n2827), .C1(n5621), 
        .C2(n5606), .ZN(branch_rega[13]) );
  INV_X1 U6091 ( .A(branch_rega[13]), .ZN(n7646) );
  OR2_X1 U6092 ( .A1(n7566), .A2(n7233), .ZN(
        \Mcontrol/Operation_decoding32/N2035 ) );
  AND2_X1 U6093 ( .A1(n6073), .A2(n7151), .ZN(n7246) );
  AND3_X1 U6094 ( .A1(n1849), .A2(n7524), .A3(n7164), .ZN(n6066) );
  AND2_X2 U6095 ( .A1(n7660), .A2(n7661), .ZN(n7626) );
  INV_X2 U6096 ( .A(n7481), .ZN(n7482) );
  CLKBUF_X1 U6097 ( .A(\Scc_coproc/x_exc_word[5] ), .Z(n7130) );
  AND2_X1 U6098 ( .A1(n2450), .A2(n2449), .ZN(n7131) );
  NOR2_X1 U6099 ( .A1(n1509), .A2(n7545), .ZN(n7132) );
  NAND2_X1 U6100 ( .A1(n7132), .A2(n7133), .ZN(n7520) );
  INV_X1 U6101 ( .A(\Mcontrol/Operation_decoding32/N1989 ), .ZN(n7134) );
  AND3_X2 U6102 ( .A1(n7524), .A2(n1849), .A3(n7164), .ZN(n7135) );
  NOR2_X2 U6103 ( .A1(n7423), .A2(n7539), .ZN(n7577) );
  INV_X1 U6104 ( .A(n7240), .ZN(n7136) );
  NAND2_X1 U6105 ( .A1(n7138), .A2(n7443), .ZN(n7137) );
  NOR2_X1 U6106 ( .A1(n7458), .A2(branch_rega[24]), .ZN(n7138) );
  CLKBUF_X1 U6107 ( .A(n7874), .Z(I_ADDR_OUTBUS[17]) );
  AND2_X1 U6108 ( .A1(n6102), .A2(n6532), .ZN(n7140) );
  AND2_X1 U6109 ( .A1(\Mcontrol/Nextpc_decoding/Bta [17]), .A2(n7356), .ZN(
        n7141) );
  AND2_X1 U6110 ( .A1(jar_in[17]), .A2(net59543), .ZN(n7142) );
  NOR3_X1 U6111 ( .A1(n7140), .A2(n7141), .A3(n7142), .ZN(n2753) );
  AND2_X1 U6112 ( .A1(n7349), .A2(n7350), .ZN(n7511) );
  NOR2_X1 U6113 ( .A1(branch_rega[28]), .A2(\Mcontrol/Nextpc_decoding/N188 ), 
        .ZN(n7350) );
  OR2_X2 U6114 ( .A1(\Mcontrol/Operation_decoding32/N1968 ), .A2(n7522), .ZN(
        \Mcontrol/Operation_decoding32/N1969 ) );
  INV_X1 U6115 ( .A(n7455), .ZN(n7145) );
  INV_X2 U6116 ( .A(n7145), .ZN(n7146) );
  NOR2_X2 U6117 ( .A1(n7357), .A2(n7147), .ZN(n1560) );
  AND2_X2 U6118 ( .A1(n6097), .A2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(
        net57810) );
  INV_X1 U6119 ( .A(n7455), .ZN(n7148) );
  NAND2_X1 U6120 ( .A1(n7256), .A2(n7148), .ZN(n7149) );
  INV_X1 U6121 ( .A(n7150), .ZN(n7151) );
  INV_X1 U6122 ( .A(n7545), .ZN(n7152) );
  OAI22_X1 U6123 ( .A1(n6404), .A2(\Mcontrol/Nextpc_decoding/N31 ), .B1(n6405), 
        .B2(\Mcontrol/Nextpc_decoding/N313 ), .ZN(n7154) );
  OAI22_X2 U6124 ( .A1(n5517), .A2(n2594), .B1(n2595), .B2(n2613), .ZN(
        break_code[3]) );
  OAI221_X4 U6125 ( .B1(n5516), .B2(n1443), .C1(\Mpath/the_alu/N453 ), .C2(
        net55850), .A(n1476), .ZN(n4373) );
  OR2_X1 U6126 ( .A1(\Mpath/the_alu/N453 ), .A2(\Alu_command[OP][5] ), .ZN(
        \Mpath/the_alu/N454 ) );
  OR2_X1 U6127 ( .A1(\Mpath/the_alu/N453 ), .A2(\Mpath/the_alu/N466 ), .ZN(
        \Mpath/the_alu/N469 ) );
  OAI22_X2 U6128 ( .A1(n2507), .A2(n2526), .B1(n5914), .B2(n2509), .ZN(
        break_code[8]) );
  INV_X2 U6129 ( .A(n7646), .ZN(n7153) );
  NAND2_X1 U6130 ( .A1(n371), .A2(\Mcontrol/f_currpc[2] ), .ZN(n7155) );
  NAND2_X1 U6131 ( .A1(n372), .A2(n7886), .ZN(n7156) );
  INV_X1 U6132 ( .A(n373), .ZN(n7157) );
  AND3_X2 U6133 ( .A1(n7155), .A2(n7156), .A3(n7157), .ZN(n859) );
  OAI22_X2 U6134 ( .A1(\Mpath/the_alu/N520 ), .A2(n2457), .B1(
        \Mpath/the_alu/N526 ), .B2(\Mpath/the_alu/N468 ), .ZN(n1696) );
  OR2_X2 U6135 ( .A1(\Mpath/the_alu/N485 ), .A2(n6500), .ZN(n1694) );
  INV_X1 U6136 ( .A(n6500), .ZN(n2446) );
  OAI221_X1 U6137 ( .B1(\Mpath/the_alu/N29 ), .B2(n1693), .C1(n1841), .C2(
        n1884), .A(n1694), .ZN(n1882) );
  OAI221_X1 U6138 ( .B1(\Mpath/the_alu/N35 ), .B2(n1693), .C1(n1841), .C2(
        n1859), .A(n1694), .ZN(n1858) );
  OAI221_X1 U6139 ( .B1(\Mpath/the_alu/N31 ), .B2(n1693), .C1(n1841), .C2(
        n1875), .A(n1694), .ZN(n1874) );
  OAI221_X1 U6140 ( .B1(\Mpath/the_alu/N25 ), .B2(n1693), .C1(n1841), .C2(
        n1902), .A(n1694), .ZN(n1900) );
  OAI221_X1 U6141 ( .B1(\Mpath/the_alu/N33 ), .B2(n1693), .C1(n1841), .C2(
        n1867), .A(n1694), .ZN(n1866) );
  OAI221_X1 U6142 ( .B1(\Mpath/the_alu/N23 ), .B2(n1693), .C1(n1841), .C2(
        n1911), .A(n1694), .ZN(n1909) );
  OAI221_X1 U6143 ( .B1(\Mpath/the_alu/N27 ), .B2(n1693), .C1(n1841), .C2(
        n1893), .A(n1694), .ZN(n1891) );
  OR3_X2 U6144 ( .A1(\regfile/N385 ), .A2(net55896), .A3(n1251), .ZN(n7158) );
  INV_X4 U6145 ( .A(n7158), .ZN(n263) );
  INV_X1 U6146 ( .A(n7351), .ZN(n5516) );
  OR2_X2 U6147 ( .A1(n7253), .A2(n7545), .ZN(
        \Mcontrol/Operation_decoding32/N2056 ) );
  AND2_X1 U6148 ( .A1(n7036), .A2(n7304), .ZN(n7159) );
  NOR2_X2 U6149 ( .A1(n7044), .A2(n6956), .ZN(n7303) );
  INV_X1 U6150 ( .A(n7254), .ZN(n7160) );
  NOR2_X1 U6151 ( .A1(n7357), .A2(n7161), .ZN(n7356) );
  INV_X1 U6152 ( .A(n7071), .ZN(n7162) );
  NAND2_X1 U6153 ( .A1(\Mcontrol/Operation_decoding32/N1963 ), .A2(
        \Mcontrol/Operation_decoding32/N1969 ), .ZN(n7544) );
  AND2_X1 U6154 ( .A1(\Scc_coproc/x_exc_word[0] ), .A2(\Scc_coproc/N579 ), 
        .ZN(n7163) );
  CLKBUF_X1 U6155 ( .A(n7272), .Z(n7164) );
  NOR2_X1 U6156 ( .A1(\Mcontrol/Operation_decoding32/N1922 ), .A2(n7247), .ZN(
        n7166) );
  NOR2_X1 U6157 ( .A1(net56922), .A2(n7247), .ZN(n7165) );
  NOR2_X1 U6158 ( .A1(\Mcontrol/Operation_decoding32/N1922 ), .A2(n7247), .ZN(
        n7539) );
  NOR2_X1 U6159 ( .A1(n7522), .A2(n7513), .ZN(n7168) );
  INV_X2 U6160 ( .A(n1222), .ZN(n1379) );
  NAND2_X1 U6161 ( .A1(\Mcontrol/Operation_decoding32/N89 ), .A2(
        \Mcontrol/Operation_decoding32/N1975 ), .ZN(n7169) );
  NAND3_X1 U6162 ( .A1(n1844), .A2(n6059), .A3(n7170), .ZN(n6094) );
  INV_X1 U6163 ( .A(n7169), .ZN(n7170) );
  OR2_X1 U6164 ( .A1(\Mcontrol/Operation_decoding32/N2087 ), .A2(
        \Mcontrol/Operation_decoding32/N1989 ), .ZN(
        \Mcontrol/Operation_decoding32/N2046 ) );
  AND2_X2 U6165 ( .A1(\Scc_coproc/x_exc_word[0] ), .A2(\Scc_coproc/N579 ), 
        .ZN(\Scc_coproc/N580 ) );
  NAND2_X1 U6166 ( .A1(n1733), .A2(n1734), .ZN(n6345) );
  NAND3_X1 U6167 ( .A1(n6428), .A2(rs1_addr[4]), .A3(n6414), .ZN(n5640) );
  INV_X2 U6168 ( .A(n1841), .ZN(n1697) );
  NOR2_X1 U6169 ( .A1(\Alu_command[OP][0] ), .A2(\Mpath/the_alu/N457 ), .ZN(
        n7171) );
  NOR2_X1 U6170 ( .A1(n7172), .A2(\Mcontrol/Operation_decoding32/N2003 ), .ZN(
        \Mcontrol/Operation_decoding32/N2007 ) );
  OR2_X1 U6171 ( .A1(\Mcontrol/d_instr [26]), .A2(n7523), .ZN(n7172) );
  NAND3_X1 U6172 ( .A1(n7687), .A2(n6416), .A3(n6413), .ZN(n5625) );
  INV_X1 U6173 ( .A(n7481), .ZN(n7483) );
  AND2_X4 U6174 ( .A1(n7326), .A2(n5903), .ZN(n7173) );
  INV_X4 U6175 ( .A(n7173), .ZN(rs1_addr[2]) );
  CLKBUF_X1 U6176 ( .A(n7135), .Z(n7174) );
  NAND2_X1 U6177 ( .A1(n7303), .A2(n7304), .ZN(n7175) );
  AND3_X4 U6178 ( .A1(n7382), .A2(rs1_addr[3]), .A3(n6433), .ZN(n2332) );
  INV_X1 U6179 ( .A(n7254), .ZN(n1509) );
  CLKBUF_X1 U6180 ( .A(n7279), .Z(n7176) );
  BUF_X2 U6181 ( .A(n6107), .Z(n7279) );
  OAI222_X4 U6182 ( .A1(n7250), .A2(n6050), .B1(n5516), .B2(n7279), .C1(n6120), 
        .C2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n6144) );
  OAI222_X4 U6183 ( .A1(n7454), .A2(n6048), .B1(n5515), .B2(n7176), .C1(n6106), 
        .C2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n6132) );
  OR2_X2 U6184 ( .A1(n7277), .A2(n7653), .ZN(n7177) );
  AND2_X1 U6185 ( .A1(n7272), .A2(\Mcontrol/Operation_decoding32/N1987 ), .ZN(
        n7178) );
  AND3_X2 U6186 ( .A1(n6057), .A2(n7505), .A3(n7178), .ZN(n6097) );
  NAND2_X1 U6187 ( .A1(n7216), .A2(n7217), .ZN(
        \Mcontrol/Operation_decoding32/N1987 ) );
  NAND2_X4 U6188 ( .A1(n6040), .A2(\Mcontrol/Operation_decoding32/N1873 ), 
        .ZN(n6034) );
  NAND2_X4 U6189 ( .A1(\BYP_BRANCH_MUXB/N4 ), .A2(byp_controlB[0]), .ZN(n5527)
         );
  NOR2_X1 U6190 ( .A1(branch_rega[3]), .A2(n7381), .ZN(n7179) );
  NAND2_X1 U6191 ( .A1(\Mpath/the_alu/diff[30] ), .A2(n1698), .ZN(n7180) );
  NAND2_X1 U6192 ( .A1(\Mpath/the_alu/sum[30] ), .A2(n7634), .ZN(n7181) );
  AND2_X2 U6193 ( .A1(n7180), .A2(n7181), .ZN(n1907) );
  INV_X2 U6194 ( .A(\Mpath/the_alu/N59 ), .ZN(n7182) );
  OAI222_X4 U6195 ( .A1(n5549), .A2(n5523), .B1(n5550), .B2(n5525), .C1(n5551), 
        .C2(n5527), .ZN(branch_regb[30]) );
  INV_X1 U6196 ( .A(\exc[ALU_OFLOW1] ), .ZN(n7183) );
  NOR2_X1 U6197 ( .A1(n2494), .A2(n1845), .ZN(n7596) );
  INV_X4 U6198 ( .A(n7184), .ZN(n7185) );
  NAND2_X4 U6199 ( .A1(n6038), .A2(\Mcontrol/Operation_decoding32/N1873 ), 
        .ZN(n6020) );
  NAND2_X1 U6200 ( .A1(\Mpath/the_alu/N474 ), .A2(n2447), .ZN(n7186) );
  NAND2_X1 U6201 ( .A1(\Mpath/the_alu/N474 ), .A2(n2447), .ZN(n7187) );
  INV_X4 U6202 ( .A(n1692), .ZN(n1713) );
  NAND2_X1 U6203 ( .A1(n7188), .A2(\Mcontrol/st_logic/N95 ), .ZN(
        \Mcontrol/st_logic/N113 ) );
  AND3_X4 U6204 ( .A1(n7190), .A2(n7191), .A3(\Mcontrol/N34 ), .ZN(n7189) );
  INV_X32 U6205 ( .A(n7214), .ZN(n7190) );
  AND2_X2 U6206 ( .A1(\Mcontrol/m_sampled_xrd[2] ), .A2(n5503), .ZN(rd_addr[2]) );
  NOR4_X2 U6207 ( .A1(n2355), .A2(n2356), .A3(n2357), .A4(n2358), .ZN(n2354)
         );
  INV_X1 U6208 ( .A(\Mpath/the_alu/N64 ), .ZN(n7192) );
  NOR2_X1 U6209 ( .A1(byp_controlA[2]), .A2(\regfile/N264 ), .ZN(n7193) );
  NOR2_X1 U6210 ( .A1(byp_controlA[2]), .A2(\regfile/N264 ), .ZN(n7194) );
  BUF_X2 U6211 ( .A(n5633), .Z(n7611) );
  AND3_X4 U6212 ( .A1(n6425), .A2(rs1_addr[3]), .A3(n7382), .ZN(n5642) );
  INV_X1 U6213 ( .A(\regfile/N358 ), .ZN(\regfile/N455 ) );
  INV_X4 U6214 ( .A(n5640), .ZN(n2336) );
  AND4_X4 U6215 ( .A1(n1673), .A2(n2490), .A3(net56319), .A4(n6041), .ZN(
        net58101) );
  OR2_X1 U6216 ( .A1(\Alu_command[OP][4] ), .A2(\Alu_command[OP][5] ), .ZN(
        \Mpath/the_alu/N517 ) );
  OR2_X1 U6217 ( .A1(\Alu_command[OP][4] ), .A2(\Alu_command[OP][5] ), .ZN(
        \Mpath/the_alu/N460 ) );
  NAND2_X1 U6218 ( .A1(n7196), .A2(n7197), .ZN(\Mpath/the_alu/N448 ) );
  INV_X4 U6219 ( .A(n6512), .ZN(n7196) );
  XNOR2_X1 U6220 ( .A(\Mpath/the_alu/N21 ), .B(\Mpath/the_alu/sum[31] ), .ZN(
        n7197) );
  NAND4_X2 U6221 ( .A1(n6021), .A2(rs2_addr[1]), .A3(rs2_addr[0]), .A4(
        rs2_addr[2]), .ZN(n5754) );
  AND2_X1 U6222 ( .A1(\Mcontrol/Nextpc_decoding/Bta [18]), .A2(n1560), .ZN(
        n7244) );
  OAI21_X1 U6223 ( .B1(net56977), .B2(n6068), .A(n7310), .ZN(n7199) );
  OAI21_X1 U6224 ( .B1(n7596), .B2(n7437), .A(n7319), .ZN(n7198) );
  OAI21_X1 U6225 ( .B1(n7437), .B2(n7596), .A(n7049), .ZN(n6297) );
  NAND2_X1 U6226 ( .A1(\Mpath/the_alu/N93 ), .A2(n2454), .ZN(n7201) );
  NAND2_X1 U6227 ( .A1(\Mpath/the_alu/N91 ), .A2(n2455), .ZN(n7202) );
  AND2_X2 U6228 ( .A1(n7201), .A2(n7202), .ZN(n2453) );
  INV_X2 U6229 ( .A(\Mpath/the_alu/N503 ), .ZN(n2455) );
  NOR2_X1 U6230 ( .A1(\Mcontrol/Nextpc_decoding/N26 ), .A2(n6399), .ZN(n7204)
         );
  NOR2_X1 U6231 ( .A1(n7334), .A2(\Mcontrol/Nextpc_decoding/N325 ), .ZN(n7205)
         );
  INV_X1 U6232 ( .A(\Mcontrol/Nextpc_decoding/N324 ), .ZN(
        \Mcontrol/Nextpc_decoding/N325 ) );
  AND2_X1 U6233 ( .A1(n7628), .A2(n7629), .ZN(n6200) );
  AND2_X2 U6234 ( .A1(\Mcontrol/bp_logicB/N2 ), .A2(\Mcontrol/bp_logicB/N8 ), 
        .ZN(\Mcontrol/bp_logicB/N15 ) );
  INV_X1 U6235 ( .A(n5655), .ZN(n5549) );
  NOR2_X2 U6236 ( .A1(branch_rega[11]), .A2(branch_rega[12]), .ZN(n7593) );
  OAI222_X4 U6237 ( .A1(n5623), .A2(n5611), .B1(n7487), .B2(n2844), .C1(n5621), 
        .C2(n5609), .ZN(branch_rega[12]) );
  AND2_X1 U6238 ( .A1(n7206), .A2(n7256), .ZN(n7622) );
  NOR2_X1 U6239 ( .A1(n7098), .A2(n7425), .ZN(n7206) );
  AOI221_X4 U6240 ( .B1(n7351), .B2(n333), .C1(n6251), .C2(n331), .A(n330), 
        .ZN(n445) );
  INV_X1 U6241 ( .A(n7325), .ZN(n6434) );
  INV_X2 U6242 ( .A(n7277), .ZN(n7278) );
  NAND2_X1 U6243 ( .A1(\exc[DMEM_MISALIGN] ), .A2(\Scc_coproc/N575 ), .ZN(
        n7208) );
  AND2_X1 U6244 ( .A1(\exc[DMEM_MISALIGN] ), .A2(\exc[ALU_OFLOW1] ), .ZN(n1684) );
  OR3_X4 U6245 ( .A1(\regfile/N324 ), .A2(net55894), .A3(n1252), .ZN(n7209) );
  INV_X4 U6246 ( .A(n7209), .ZN(n317) );
  OR3_X4 U6247 ( .A1(\regfile/N318 ), .A2(net55890), .A3(n1108), .ZN(n7210) );
  INV_X4 U6248 ( .A(n7210), .ZN(n314) );
  NOR2_X1 U6249 ( .A1(n7634), .A2(n2452), .ZN(n7211) );
  NOR2_X1 U6250 ( .A1(n2453), .A2(n7212), .ZN(n2451) );
  INV_X1 U6251 ( .A(n7211), .ZN(n7212) );
  NAND2_X2 U6252 ( .A1(\Mpath/the_alu/N515 ), .A2(\Mpath/the_alu/N509 ), .ZN(
        n2452) );
  OR2_X2 U6253 ( .A1(n7403), .A2(\Mcontrol/Operation_decoding32/N1880 ), .ZN(
        \Mcontrol/Operation_decoding32/N1881 ) );
  NOR4_X2 U6254 ( .A1(n2849), .A2(n2850), .A3(n2851), .A4(n2852), .ZN(n2848)
         );
  AND2_X4 U6255 ( .A1(n6433), .A2(n7686), .ZN(n6429) );
  NOR2_X1 U6256 ( .A1(\Mcontrol/Operation_decoding32/N1984 ), .A2(n7308), .ZN(
        n7216) );
  NOR2_X1 U6257 ( .A1(n7305), .A2(n7447), .ZN(n7217) );
  CLKBUF_X1 U6258 ( .A(\Mcontrol/Operation_decoding32/N1957 ), .Z(n7218) );
  NOR2_X1 U6259 ( .A1(n7403), .A2(n7088), .ZN(n7219) );
  NAND2_X1 U6260 ( .A1(n7219), .A2(n7220), .ZN(n7505) );
  AND2_X1 U6261 ( .A1(net58000), .A2(n7221), .ZN(n7220) );
  INV_X1 U6262 ( .A(net56678), .ZN(net58000) );
  INV_X1 U6263 ( .A(\Mcontrol/d_instr [28]), .ZN(
        \Mcontrol/Operation_decoding32/N1989 ) );
  AND2_X1 U6264 ( .A1(n7263), .A2(n7652), .ZN(n7431) );
  INV_X2 U6265 ( .A(n7194), .ZN(n7487) );
  NAND2_X1 U6266 ( .A1(\Mcontrol/bp_logicA/memory_main ), .A2(n2488), .ZN(
        \Mcontrol/st_logic/N47 ) );
  AND3_X4 U6267 ( .A1(n7173), .A2(n7686), .A3(n6431), .ZN(n7642) );
  NOR2_X1 U6268 ( .A1(n7686), .A2(n7173), .ZN(n6428) );
  NAND2_X1 U6269 ( .A1(n7522), .A2(n7403), .ZN(n7398) );
  NOR2_X1 U6270 ( .A1(n7165), .A2(n7093), .ZN(n7420) );
  INV_X1 U6271 ( .A(n1509), .ZN(n7222) );
  NAND3_X2 U6272 ( .A1(n7598), .A2(net57341), .A3(n1474), .ZN(n1523) );
  NAND2_X1 U6273 ( .A1(n7146), .A2(n7223), .ZN(n7414) );
  AND2_X1 U6274 ( .A1(n7043), .A2(n7053), .ZN(n7223) );
  INV_X1 U6275 ( .A(n2774), .ZN(n7224) );
  OAI22_X1 U6276 ( .A1(n6093), .A2(n5914), .B1(n6200), .B2(n6171), .ZN(n6199)
         );
  AND2_X2 U6277 ( .A1(n7135), .A2(n7438), .ZN(n7424) );
  NAND2_X1 U6278 ( .A1(n7224), .A2(n7047), .ZN(n7226) );
  CLKBUF_X1 U6279 ( .A(n7165), .Z(n7227) );
  NOR2_X1 U6280 ( .A1(n7446), .A2(net56922), .ZN(n7228) );
  NOR2_X1 U6281 ( .A1(n7058), .A2(n7088), .ZN(
        \Mcontrol/Operation_decoding32/N2001 ) );
  NAND2_X1 U6282 ( .A1(n7146), .A2(n7078), .ZN(n7551) );
  OR2_X1 U6283 ( .A1(\Mcontrol/Operation_decoding32/N1922 ), .A2(n7513), .ZN(
        net57313) );
  INV_X1 U6284 ( .A(net57810), .ZN(n6054) );
  INV_X1 U6285 ( .A(n6076), .ZN(n7229) );
  INV_X1 U6286 ( .A(n7647), .ZN(n7230) );
  NAND2_X1 U6287 ( .A1(\Mcontrol/Operation_decoding32/N1975 ), .A2(
        \Mcontrol/Operation_decoding32/N89 ), .ZN(n7231) );
  NAND3_X1 U6288 ( .A1(net57942), .A2(n7232), .A3(n6059), .ZN(n7442) );
  INV_X1 U6289 ( .A(n7231), .ZN(n7232) );
  INV_X1 U6290 ( .A(n7177), .ZN(n7462) );
  CLKBUF_X1 U6291 ( .A(n7551), .Z(n7233) );
  OR2_X1 U6292 ( .A1(n7160), .A2(\Mcontrol/d_instr [28]), .ZN(n7234) );
  NOR2_X1 U6293 ( .A1(n7544), .A2(n6068), .ZN(net57942) );
  CLKBUF_X1 U6294 ( .A(n7250), .Z(n7454) );
  OR2_X2 U6295 ( .A1(n7124), .A2(n6956), .ZN(n7426) );
  NAND3_X1 U6296 ( .A1(\Mcontrol/Operation_decoding32/N2036 ), .A2(n7301), 
        .A3(\Mcontrol/Operation_decoding32/N2030 ), .ZN(n7235) );
  NAND3_X1 U6297 ( .A1(\Mcontrol/Operation_decoding32/N2036 ), .A2(n7301), 
        .A3(\Mcontrol/Operation_decoding32/N2030 ), .ZN(n6063) );
  INV_X1 U6298 ( .A(n1471), .ZN(n7236) );
  NOR2_X2 U6299 ( .A1(n7237), .A2(n7238), .ZN(n7580) );
  OR2_X1 U6300 ( .A1(n7239), .A2(branch_rega[1]), .ZN(n7238) );
  INV_X1 U6301 ( .A(n7445), .ZN(n7239) );
  OR2_X1 U6302 ( .A1(n7241), .A2(branch_rega[7]), .ZN(n7240) );
  INV_X1 U6303 ( .A(n7444), .ZN(n7241) );
  CLKBUF_X1 U6304 ( .A(n7873), .Z(I_ADDR_OUTBUS[18]) );
  AND2_X1 U6305 ( .A1(jar_in[18]), .A2(n1561), .ZN(n7245) );
  NOR3_X2 U6306 ( .A1(n7243), .A2(n7244), .A3(n7245), .ZN(n2735) );
  NAND2_X1 U6307 ( .A1(n7041), .A2(n7435), .ZN(n7247) );
  AND3_X2 U6308 ( .A1(n7677), .A2(n7678), .A3(n7679), .ZN(
        \Mcontrol/bp_logicA/N3 ) );
  OR2_X1 U6309 ( .A1(branch_rega[21]), .A2(branch_rega[20]), .ZN(n7662) );
  OAI222_X1 U6310 ( .A1(n5623), .A2(n5578), .B1(n7486), .B2(n2666), .C1(n5621), 
        .C2(n5576), .ZN(branch_rega[22]) );
  AOI221_X1 U6311 ( .B1(n371), .B2(\Mcontrol/f_currpc[4] ), .C1(n372), .C2(
        I_ADDR_OUTBUS[4]), .A(n373), .ZN(n837) );
  NAND2_X1 U6312 ( .A1(net56765), .A2(n7248), .ZN(
        \Mcontrol/Operation_decoding32/N1951 ) );
  AND2_X1 U6313 ( .A1(n7419), .A2(n7401), .ZN(n7248) );
  OAI222_X1 U6314 ( .A1(n7454), .A2(n5846), .B1(n6106), .B2(n7176), .C1(n5904), 
        .C2(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n6104) );
  OR2_X2 U6315 ( .A1(n7060), .A2(n7536), .ZN(
        \Mcontrol/Operation_decoding32/N2021 ) );
  OR2_X1 U6316 ( .A1(\Mcontrol/d_jump_type[1] ), .A2(\Mcontrol/st_logic/N74 ), 
        .ZN(\Mcontrol/st_logic/N75 ) );
  OR2_X1 U6317 ( .A1(\Mcontrol/st_logic/N58 ), .A2(\Mcontrol/st_logic/N73 ), 
        .ZN(\Mcontrol/st_logic/N74 ) );
  XNOR2_X1 U6318 ( .A(n7249), .B(n7658), .ZN(n7280) );
  INV_X32 U6319 ( .A(\Mpath/the_alu/N21 ), .ZN(n7249) );
  NAND4_X1 U6320 ( .A1(n1844), .A2(\Mcontrol/Operation_decoding32/N89 ), .A3(
        n6059), .A4(\Mcontrol/Operation_decoding32/N1975 ), .ZN(n7250) );
  INV_X1 U6321 ( .A(n7263), .ZN(n7252) );
  NOR3_X1 U6322 ( .A1(\Mcontrol/Operation_decoding32/N2001 ), .A2(n7453), .A3(
        \Mcontrol/Operation_decoding32/N2007 ), .ZN(n6057) );
  NOR2_X4 U6323 ( .A1(n7675), .A2(rs1_addr[4]), .ZN(n6433) );
  OR2_X2 U6324 ( .A1(n7673), .A2(n7631), .ZN(n7254) );
  AND2_X4 U6325 ( .A1(\Mcontrol/d_sampled_finstr [26]), .A2(n7278), .ZN(
        \Mcontrol/d_instr [26]) );
  INV_X1 U6326 ( .A(n7225), .ZN(n1471) );
  CLKBUF_X1 U6327 ( .A(n7250), .Z(n7255) );
  INV_X4 U6328 ( .A(n7256), .ZN(\Mcontrol/d_instr [28]) );
  NAND2_X1 U6329 ( .A1(n7258), .A2(n7464), .ZN(n7257) );
  AND2_X2 U6330 ( .A1(n7680), .A2(n7689), .ZN(n7258) );
  NAND2_X1 U6331 ( .A1(n371), .A2(\Mcontrol/f_currpc[8] ), .ZN(n7259) );
  NAND2_X1 U6332 ( .A1(n372), .A2(I_ADDR_OUTBUS[8]), .ZN(n7260) );
  INV_X1 U6333 ( .A(n373), .ZN(n7261) );
  AND3_X1 U6334 ( .A1(n7259), .A2(n7260), .A3(n7261), .ZN(n826) );
  OR2_X2 U6335 ( .A1(n7267), .A2(n7580), .ZN(\Mcontrol/Nextpc_decoding/N31 )
         );
  NAND2_X1 U6336 ( .A1(n7198), .A2(\Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n7262) );
  OR2_X1 U6337 ( .A1(\Mpath/out_regA[4] ), .A2(n7707), .ZN(
        \Mpath/the_alu/N153 ) );
  AND2_X1 U6338 ( .A1(\Mpath/out_regA[4] ), .A2(n7707), .ZN(
        \Mpath/the_alu/N121 ) );
  NOR2_X4 U6339 ( .A1(n1523), .A2(n7159), .ZN(n1533) );
  OR2_X2 U6340 ( .A1(n7252), .A2(n7462), .ZN(
        \Mcontrol/Operation_decoding32/N2062 ) );
  INV_X1 U6341 ( .A(n7469), .ZN(n7264) );
  INV_X1 U6342 ( .A(net56617), .ZN(net57843) );
  CLKBUF_X1 U6343 ( .A(n7881), .Z(I_ADDR_OUTBUS[10]) );
  CLKBUF_X1 U6344 ( .A(n7086), .Z(n7267) );
  AND2_X1 U6345 ( .A1(n6102), .A2(n6515), .ZN(n7268) );
  AND2_X1 U6346 ( .A1(\Mcontrol/Nextpc_decoding/Bta [10]), .A2(net58826), .ZN(
        n7269) );
  AND2_X1 U6347 ( .A1(jar_in[10]), .A2(n1561), .ZN(n7270) );
  NOR3_X2 U6348 ( .A1(n7268), .A2(n7269), .A3(n7270), .ZN(n2876) );
  OR3_X2 U6349 ( .A1(\regfile/N360 ), .A2(net55894), .A3(n1251), .ZN(n7271) );
  INV_X4 U6350 ( .A(n7271), .ZN(n252) );
  NAND3_X1 U6351 ( .A1(n7273), .A2(n7052), .A3(n7305), .ZN(n7272) );
  NAND2_X1 U6352 ( .A1(net56996), .A2(\Mcontrol/d_instr [7]), .ZN(n7274) );
  NAND2_X1 U6353 ( .A1(net56605), .A2(n7275), .ZN(n2459) );
  INV_X1 U6354 ( .A(n7274), .ZN(n7275) );
  INV_X2 U6355 ( .A(n6106), .ZN(\Mcontrol/d_instr [7]) );
  CLKBUF_X1 U6356 ( .A(n6080), .Z(net56605) );
  OR3_X4 U6357 ( .A1(\regfile/N415 ), .A2(net55890), .A3(n1108), .ZN(n7276) );
  INV_X4 U6358 ( .A(n7276), .ZN(n278) );
  OAI222_X4 U6359 ( .A1(n5567), .A2(n5621), .B1(n5512), .B2(n7486), .C1(n5569), 
        .C2(n5623), .ZN(branch_rega[25]) );
  NAND2_X1 U6360 ( .A1(n6297), .A2(\Mcontrol/Operation_decoding32/N1975 ), 
        .ZN(n6107) );
  OAI222_X4 U6361 ( .A1(n5570), .A2(n5621), .B1(n5513), .B2(n7486), .C1(n5572), 
        .C2(n5623), .ZN(branch_rega[24]) );
  AND3_X1 U6362 ( .A1(n7870), .A2(n7869), .A3(n7868), .ZN(n7677) );
  OAI222_X4 U6363 ( .A1(n5558), .A2(n5621), .B1(n5509), .B2(n7486), .C1(n5560), 
        .C2(n5623), .ZN(branch_rega[28]) );
  OAI222_X1 U6364 ( .A1(n5623), .A2(n5602), .B1(n7486), .B2(n2793), .C1(n5621), 
        .C2(n5600), .ZN(branch_rega[15]) );
  NAND2_X1 U6365 ( .A1(n7541), .A2(n7542), .ZN(
        \Mcontrol/Operation_decoding32/N1939 ) );
  INV_X1 U6366 ( .A(n7671), .ZN(n7282) );
  CLKBUF_X1 U6367 ( .A(n7882), .Z(I_ADDR_OUTBUS[9]) );
  AND2_X1 U6368 ( .A1(n6102), .A2(n6536), .ZN(n7284) );
  AND2_X1 U6369 ( .A1(\Mcontrol/Nextpc_decoding/Bta [9]), .A2(n1560), .ZN(
        n7285) );
  AND2_X1 U6370 ( .A1(jar_in[9]), .A2(n1561), .ZN(n7286) );
  NOR3_X2 U6371 ( .A1(n7284), .A2(n7285), .A3(n7286), .ZN(n2506) );
  OR2_X1 U6372 ( .A1(n7100), .A2(n7287), .ZN(n5517) );
  NOR2_X2 U6373 ( .A1(n6022), .A2(rs2_addr[1]), .ZN(n6025) );
  OR2_X1 U6374 ( .A1(rs2_addr[1]), .A2(\regfile/N266 ), .ZN(\regfile/N267 ) );
  NOR2_X2 U6375 ( .A1(n7636), .A2(n7089), .ZN(n7289) );
  CLKBUF_X1 U6376 ( .A(n7883), .Z(I_ADDR_OUTBUS[7]) );
  AND2_X1 U6377 ( .A1(n2447), .A2(\Mpath/the_alu/N473 ), .ZN(n1710) );
  AND3_X4 U6378 ( .A1(n7292), .A2(net57757), .A3(n7291), .ZN(n237) );
  NOR2_X1 U6379 ( .A1(rd_addr[2]), .A2(\regfile/N329 ), .ZN(n7292) );
  INV_X1 U6380 ( .A(\Mpath/the_alu/N473 ), .ZN(\Mpath/the_alu/N474 ) );
  AND2_X1 U6381 ( .A1(n1697), .A2(n6512), .ZN(n7295) );
  AND2_X1 U6382 ( .A1(\Mpath/the_alu/diff[31] ), .A2(n1698), .ZN(n7296) );
  NOR3_X2 U6383 ( .A1(n7294), .A2(n7295), .A3(n7296), .ZN(n1685) );
  CLKBUF_X1 U6384 ( .A(n7884), .Z(I_ADDR_OUTBUS[6]) );
  CLKBUF_X1 U6385 ( .A(n7267), .Z(n7298) );
  OAI222_X1 U6386 ( .A1(n5546), .A2(n5621), .B1(n5506), .B2(n7485), .C1(n5548), 
        .C2(n5623), .ZN(branch_rega[31]) );
  NAND2_X1 U6387 ( .A1(\Mcontrol/d_instr [27]), .A2(\Mcontrol/d_instr [28]), 
        .ZN(n7299) );
  NAND2_X1 U6388 ( .A1(n7300), .A2(n7052), .ZN(
        \Mcontrol/Operation_decoding32/N1968 ) );
  NAND2_X1 U6389 ( .A1(n7256), .A2(n7409), .ZN(n7302) );
  NOR2_X1 U6390 ( .A1(\Mcontrol/d_instr [26]), .A2(n7041), .ZN(n7304) );
  OR2_X1 U6391 ( .A1(n7451), .A2(n7547), .ZN(net57730) );
  INV_X1 U6392 ( .A(n7053), .ZN(n7305) );
  NAND2_X1 U6393 ( .A1(n7306), .A2(\Mcontrol/d_instr [28]), .ZN(
        \Mcontrol/Operation_decoding32/N2064 ) );
  NOR2_X1 U6394 ( .A1(\Mcontrol/Operation_decoding32/N2062 ), .A2(n7536), .ZN(
        n7306) );
  INV_X1 U6395 ( .A(\Mcontrol/Operation_decoding32/N1989 ), .ZN(n7308) );
  AND2_X1 U6396 ( .A1(n7383), .A2(n7452), .ZN(n7309) );
  AND2_X1 U6397 ( .A1(\Mcontrol/Operation_decoding32/N1922 ), .A2(n7072), .ZN(
        n7383) );
  INV_X1 U6398 ( .A(branch_rega[6]), .ZN(n7489) );
  AND2_X1 U6399 ( .A1(\Mpath/out_regA[0] ), .A2(n7715), .ZN(
        \Mpath/the_alu/N125 ) );
  OR2_X1 U6400 ( .A1(\Mpath/out_regA[0] ), .A2(n7715), .ZN(
        \Mpath/the_alu/N157 ) );
  INV_X1 U6401 ( .A(n7162), .ZN(n7310) );
  CLKBUF_X1 U6402 ( .A(break_code[3]), .Z(n7311) );
  AOI21_X1 U6403 ( .B1(n6401), .B2(n6402), .A(n6403), .ZN(n6400) );
  INV_X1 U6404 ( .A(n7310), .ZN(n6067) );
  OR2_X1 U6405 ( .A1(\Mpath/out_regA[2] ), .A2(n7711), .ZN(
        \Mpath/the_alu/N155 ) );
  AND2_X1 U6406 ( .A1(\Mpath/out_regA[2] ), .A2(n7711), .ZN(
        \Mpath/the_alu/N123 ) );
  AND2_X2 U6407 ( .A1(n7676), .A2(n7312), .ZN(n7661) );
  NOR2_X1 U6408 ( .A1(branch_rega[11]), .A2(n7354), .ZN(n7312) );
  INV_X1 U6409 ( .A(n1694), .ZN(n7313) );
  INV_X1 U6410 ( .A(n1695), .ZN(n7314) );
  INV_X1 U6411 ( .A(n7314), .ZN(n7315) );
  OR2_X2 U6412 ( .A1(n7474), .A2(n7355), .ZN(n7354) );
  INV_X2 U6413 ( .A(n1694), .ZN(n1714) );
  AND3_X4 U6414 ( .A1(n7317), .A2(net57683), .A3(n7316), .ZN(n292) );
  INV_X32 U6415 ( .A(net55892), .ZN(net57683) );
  NOR2_X1 U6416 ( .A1(rd_addr[2]), .A2(\regfile/N279 ), .ZN(n7317) );
  OR2_X1 U6417 ( .A1(\Mpath/the_alu/N453 ), .A2(\Alu_command[OP][5] ), .ZN(
        \Mpath/the_alu/N505 ) );
  OR2_X1 U6418 ( .A1(\Mpath/the_alu/N453 ), .A2(\Alu_command[OP][5] ), .ZN(
        \Mpath/the_alu/N511 ) );
  OR2_X1 U6419 ( .A1(\Mpath/the_alu/N453 ), .A2(\Mpath/the_alu/N466 ), .ZN(
        \Mpath/the_alu/N487 ) );
  OR2_X1 U6420 ( .A1(\Mpath/the_alu/N453 ), .A2(\Mpath/the_alu/N466 ), .ZN(
        \Mpath/the_alu/N481 ) );
  OR2_X1 U6421 ( .A1(\Mpath/the_alu/N453 ), .A2(\Mpath/the_alu/N466 ), .ZN(
        \Mpath/the_alu/N475 ) );
  OR3_X2 U6422 ( .A1(\regfile/N336 ), .A2(net55896), .A3(n1251), .ZN(n7318) );
  INV_X4 U6423 ( .A(n7318), .ZN(n240) );
  OR2_X1 U6424 ( .A1(\regfile/N315 ), .A2(n7195), .ZN(\regfile/N456 ) );
  OR2_X1 U6425 ( .A1(\regfile/N315 ), .A2(n7195), .ZN(\regfile/N438 ) );
  OR2_X1 U6426 ( .A1(\regfile/N315 ), .A2(n7195), .ZN(\regfile/N444 ) );
  OR2_X1 U6427 ( .A1(\regfile/N315 ), .A2(n7195), .ZN(\regfile/N414 ) );
  OR2_X1 U6428 ( .A1(\regfile/N315 ), .A2(\regfile/N455 ), .ZN(\regfile/N420 )
         );
  OR2_X1 U6429 ( .A1(\regfile/N315 ), .A2(\regfile/N455 ), .ZN(\regfile/N426 )
         );
  OR2_X1 U6430 ( .A1(\regfile/N315 ), .A2(\regfile/N455 ), .ZN(\regfile/N432 )
         );
  AND2_X1 U6431 ( .A1(\Mpath/out_regA[22] ), .A2(\Mpath/out_regB[22] ), .ZN(
        \Mpath/the_alu/N103 ) );
  OR2_X1 U6432 ( .A1(\Mpath/out_regA[22] ), .A2(\Mpath/out_regB[22] ), .ZN(
        \Mpath/the_alu/N135 ) );
  AND2_X2 U6433 ( .A1(\Mcontrol/Operation_decoding32/N1969 ), .A2(
        \Mcontrol/Operation_decoding32/N1963 ), .ZN(n7319) );
  NOR2_X2 U6434 ( .A1(n1710), .A2(n7313), .ZN(n1695) );
  NOR2_X1 U6435 ( .A1(n7600), .A2(n7459), .ZN(n7320) );
  AOI22_X2 U6436 ( .A1(n7503), .A2(\regfile/reg_out[21][22] ), .B1(n7612), 
        .B2(\regfile/reg_out[20][22] ), .ZN(n6229) );
  NOR2_X1 U6437 ( .A1(n7352), .A2(n7673), .ZN(n7351) );
  NOR2_X4 U6438 ( .A1(n2500), .A2(\Mcontrol/Operation_decoding32/N1976 ), .ZN(
        n1673) );
  INV_X2 U6439 ( .A(n2792), .ZN(n1474) );
  NAND2_X2 U6440 ( .A1(n1533), .A2(n7430), .ZN(n2500) );
  INV_X1 U6441 ( .A(branch_rega[15]), .ZN(n7650) );
  AOI221_X4 U6442 ( .B1(n7623), .B2(n333), .C1(n6239), .C2(n331), .A(n330), 
        .ZN(n410) );
  OR2_X1 U6443 ( .A1(\Mcontrol/Operation_decoding32/N1900 ), .A2(n7623), .ZN(
        \Mcontrol/Operation_decoding32/N1902 ) );
  AND2_X2 U6444 ( .A1(\Mcontrol/bp_logicA/N3 ), .A2(\Mcontrol/bp_logicA/N13 ), 
        .ZN(\Mcontrol/bp_logicA/N16 ) );
  NAND4_X1 U6445 ( .A1(n6417), .A2(rs1_addr[1]), .A3(rs1_addr[0]), .A4(
        rs1_addr[2]), .ZN(n5629) );
  INV_X1 U6446 ( .A(\Mpath/out_regB[18] ), .ZN(n7358) );
  INV_X1 U6447 ( .A(n7692), .ZN(n7693) );
  OAI222_X1 U6448 ( .A1(n5623), .A2(n5530), .B1(n7487), .B2(n2527), .C1(n5621), 
        .C2(n5528), .ZN(branch_rega[8]) );
  NOR2_X4 U6449 ( .A1(n1916), .A2(\Mpath/the_shift/N118 ), .ZN(n1704) );
  INV_X1 U6450 ( .A(n7556), .ZN(n7557) );
  INV_X2 U6451 ( .A(\Mpath/out_regB[15] ), .ZN(n7321) );
  INV_X1 U6452 ( .A(n7321), .ZN(n7322) );
  INV_X2 U6453 ( .A(n7321), .ZN(n7323) );
  CLKBUF_X1 U6454 ( .A(byp_controlA[0]), .Z(n7324) );
  NAND2_X2 U6455 ( .A1(n7645), .A2(\Mcontrol/Operation_decoding32/N1887 ), 
        .ZN(n7326) );
  NAND2_X1 U6456 ( .A1(n7645), .A2(\Mcontrol/Operation_decoding32/N1887 ), 
        .ZN(n7325) );
  INV_X1 U6457 ( .A(\Mcontrol/st_logic/N47 ), .ZN(byp_controlA[0]) );
  NOR2_X4 U6458 ( .A1(n7569), .A2(\Mcontrol/Operation_decoding32/N1881 ), .ZN(
        n7645) );
  NAND2_X1 U6459 ( .A1(n7645), .A2(\Mcontrol/Operation_decoding32/N1887 ), 
        .ZN(\Mcontrol/Operation_decoding32/N1871 ) );
  NOR2_X1 U6460 ( .A1(n7686), .A2(rs1_addr[2]), .ZN(n7328) );
  NOR2_X1 U6461 ( .A1(n7686), .A2(rs1_addr[2]), .ZN(n7327) );
  NOR2_X1 U6462 ( .A1(n7686), .A2(rs1_addr[2]), .ZN(n6426) );
  NOR2_X2 U6463 ( .A1(n7329), .A2(\Mcontrol/x_sampled_dwe ), .ZN(
        \Mcontrol/bp_logicA/exec_main ) );
  NAND2_X1 U6464 ( .A1(\Mcontrol/bp_logicA/N2 ), .A2(\Mcontrol/bp_logicA/N8 ), 
        .ZN(n7329) );
  NAND2_X4 U6465 ( .A1(\Mcontrol/Operation_decoding32/N1873 ), .A2(n6041), 
        .ZN(n6026) );
  OR2_X4 U6466 ( .A1(\BYP_BRANCH_MUXB/N4 ), .A2(\regfile/N269 ), .ZN(n5525) );
  INV_X2 U6467 ( .A(\Mpath/out_regB[19] ), .ZN(n7330) );
  INV_X1 U6468 ( .A(n7330), .ZN(n7331) );
  INV_X1 U6469 ( .A(n7330), .ZN(n7333) );
  INV_X1 U6470 ( .A(n7330), .ZN(n7332) );
  INV_X4 U6471 ( .A(n1252), .ZN(n7368) );
  OR3_X1 U6472 ( .A1(\regfile/N397 ), .A2(net55896), .A3(n1252), .ZN(n7406) );
  OR2_X1 U6473 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N460 ), .ZN(
        \Mpath/the_alu/N461 ) );
  OR2_X1 U6474 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N454 ), .ZN(
        \Mpath/the_alu/N455 ) );
  OR2_X1 U6475 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N469 ), .ZN(
        \Mpath/the_alu/N470 ) );
  OR2_X1 U6476 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N475 ), .ZN(
        \Mpath/the_alu/N476 ) );
  OR2_X1 U6477 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N481 ), .ZN(
        \Mpath/the_alu/N482 ) );
  OR2_X1 U6478 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N493 ), .ZN(
        \Mpath/the_alu/N494 ) );
  OR2_X1 U6479 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N487 ), .ZN(
        \Mpath/the_alu/N488 ) );
  OR2_X1 U6480 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N499 ), .ZN(
        \Mpath/the_alu/N500 ) );
  OR2_X1 U6481 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N511 ), .ZN(
        \Mpath/the_alu/N512 ) );
  OR2_X1 U6482 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N505 ), .ZN(
        \Mpath/the_alu/N506 ) );
  OR2_X1 U6483 ( .A1(\Alu_command[OP][3] ), .A2(\Mpath/the_alu/N517 ), .ZN(
        \Mpath/the_alu/N518 ) );
  INV_X4 U6484 ( .A(n1108), .ZN(n7439) );
  OR3_X4 U6485 ( .A1(\regfile/N342 ), .A2(net55892), .A3(n1108), .ZN(n7370) );
  OR2_X1 U6486 ( .A1(\Mcontrol/d_instr [3]), .A2(
        \Mcontrol/Operation_decoding32/N1902 ), .ZN(
        \Mcontrol/Operation_decoding32/N1903 ) );
  OR2_X1 U6487 ( .A1(n7324), .A2(\Mcontrol/st_logic/N55 ), .ZN(
        \Mcontrol/st_logic/N18 ) );
  OR2_X1 U6488 ( .A1(byp_controlA[0]), .A2(\Mcontrol/st_logic/N55 ), .ZN(
        \Mcontrol/st_logic/N56 ) );
  OR2_X1 U6489 ( .A1(\Mcontrol/st_logic/N47 ), .A2(\Mcontrol/st_logic/N55 ), 
        .ZN(\Mcontrol/st_logic/N49 ) );
  OR2_X1 U6490 ( .A1(\Mcontrol/d_instr [3]), .A2(
        \Mcontrol/Operation_decoding32/N1908 ), .ZN(
        \Mcontrol/Operation_decoding32/N1909 ) );
  AND2_X1 U6491 ( .A1(\Mcontrol/d_instr [3]), .A2(
        \Mcontrol/Operation_decoding32/N1894 ), .ZN(
        \Mcontrol/Operation_decoding32/N1895 ) );
  NAND2_X2 U6492 ( .A1(n6499), .A2(n6501), .ZN(n6500) );
  NOR2_X2 U6493 ( .A1(n7173), .A2(rs1_addr[1]), .ZN(n7382) );
  INV_X2 U6494 ( .A(n7500), .ZN(n7502) );
  AOI21_X1 U6495 ( .B1(n7154), .B2(n6402), .A(n6403), .ZN(n7334) );
  AND2_X4 U6496 ( .A1(n6429), .A2(n7382), .ZN(n5649) );
  AND2_X1 U6497 ( .A1(\Mcontrol/st_logic/N57 ), .A2(\Mcontrol/st_logic/N51 ), 
        .ZN(\Mcontrol/st_logic/N118 ) );
  OAI21_X1 U6498 ( .B1(n6067), .B2(n2499), .A(n1673), .ZN(
        \Mcontrol/d_jump_type[0] ) );
  OAI21_X2 U6499 ( .B1(n5743), .B2(n2493), .A(n1673), .ZN(
        \Mcontrol/d_jump_type[2] ) );
  INV_X4 U6500 ( .A(branch_rega[22]), .ZN(net56617) );
  AND2_X4 U6501 ( .A1(\Mcontrol/m_sampled_xrd[3] ), .A2(n5503), .ZN(rd_addr[3]) );
  CLKBUF_X1 U6502 ( .A(n7875), .Z(I_ADDR_OUTBUS[16]) );
  AND2_X1 U6503 ( .A1(n6102), .A2(n6534), .ZN(n7336) );
  AND2_X1 U6504 ( .A1(\Mcontrol/Nextpc_decoding/Bta [16]), .A2(net58826), .ZN(
        n7337) );
  AND2_X1 U6505 ( .A1(jar_in[16]), .A2(n1561), .ZN(n7338) );
  NOR3_X2 U6506 ( .A1(n7336), .A2(n7337), .A3(n7338), .ZN(n2771) );
  AND2_X1 U6507 ( .A1(n6102), .A2(n6528), .ZN(n7339) );
  AND2_X1 U6508 ( .A1(\Mcontrol/Nextpc_decoding/Bta [19]), .A2(net58826), .ZN(
        n7340) );
  AND2_X1 U6509 ( .A1(jar_in[19]), .A2(n1561), .ZN(n7341) );
  INV_X1 U6510 ( .A(\Mpath/out_regB[17] ), .ZN(n7342) );
  INV_X1 U6511 ( .A(n7342), .ZN(n7343) );
  INV_X2 U6512 ( .A(n7342), .ZN(n7344) );
  OAI222_X4 U6513 ( .A1(n5523), .A2(n5546), .B1(n5547), .B2(n5525), .C1(n5548), 
        .C2(n5527), .ZN(branch_regb[31]) );
  OAI221_X4 U6514 ( .B1(net55834), .B2(n3052), .C1(n5517), .C2(net55918), .A(
        n1456), .ZN(n4371) );
  OAI221_X4 U6515 ( .B1(n2500), .B2(n2717), .C1(n5517), .C2(n2718), .A(n2719), 
        .ZN(break_code[19]) );
  INV_X4 U6516 ( .A(branch_rega[27]), .ZN(n7349) );
  CLKBUF_X1 U6517 ( .A(n7872), .Z(I_ADDR_OUTBUS[20]) );
  NAND2_X1 U6518 ( .A1(\Mcontrol/Nextpc_decoding/Bta [20]), .A2(net58826), 
        .ZN(n7347) );
  NAND2_X1 U6519 ( .A1(n1561), .A2(jar_in[20]), .ZN(n7348) );
  AND3_X2 U6520 ( .A1(n7346), .A2(n7347), .A3(n7348), .ZN(n2698) );
  NOR3_X4 U6521 ( .A1(\Mpath/the_alu/N486 ), .A2(n6500), .A3(
        \Mpath/the_alu/N480 ), .ZN(n2447) );
  INV_X1 U6522 ( .A(n5913), .ZN(n7703) );
  CLKBUF_X1 U6523 ( .A(break_code[2]), .Z(n7353) );
  INV_X1 U6524 ( .A(n7371), .ZN(n7355) );
  AND2_X1 U6525 ( .A1(\Mcontrol/Nextpc_decoding/Bta [11]), .A2(n1560), .ZN(
        n7701) );
  INV_X1 U6526 ( .A(n7358), .ZN(n7359) );
  INV_X1 U6527 ( .A(n7358), .ZN(n7361) );
  INV_X1 U6528 ( .A(n7358), .ZN(n7360) );
  OR3_X2 U6529 ( .A1(\regfile/N409 ), .A2(net55896), .A3(n1251), .ZN(n7363) );
  INV_X4 U6530 ( .A(n7363), .ZN(n275) );
  AND3_X4 U6531 ( .A1(n7365), .A2(net57474), .A3(n7364), .ZN(n272) );
  INV_X32 U6532 ( .A(net55888), .ZN(net57474) );
  NOR2_X1 U6533 ( .A1(\regfile/N290 ), .A2(\regfile/N402 ), .ZN(n7365) );
  AOI21_X1 U6534 ( .B1(\Mcontrol/Nextpc_decoding/condition ), .B2(
        \Mcontrol/st_logic/N103 ), .A(\Mcontrol/d_jump_type[3] ), .ZN(n6398)
         );
  OR2_X2 U6535 ( .A1(branch_rega[30]), .A2(branch_rega[31]), .ZN(
        \Mcontrol/Nextpc_decoding/N252 ) );
  OR2_X4 U6536 ( .A1(branch_rega[20]), .A2(branch_rega[19]), .ZN(n7694) );
  INV_X4 U6537 ( .A(n5629), .ZN(n2334) );
  OR2_X1 U6538 ( .A1(rd_addr[3]), .A2(n7195), .ZN(\regfile/N396 ) );
  OR2_X1 U6539 ( .A1(rd_addr[3]), .A2(n7195), .ZN(\regfile/N390 ) );
  OR2_X1 U6540 ( .A1(rd_addr[3]), .A2(\regfile/N455 ), .ZN(\regfile/N384 ) );
  OR2_X1 U6541 ( .A1(rd_addr[3]), .A2(\regfile/N455 ), .ZN(\regfile/N372 ) );
  OR2_X1 U6542 ( .A1(rd_addr[3]), .A2(\regfile/N455 ), .ZN(\regfile/N378 ) );
  OR2_X1 U6543 ( .A1(rd_addr[3]), .A2(n7195), .ZN(\regfile/N366 ) );
  OR2_X1 U6544 ( .A1(rd_addr[3]), .A2(n7195), .ZN(\regfile/N402 ) );
  AND3_X4 U6545 ( .A1(n7367), .A2(net57465), .A3(n7366), .ZN(n249) );
  NOR2_X1 U6546 ( .A1(\regfile/N290 ), .A2(\regfile/N353 ), .ZN(n7367) );
  AND3_X4 U6547 ( .A1(n7369), .A2(net57460), .A3(n7368), .ZN(n246) );
  INV_X32 U6548 ( .A(net55896), .ZN(net57460) );
  NOR2_X1 U6549 ( .A1(\regfile/N290 ), .A2(\regfile/N347 ), .ZN(n7369) );
  INV_X4 U6550 ( .A(n7370), .ZN(n243) );
  NOR2_X1 U6551 ( .A1(n7473), .A2(branch_rega[7]), .ZN(n7371) );
  INV_X1 U6552 ( .A(\Mcontrol/Nextpc_decoding/N219 ), .ZN(n7594) );
  INV_X1 U6553 ( .A(\Mcontrol/Nextpc_decoding/N219 ), .ZN(n7668) );
  CLKBUF_X1 U6554 ( .A(n7871), .Z(I_ADDR_OUTBUS[21]) );
  NAND2_X1 U6555 ( .A1(\Mcontrol/Nextpc_decoding/Bta [21]), .A2(net58826), 
        .ZN(n7374) );
  NAND2_X1 U6556 ( .A1(jar_in[21]), .A2(n1561), .ZN(n7375) );
  AND3_X2 U6557 ( .A1(n7374), .A2(n7373), .A3(n7375), .ZN(n2681) );
  OR2_X4 U6558 ( .A1(n6956), .A2(n7376), .ZN(
        \Mcontrol/Operation_decoding32/N1975 ) );
  NAND2_X1 U6559 ( .A1(n7377), .A2(n7549), .ZN(n7376) );
  NOR2_X1 U6560 ( .A1(n7063), .A2(\Mcontrol/Operation_decoding32/N1990 ), .ZN(
        n7377) );
  CLKBUF_X1 U6561 ( .A(\Mcontrol/Operation_decoding32/N1987 ), .Z(n7378) );
  INV_X1 U6562 ( .A(n7229), .ZN(\Mcontrol/Operation_decoding32/N2060 ) );
  INV_X1 U6563 ( .A(n7465), .ZN(n7380) );
  NAND2_X1 U6564 ( .A1(branch_rega[0]), .A2(n7380), .ZN(n7381) );
  INV_X1 U6565 ( .A(n7662), .ZN(n7663) );
  INV_X2 U6566 ( .A(rd_addr[1]), .ZN(n1221) );
  CLKBUF_X1 U6567 ( .A(\Mcontrol/Operation_decoding32/N2007 ), .Z(n7384) );
  INV_X2 U6568 ( .A(\Mpath/out_regB[16] ), .ZN(n7385) );
  INV_X1 U6569 ( .A(n7385), .ZN(n7386) );
  INV_X1 U6570 ( .A(n7385), .ZN(n7388) );
  INV_X1 U6571 ( .A(n7385), .ZN(n7387) );
  OR2_X2 U6572 ( .A1(n7521), .A2(n7123), .ZN(n7389) );
  NAND2_X1 U6573 ( .A1(n7390), .A2(n7401), .ZN(
        \Mcontrol/Operation_decoding32/N2017 ) );
  CLKBUF_X1 U6574 ( .A(\Mcontrol/Operation_decoding32/N1963 ), .Z(n7391) );
  INV_X2 U6575 ( .A(\Mpath/out_regB[14] ), .ZN(n7392) );
  INV_X1 U6576 ( .A(n7392), .ZN(n7393) );
  INV_X1 U6577 ( .A(n7392), .ZN(n7395) );
  NAND2_X1 U6578 ( .A1(n7390), .A2(n7396), .ZN(n7504) );
  NOR2_X1 U6579 ( .A1(n7569), .A2(n7052), .ZN(n7396) );
  INV_X1 U6580 ( .A(\Mcontrol/d_instr [27]), .ZN(
        \Mcontrol/Operation_decoding32/N1921 ) );
  NAND2_X1 U6581 ( .A1(n7174), .A2(n7378), .ZN(n6252) );
  AOI221_X1 U6582 ( .B1(n1436), .B2(n1437), .C1(n7226), .C2(n7598), .A(n7449), 
        .ZN(n1430) );
  NAND2_X1 U6583 ( .A1(net58533), .A2(n7400), .ZN(net57386) );
  INV_X1 U6584 ( .A(n7043), .ZN(n7401) );
  CLKBUF_X1 U6585 ( .A(net58543), .Z(net57379) );
  CLKBUF_X1 U6586 ( .A(n7389), .Z(n7402) );
  INV_X1 U6587 ( .A(n7043), .ZN(n7403) );
  INV_X1 U6588 ( .A(\Mcontrol/Operation_decoding32/N1921 ), .ZN(n7447) );
  AND2_X2 U6589 ( .A1(n7404), .A2(n7405), .ZN(n2594) );
  OR3_X1 U6590 ( .A1(net56846), .A2(n6168), .A3(n7035), .ZN(n7404) );
  NAND2_X1 U6591 ( .A1(n7035), .A2(n5521), .ZN(n7405) );
  INV_X1 U6592 ( .A(net57236), .ZN(net57368) );
  INV_X1 U6593 ( .A(net56922), .ZN(net57366) );
  OR2_X1 U6594 ( .A1(rd_addr[3]), .A2(n6967), .ZN(\regfile/N279 ) );
  OR2_X1 U6595 ( .A1(rd_addr[3]), .A2(\regfile/N358 ), .ZN(\regfile/N285 ) );
  OR2_X1 U6596 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N317 ) );
  OR2_X1 U6597 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N323 ) );
  OR2_X1 U6598 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N335 ) );
  OR2_X1 U6599 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N329 ) );
  OR2_X1 U6600 ( .A1(rd_addr[3]), .A2(n6967), .ZN(\regfile/N298 ) );
  OR2_X1 U6601 ( .A1(rd_addr[3]), .A2(n6967), .ZN(\regfile/N310 ) );
  OR2_X1 U6602 ( .A1(rd_addr[3]), .A2(n6967), .ZN(\regfile/N292 ) );
  OR2_X1 U6603 ( .A1(rd_addr[3]), .A2(n6967), .ZN(\regfile/N304 ) );
  OR2_X1 U6604 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N347 ) );
  OR2_X1 U6605 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N341 ) );
  OR2_X1 U6606 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N359 ) );
  OR2_X1 U6607 ( .A1(\regfile/N315 ), .A2(n6967), .ZN(\regfile/N353 ) );
  NOR2_X1 U6608 ( .A1(net56678), .A2(n7041), .ZN(n7409) );
  NOR3_X1 U6609 ( .A1(n7228), .A2(n7384), .A3(n7527), .ZN(n7410) );
  NAND2_X1 U6610 ( .A1(net58533), .A2(n7411), .ZN(
        \Mcontrol/Operation_decoding32/N1957 ) );
  NOR2_X1 U6611 ( .A1(n7052), .A2(\Mcontrol/Operation_decoding32/N1955 ), .ZN(
        n7411) );
  AND3_X4 U6612 ( .A1(n7413), .A2(net57346), .A3(n7412), .ZN(n298) );
  INV_X32 U6613 ( .A(net55892), .ZN(net57346) );
  INV_X32 U6614 ( .A(n1251), .ZN(n7412) );
  NOR2_X1 U6615 ( .A1(\regfile/N290 ), .A2(\regfile/N456 ), .ZN(n7413) );
  INV_X1 U6616 ( .A(net56846), .ZN(net57341) );
  INV_X2 U6617 ( .A(n5521), .ZN(net56846) );
  OR2_X2 U6618 ( .A1(n7566), .A2(n7414), .ZN(
        \Mcontrol/Operation_decoding32/N2036 ) );
  INV_X1 U6619 ( .A(n7534), .ZN(n7416) );
  AND3_X4 U6620 ( .A1(n7418), .A2(net57331), .A3(n7417), .ZN(n295) );
  NOR2_X1 U6621 ( .A1(\regfile/N290 ), .A2(\regfile/N444 ), .ZN(n7418) );
  OAI222_X1 U6622 ( .A1(n6044), .A2(n7255), .B1(n7176), .B2(n6050), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n6047), .ZN(n6334) );
  OAI222_X1 U6623 ( .A1(n6049), .A2(n7454), .B1(n7176), .B2(n5904), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n6051), .ZN(n6370) );
  OAI222_X1 U6624 ( .A1(n6046), .A2(n7454), .B1(n7176), .B2(n6051), .C1(
        \Mcontrol/Operation_decoding32/N1975 ), .C2(n6048), .ZN(n6346) );
  INV_X1 U6625 ( .A(n5521), .ZN(net57323) );
  NAND2_X1 U6626 ( .A1(n1478), .A2(n7040), .ZN(n7421) );
  NAND2_X1 U6627 ( .A1(n1478), .A2(n7550), .ZN(n6074) );
  NAND2_X1 U6628 ( .A1(n7568), .A2(\Mcontrol/Operation_decoding32/N2054 ), 
        .ZN(n7423) );
  NAND2_X1 U6629 ( .A1(n7092), .A2(n7389), .ZN(n7422) );
  INV_X1 U6630 ( .A(n7062), .ZN(n7425) );
  OR2_X2 U6631 ( .A1(n7426), .A2(net57313), .ZN(
        \Mcontrol/Operation_decoding32/N2084 ) );
  CLKBUF_X1 U6632 ( .A(n7038), .Z(n7427) );
  AND3_X4 U6633 ( .A1(n7429), .A2(net57297), .A3(n7428), .ZN(n290) );
  INV_X32 U6634 ( .A(net55892), .ZN(net57297) );
  NOR2_X1 U6635 ( .A1(\regfile/N290 ), .A2(\regfile/N444 ), .ZN(n7429) );
  INV_X1 U6636 ( .A(n7450), .ZN(n7430) );
  BUF_X4 U6637 ( .A(n7254), .Z(n7455) );
  CLKBUF_X1 U6638 ( .A(n7235), .Z(n7432) );
  INV_X1 U6639 ( .A(n7430), .ZN(n7433) );
  INV_X1 U6640 ( .A(n7433), .ZN(n7434) );
  INV_X1 U6641 ( .A(n7159), .ZN(n7436) );
  NAND2_X1 U6642 ( .A1(\Mcontrol/Operation_decoding32/N1951 ), .A2(
        \Mcontrol/Operation_decoding32/N1957 ), .ZN(n7437) );
  NOR2_X1 U6643 ( .A1(n1524), .A2(\Mcontrol/Operation_decoding32/N1982 ), .ZN(
        n7438) );
  AND3_X4 U6644 ( .A1(n7440), .A2(net57255), .A3(n7439), .ZN(n288) );
  NOR2_X1 U6645 ( .A1(\regfile/N290 ), .A2(\regfile/N438 ), .ZN(n7440) );
  CLKBUF_X1 U6646 ( .A(n6068), .Z(n7441) );
  INV_X32 U6647 ( .A(branch_rega[0]), .ZN(n7445) );
  INV_X1 U6648 ( .A(n7059), .ZN(n7446) );
  INV_X1 U6649 ( .A(net58594), .ZN(n6171) );
  NOR2_X1 U6650 ( .A1(n7401), .A2(\Mcontrol/Operation_decoding32/N2064 ), .ZN(
        n7448) );
  CLKBUF_X1 U6651 ( .A(n7093), .Z(n7449) );
  INV_X1 U6652 ( .A(n7061), .ZN(n7450) );
  INV_X1 U6653 ( .A(n6103), .ZN(n6173) );
  NAND2_X1 U6654 ( .A1(n1846), .A2(n7585), .ZN(n7451) );
  OR2_X2 U6655 ( .A1(\Mcontrol/Operation_decoding32/N1996 ), .A2(n7536), .ZN(
        \Mcontrol/Operation_decoding32/N2003 ) );
  NOR2_X1 U6656 ( .A1(n7126), .A2(\Mcontrol/Operation_decoding32/N2021 ), .ZN(
        n7453) );
  INV_X1 U6657 ( .A(n7532), .ZN(n7456) );
  OR2_X1 U6658 ( .A1(\Mpath/out_regA[21] ), .A2(\Mpath/out_regB[21] ), .ZN(
        \Mpath/the_alu/N136 ) );
  NAND2_X1 U6659 ( .A1(n7511), .A2(n7512), .ZN(n7457) );
  INV_X1 U6660 ( .A(n7691), .ZN(n7458) );
  OR2_X1 U6661 ( .A1(n7460), .A2(branch_rega[10]), .ZN(n7459) );
  INV_X1 U6662 ( .A(n7693), .ZN(n7460) );
  CLKBUF_X1 U6663 ( .A(n5628), .Z(n7461) );
  INV_X1 U6664 ( .A(n7230), .ZN(n7463) );
  NOR2_X1 U6665 ( .A1(branch_rega[8]), .A2(branch_rega[7]), .ZN(n7464) );
  OR2_X1 U6666 ( .A1(n7466), .A2(branch_rega[2]), .ZN(n7465) );
  INV_X1 U6667 ( .A(n7467), .ZN(n7466) );
  AND2_X2 U6668 ( .A1(n7618), .A2(n7617), .ZN(n6412) );
  OR3_X2 U6669 ( .A1(n6398), .A2(\Mcontrol/Nextpc_decoding/N171 ), .A3(n2877), 
        .ZN(net55921) );
  AND3_X1 U6670 ( .A1(n7382), .A2(rs1_addr[0]), .A3(n6417), .ZN(n5632) );
  AND2_X1 U6671 ( .A1(\Mcontrol/bp_logicB/N3 ), .A2(\Mcontrol/bp_logicB/N13 ), 
        .ZN(\Mcontrol/bp_logicB/N16 ) );
  NAND2_X1 U6672 ( .A1(n7563), .A2(n7564), .ZN(n7468) );
  OR2_X1 U6673 ( .A1(n7470), .A2(branch_rega[16]), .ZN(n7469) );
  INV_X1 U6674 ( .A(n7684), .ZN(n7470) );
  INV_X1 U6675 ( .A(branch_rega[27]), .ZN(n7471) );
  NAND2_X1 U6676 ( .A1(n7480), .A2(n7471), .ZN(n7472) );
  INV_X1 U6677 ( .A(n7489), .ZN(n7473) );
  INV_X1 U6678 ( .A(n7557), .ZN(n7475) );
  INV_X1 U6679 ( .A(\Mpath/the_alu/N44 ), .ZN(n7476) );
  AND2_X1 U6680 ( .A1(\Mcontrol/Nextpc_decoding/Bta [1]), .A2(n1560), .ZN(
        n7478) );
  INV_X1 U6681 ( .A(byp_controlB[2]), .ZN(\BYP_BRANCH_MUXB/N39 ) );
  INV_X4 U6682 ( .A(n5625), .ZN(n2324) );
  INV_X4 U6683 ( .A(n249), .ZN(n251) );
  INV_X1 U6684 ( .A(n7351), .ZN(\Mcontrol/Operation_decoding32/N1900 ) );
  NOR2_X1 U6685 ( .A1(n7173), .A2(rs1_addr[1]), .ZN(n6421) );
  NAND3_X1 U6686 ( .A1(rs1_addr[1]), .A2(n7173), .A3(n6429), .ZN(n5645) );
  OAI22_X2 U6687 ( .A1(n5518), .A2(n2594), .B1(n2630), .B2(n2595), .ZN(
        break_code[2]) );
  AOI211_X2 U6688 ( .C1(\regfile/reg_out[16][31] ), .C2(n2324), .A(n2432), .B(
        n2433), .ZN(n2425) );
  INV_X2 U6689 ( .A(n5653), .ZN(n7481) );
  INV_X4 U6690 ( .A(n7481), .ZN(n7484) );
  INV_X1 U6691 ( .A(n7194), .ZN(n7485) );
  INV_X2 U6692 ( .A(n7193), .ZN(n7486) );
  INV_X4 U6693 ( .A(n272), .ZN(n274) );
  INV_X4 U6694 ( .A(n268), .ZN(n269) );
  INV_X4 U6695 ( .A(n372), .ZN(n371) );
  NAND2_X4 U6696 ( .A1(n1655), .A2(n6547), .ZN(n372) );
  NAND2_X1 U6697 ( .A1(n6431), .A2(n6428), .ZN(n5651) );
  NAND3_X1 U6698 ( .A1(n6425), .A2(n6428), .A3(rs1_addr[1]), .ZN(n5639) );
  NAND2_X4 U6699 ( .A1(\Mcontrol/Operation_decoding32/N1873 ), .A2(n6042), 
        .ZN(rs2_addr[0]) );
  INV_X2 U6700 ( .A(n6034), .ZN(rs2_addr[3]) );
  OAI222_X4 U6701 ( .A1(n5576), .A2(n5523), .B1(n6987), .B2(n5525), .C1(n5578), 
        .C2(n5527), .ZN(branch_regb[22]) );
  OAI222_X4 U6702 ( .A1(n5615), .A2(n5523), .B1(n5616), .B2(n5525), .C1(n5617), 
        .C2(n5527), .ZN(branch_regb[10]) );
  AND2_X4 U6703 ( .A1(n6033), .A2(n6025), .ZN(n5774) );
  OAI22_X1 U6704 ( .A1(\Mcontrol/Nextpc_decoding/N26 ), .A2(n6399), .B1(n6400), 
        .B2(\Mcontrol/Nextpc_decoding/N325 ), .ZN(
        \Mcontrol/Nextpc_decoding/condition ) );
  AND3_X4 U6705 ( .A1(rs2_addr[3]), .A2(rs2_addr[4]), .A3(n6024), .ZN(n5768)
         );
  AND3_X1 U6706 ( .A1(n6397), .A2(n2878), .A3(\Mcontrol/st_logic/N103 ), .ZN(
        n7488) );
  INV_X1 U6707 ( .A(\Mcontrol/d_jump_type[3] ), .ZN(\Mcontrol/st_logic/N103 )
         );
  AND2_X2 U6708 ( .A1(n1685), .A2(n1686), .ZN(n6437) );
  AND3_X2 U6709 ( .A1(n7173), .A2(n7686), .A3(n6431), .ZN(n7641) );
  AND3_X4 U6710 ( .A1(n6034), .A2(n6026), .A3(n6024), .ZN(n5775) );
  NOR2_X2 U6711 ( .A1(\Mcontrol/Nextpc_decoding/N29 ), .A2(n6402), .ZN(n6403)
         );
  AND2_X4 U6712 ( .A1(n6021), .A2(n6024), .ZN(n5758) );
  OAI222_X4 U6713 ( .A1(n5561), .A2(n5523), .B1(n5562), .B2(n5525), .C1(n5563), 
        .C2(n5527), .ZN(branch_regb[27]) );
  INV_X2 U6714 ( .A(n5771), .ZN(n7490) );
  INV_X1 U6715 ( .A(n7490), .ZN(n7491) );
  INV_X1 U6716 ( .A(n7490), .ZN(n7493) );
  INV_X2 U6717 ( .A(n7490), .ZN(n7492) );
  NOR2_X1 U6718 ( .A1(branch_rega[22]), .A2(n7635), .ZN(n7494) );
  OR2_X1 U6719 ( .A1(n6074), .A2(n7397), .ZN(net57038) );
  OAI222_X4 U6720 ( .A1(n5618), .A2(n5621), .B1(n5514), .B2(n7486), .C1(n5620), 
        .C2(n5623), .ZN(branch_rega[0]) );
  NOR3_X4 U6721 ( .A1(\Mpath/N186 ), .A2(\Mpath/N190 ), .A3(\Mpath/N183 ), 
        .ZN(n6091) );
  INV_X1 U6722 ( .A(n7593), .ZN(n7495) );
  NAND2_X1 U6723 ( .A1(n7663), .A2(n7494), .ZN(n7496) );
  NAND2_X1 U6724 ( .A1(n371), .A2(\Mcontrol/f_currpc[5] ), .ZN(n7497) );
  NAND2_X1 U6725 ( .A1(n372), .A2(I_ADDR_OUTBUS[5]), .ZN(n7498) );
  INV_X1 U6726 ( .A(n373), .ZN(n7499) );
  AND3_X2 U6727 ( .A1(n7498), .A2(n7497), .A3(n7499), .ZN(n878) );
  INV_X2 U6728 ( .A(n5632), .ZN(n7500) );
  INV_X1 U6729 ( .A(n7500), .ZN(n7501) );
  INV_X2 U6730 ( .A(n7500), .ZN(n7503) );
  INV_X1 U6731 ( .A(n7604), .ZN(n7575) );
  INV_X2 U6732 ( .A(n5630), .ZN(n2335) );
  CLKBUF_X1 U6733 ( .A(net56996), .Z(net56982) );
  NAND2_X1 U6734 ( .A1(n7504), .A2(n7175), .ZN(n7584) );
  INV_X1 U6735 ( .A(net57730), .ZN(net56977) );
  CLKBUF_X1 U6736 ( .A(n6252), .Z(n7506) );
  NOR2_X1 U6737 ( .A1(\Mcontrol/Operation_decoding32/N1922 ), .A2(n7446), .ZN(
        n7507) );
  NAND2_X1 U6738 ( .A1(n7508), .A2(n7078), .ZN(
        \Mcontrol/Operation_decoding32/N2041 ) );
  NOR2_X1 U6739 ( .A1(n7540), .A2(\Mcontrol/d_instr [28]), .ZN(n7508) );
  INV_X1 U6740 ( .A(\Mcontrol/Operation_decoding32/N1982 ), .ZN(n7509) );
  CLKBUF_X1 U6741 ( .A(n7509), .Z(n7510) );
  NOR2_X1 U6742 ( .A1(branch_rega[26]), .A2(branch_rega[25]), .ZN(n7512) );
  AND2_X1 U6743 ( .A1(n6417), .A2(n6420), .ZN(n7514) );
  AND2_X4 U6744 ( .A1(n6417), .A2(n6420), .ZN(n5633) );
  INV_X1 U6745 ( .A(n7516), .ZN(n7517) );
  INV_X4 U6746 ( .A(n7516), .ZN(n7518) );
  OR2_X1 U6747 ( .A1(\Mcontrol/d_instr [26]), .A2(n7043), .ZN(n7521) );
  OR2_X1 U6748 ( .A1(n7256), .A2(n7526), .ZN(n7523) );
  INV_X1 U6749 ( .A(n6052), .ZN(n7705) );
  CLKBUF_X1 U6750 ( .A(n1846), .Z(n7525) );
  INV_X1 U6751 ( .A(n7524), .ZN(n7527) );
  INV_X1 U6752 ( .A(\Mcontrol/d_instr [28]), .ZN(n7528) );
  CLKBUF_X1 U6753 ( .A(n7507), .Z(n7529) );
  CLKBUF_X1 U6754 ( .A(n7384), .Z(n7530) );
  CLKBUF_X1 U6755 ( .A(n7527), .Z(n7531) );
  AND2_X4 U6756 ( .A1(n6017), .A2(n6018), .ZN(n5753) );
  CLKBUF_X1 U6757 ( .A(n7164), .Z(n7532) );
  INV_X1 U6758 ( .A(n7525), .ZN(n7533) );
  INV_X1 U6759 ( .A(n7533), .ZN(n7534) );
  NAND2_X1 U6760 ( .A1(n7537), .A2(n7538), .ZN(
        \Mcontrol/Operation_decoding32/N2029 ) );
  NOR2_X1 U6761 ( .A1(\Mcontrol/d_instr [28]), .A2(\Mcontrol/d_instr [27]), 
        .ZN(n7538) );
  NAND2_X1 U6762 ( .A1(n7143), .A2(n7160), .ZN(n7540) );
  NOR2_X1 U6763 ( .A1(\Mcontrol/d_instr [27]), .A2(
        \Mcontrol/Operation_decoding32/N1922 ), .ZN(n7542) );
  OR2_X1 U6764 ( .A1(n7513), .A2(\Mcontrol/Operation_decoding32/N1891 ), .ZN(
        \Mcontrol/Operation_decoding32/N1892 ) );
  OR2_X1 U6765 ( .A1(n6907), .A2(\Mcontrol/Operation_decoding32/N1890 ), .ZN(
        \Mcontrol/Operation_decoding32/N1891 ) );
  OAI21_X2 U6766 ( .B1(n6494), .B2(n6495), .A(N80), .ZN(\exc[DMEM_MISALIGN] )
         );
  INV_X1 U6767 ( .A(n7177), .ZN(n7545) );
  NAND2_X1 U6768 ( .A1(\Mcontrol/Operation_decoding32/N1939 ), .A2(
        \Mcontrol/Operation_decoding32/N1933 ), .ZN(n7547) );
  NAND2_X1 U6769 ( .A1(\Mcontrol/Operation_decoding32/N1939 ), .A2(
        \Mcontrol/Operation_decoding32/N1933 ), .ZN(n1845) );
  INV_X1 U6770 ( .A(n7647), .ZN(n7652) );
  NAND2_X1 U6771 ( .A1(n7535), .A2(n7379), .ZN(n7548) );
  NOR2_X1 U6772 ( .A1(n7043), .A2(\Mcontrol/d_instr [26]), .ZN(n7549) );
  AND2_X2 U6773 ( .A1(\Mcontrol/Operation_decoding32/N2066 ), .A2(n7570), .ZN(
        n7550) );
  NAND2_X1 U6774 ( .A1(n7383), .A2(n7452), .ZN(
        \Mcontrol/Operation_decoding32/N1933 ) );
  INV_X1 U6775 ( .A(n7226), .ZN(n6065) );
  OR2_X1 U6776 ( .A1(net58533), .A2(\Mcontrol/Operation_decoding32/N2029 ), 
        .ZN(n7552) );
  INV_X1 U6777 ( .A(n7698), .ZN(n7553) );
  NOR2_X1 U6778 ( .A1(n7574), .A2(n7553), .ZN(n7555) );
  NAND2_X1 U6779 ( .A1(n7654), .A2(n7655), .ZN(n7558) );
  NAND2_X1 U6780 ( .A1(net56316), .A2(n7559), .ZN(n7565) );
  INV_X1 U6781 ( .A(n7558), .ZN(n7559) );
  NAND2_X1 U6782 ( .A1(\Mcontrol/f_currpc[22] ), .A2(n371), .ZN(n7560) );
  INV_X1 U6783 ( .A(n373), .ZN(n7561) );
  NAND2_X4 U6784 ( .A1(\Mcontrol/Operation_decoding32/N1873 ), .A2(n6039), 
        .ZN(rs2_addr[2]) );
  OAI222_X4 U6785 ( .A1(n5623), .A2(n5545), .B1(n7487), .B2(n2614), .C1(n5621), 
        .C2(n5543), .ZN(branch_rega[3]) );
  INV_X1 U6786 ( .A(n7643), .ZN(n7562) );
  NOR2_X2 U6787 ( .A1(n7579), .A2(n7562), .ZN(n7564) );
  INV_X2 U6788 ( .A(n6026), .ZN(rs2_addr[4]) );
  OR2_X4 U6789 ( .A1(\Mcontrol/Operation_decoding32/N1893 ), .A2(
        \Mcontrol/Operation_decoding32/N1899 ), .ZN(
        \Mcontrol/Operation_decoding32/N1873 ) );
  OAI222_X4 U6790 ( .A1(n5623), .A2(n5614), .B1(n7487), .B2(n2861), .C1(n5621), 
        .C2(n5612), .ZN(branch_rega[11]) );
  INV_X4 U6791 ( .A(n5770), .ZN(n1927) );
  CLKBUF_X1 U6792 ( .A(n7199), .Z(n7567) );
  INV_X1 U6793 ( .A(net58533), .ZN(net56765) );
  OR2_X1 U6794 ( .A1(n6891), .A2(\Mcontrol/Operation_decoding32/N2046 ), .ZN(
        \Mcontrol/Operation_decoding32/N2047 ) );
  OAI222_X4 U6795 ( .A1(n5623), .A2(n5536), .B1(n7486), .B2(n2561), .C1(n5621), 
        .C2(n5534), .ZN(branch_rega[6]) );
  INV_X2 U6796 ( .A(n6020), .ZN(rs2_addr[1]) );
  NOR2_X4 U6797 ( .A1(n6026), .A2(rs2_addr[3]), .ZN(n6021) );
  OR2_X1 U6798 ( .A1(n6891), .A2(\Mcontrol/Operation_decoding32/N2070 ), .ZN(
        \Mcontrol/Operation_decoding32/N2071 ) );
  INV_X1 U6799 ( .A(n6060), .ZN(n7571) );
  INV_X4 U6800 ( .A(branch_rega[9]), .ZN(n7689) );
  NOR2_X1 U6801 ( .A1(n7581), .A2(branch_rega[27]), .ZN(n7572) );
  NOR2_X1 U6802 ( .A1(branch_rega[28]), .A2(\Mcontrol/Nextpc_decoding/N253 ), 
        .ZN(n7573) );
  OAI222_X4 U6803 ( .A1(n5561), .A2(n5621), .B1(n5510), .B2(n7487), .C1(n5563), 
        .C2(n5623), .ZN(branch_rega[27]) );
  NAND2_X1 U6804 ( .A1(n2751), .A2(n7575), .ZN(n7574) );
  OR2_X1 U6805 ( .A1(n7305), .A2(\Mcontrol/Operation_decoding32/N1944 ), .ZN(
        n7576) );
  NAND2_X1 U6806 ( .A1(n2459), .A2(n2458), .ZN(break_code[1]) );
  INV_X1 U6807 ( .A(n7576), .ZN(n2497) );
  NOR2_X1 U6808 ( .A1(n7422), .A2(n7166), .ZN(n1478) );
  INV_X1 U6809 ( .A(branch_rega[18]), .ZN(n7578) );
  NAND2_X1 U6810 ( .A1(n7582), .A2(n7578), .ZN(n7579) );
  INV_X1 U6811 ( .A(n5883), .ZN(n7659) );
  OAI222_X4 U6812 ( .A1(n5623), .A2(n5584), .B1(n7487), .B2(n2700), .C1(n5621), 
        .C2(n5582), .ZN(branch_rega[20]) );
  INV_X1 U6813 ( .A(branch_rega[10]), .ZN(n7680) );
  OR2_X1 U6814 ( .A1(branch_rega[25]), .A2(branch_rega[26]), .ZN(n7581) );
  AND2_X2 U6815 ( .A1(n6421), .A2(n7687), .ZN(n6420) );
  AND2_X1 U6816 ( .A1(n7583), .A2(n7589), .ZN(n7582) );
  INV_X1 U6817 ( .A(branch_rega[19]), .ZN(n7583) );
  INV_X1 U6818 ( .A(n7588), .ZN(n7589) );
  INV_X1 U6819 ( .A(\Mcontrol/st_logic/N82 ), .ZN(\Mcontrol/st_logic/N83 ) );
  NOR4_X4 U6820 ( .A1(n2455), .A2(n2452), .A3(n7633), .A4(\Mpath/the_alu/N498 ), .ZN(n6499) );
  NAND2_X4 U6821 ( .A1(n359), .A2(\Scc_coproc/N551 ), .ZN(n357) );
  NOR2_X4 U6822 ( .A1(n1600), .A2(serve_exception), .ZN(n359) );
  CLKBUF_X1 U6823 ( .A(break_code[1]), .Z(n7586) );
  NAND2_X1 U6824 ( .A1(n7420), .A2(n7543), .ZN(n7587) );
  NAND2_X1 U6825 ( .A1(n7577), .A2(n7543), .ZN(net56668) );
  INV_X4 U6826 ( .A(n5634), .ZN(n2333) );
  NAND2_X1 U6827 ( .A1(n5642), .A2(\regfile/reg_out[29][31] ), .ZN(n7590) );
  NAND2_X1 U6828 ( .A1(n5643), .A2(\regfile/reg_out[28][31] ), .ZN(n7591) );
  AND2_X1 U6829 ( .A1(n7590), .A2(n7591), .ZN(n6427) );
  INV_X1 U6830 ( .A(branch_rega[17]), .ZN(n7643) );
  AND2_X4 U6831 ( .A1(n6413), .A2(n6414), .ZN(n7592) );
  NOR4_X2 U6832 ( .A1(n2415), .A2(n2416), .A3(n2417), .A4(n2418), .ZN(n2414)
         );
  NAND3_X1 U6833 ( .A1(n6414), .A2(rs1_addr[4]), .A3(n7328), .ZN(n5635) );
  NOR2_X1 U6834 ( .A1(n7547), .A2(n7451), .ZN(n6059) );
  INV_X1 U6835 ( .A(branch_rega[16]), .ZN(n7670) );
  NOR2_X4 U6836 ( .A1(n1915), .A2(\Mpath/the_shift/N107 ), .ZN(n1701) );
  AND3_X1 U6837 ( .A1(n7415), .A2(n7552), .A3(n7225), .ZN(n7598) );
  INV_X1 U6838 ( .A(n7177), .ZN(n7599) );
  OAI222_X4 U6839 ( .A1(n5623), .A2(n5605), .B1(n7486), .B2(n2810), .C1(n5621), 
        .C2(n5603), .ZN(branch_rega[14]) );
  INV_X4 U6840 ( .A(n5635), .ZN(n2337) );
  OR2_X1 U6841 ( .A1(branch_rega[12]), .A2(branch_rega[11]), .ZN(n7600) );
  OR2_X1 U6842 ( .A1(branch_rega[3]), .A2(branch_rega[2]), .ZN(n7601) );
  INV_X32 U6843 ( .A(n7601), .ZN(n7602) );
  AND2_X4 U6844 ( .A1(n6413), .A2(n7619), .ZN(n7603) );
  OR2_X1 U6845 ( .A1(n7605), .A2(branch_rega[16]), .ZN(n7604) );
  INV_X1 U6846 ( .A(n7650), .ZN(n7605) );
  AND2_X1 U6847 ( .A1(n6413), .A2(n7619), .ZN(n5627) );
  OR2_X1 U6848 ( .A1(rs1_addr[2]), .A2(\regfile/N260 ), .ZN(\regfile/N261 ) );
  NAND2_X1 U6849 ( .A1(n5649), .A2(\regfile/reg_out[5][31] ), .ZN(n7606) );
  NAND2_X1 U6850 ( .A1(n5650), .A2(\regfile/reg_out[4][31] ), .ZN(n7607) );
  AND2_X1 U6851 ( .A1(n7606), .A2(n7607), .ZN(n6432) );
  AND2_X1 U6852 ( .A1(n7686), .A2(n6422), .ZN(n7608) );
  AND2_X4 U6853 ( .A1(n6420), .A2(n7608), .ZN(n5650) );
  NAND2_X1 U6854 ( .A1(n7501), .A2(\regfile/reg_out[21][31] ), .ZN(n7609) );
  NAND2_X1 U6855 ( .A1(n7514), .A2(\regfile/reg_out[20][31] ), .ZN(n7610) );
  AND2_X1 U6856 ( .A1(n7610), .A2(n7609), .ZN(n6419) );
  BUF_X4 U6857 ( .A(n5633), .Z(n7612) );
  INV_X1 U6858 ( .A(n7613), .ZN(n7614) );
  INV_X1 U6859 ( .A(n7613), .ZN(n7616) );
  INV_X1 U6860 ( .A(n7613), .ZN(n7615) );
  NAND2_X1 U6861 ( .A1(n5627), .A2(\regfile/reg_out[19][31] ), .ZN(n7617) );
  NAND2_X1 U6862 ( .A1(n5628), .A2(\regfile/reg_out[18][31] ), .ZN(n7618) );
  AND2_X1 U6863 ( .A1(rs1_addr[0]), .A2(rs1_addr[1]), .ZN(n7619) );
  AND2_X1 U6864 ( .A1(n7351), .A2(n7623), .ZN(
        \Mcontrol/Operation_decoding32/N1894 ) );
  INV_X1 U6865 ( .A(n7592), .ZN(n7620) );
  INV_X1 U6866 ( .A(n7620), .ZN(n7621) );
  NAND2_X1 U6867 ( .A1(n7050), .A2(n7622), .ZN(
        \Mcontrol/Operation_decoding32/N1880 ) );
  AND2_X2 U6868 ( .A1(n7672), .A2(\Mcontrol/Nextpc_decoding/N307 ), .ZN(n6408)
         );
  AND3_X1 U6869 ( .A1(n7867), .A2(n7866), .A3(n7865), .ZN(n7681) );
  OAI22_X4 U6870 ( .A1(n2507), .A2(n2860), .B1(n6051), .B2(n2509), .ZN(
        break_code[11]) );
  INV_X32 U6871 ( .A(branch_rega[5]), .ZN(n7624) );
  INV_X1 U6872 ( .A(n7630), .ZN(n7625) );
  NAND2_X1 U6873 ( .A1(n7626), .A2(n7627), .ZN(\Mcontrol/Nextpc_decoding/N249 ) );
  NOR2_X1 U6874 ( .A1(n7657), .A2(n7625), .ZN(n7627) );
  NAND2_X1 U6875 ( .A1(n6201), .A2(n7424), .ZN(n7628) );
  NAND2_X1 U6876 ( .A1(\Mcontrol/d_instr [2]), .A2(n6173), .ZN(n7629) );
  AND2_X1 U6877 ( .A1(n1556), .A2(n7685), .ZN(n7630) );
  AND3_X4 U6878 ( .A1(n6420), .A2(n2896), .A3(rs1_addr[3]), .ZN(n2331) );
  INV_X2 U6879 ( .A(n1696), .ZN(n7632) );
  INV_X8 U6880 ( .A(n7632), .ZN(n7634) );
  OR2_X1 U6881 ( .A1(branch_rega[18]), .A2(n7637), .ZN(n7636) );
  INV_X1 U6882 ( .A(n7648), .ZN(n7637) );
  AND2_X1 U6883 ( .A1(\Mcontrol/Nextpc_decoding/N295 ), .A2(n7298), .ZN(n7638)
         );
  NOR2_X1 U6884 ( .A1(n6411), .A2(n7638), .ZN(n6410) );
  OR2_X1 U6885 ( .A1(n5646), .A2(n1354), .ZN(n7639) );
  OR2_X1 U6886 ( .A1(n5647), .A2(n1210), .ZN(n7640) );
  NAND3_X1 U6887 ( .A1(n7639), .A2(n7640), .A3(n2431), .ZN(n2427) );
  INV_X1 U6888 ( .A(\Mcontrol/Nextpc_decoding/N294 ), .ZN(
        \Mcontrol/Nextpc_decoding/N295 ) );
  NAND2_X1 U6889 ( .A1(n6499), .A2(\Mpath/the_alu/N492 ), .ZN(n1693) );
  INV_X4 U6890 ( .A(n5639), .ZN(n2338) );
  OAI222_X4 U6891 ( .A1(n5623), .A2(n5539), .B1(n7487), .B2(n2578), .C1(n5621), 
        .C2(n5537), .ZN(branch_rega[5]) );
  NAND3_X4 U6892 ( .A1(n2446), .A2(n2445), .A3(\Mpath/the_alu/N480 ), .ZN(
        n1841) );
  AOI221_X1 U6893 ( .B1(n1687), .B2(n1688), .C1(n1689), .C2(n1690), .A(n1691), 
        .ZN(n1686) );
  NOR2_X1 U6894 ( .A1(n7664), .A2(branch_rega[17]), .ZN(n7648) );
  BUF_X8 U6895 ( .A(\Mpath/out_regB[3] ), .Z(n7708) );
  INV_X1 U6896 ( .A(branch_rega[24]), .ZN(n7671) );
  AOI211_X4 U6897 ( .C1(n1673), .C2(n6077), .A(n1672), .B(net55898), .ZN(n1676) );
  OR2_X1 U6898 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N321 ) );
  OR2_X1 U6899 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N315 ) );
  OR2_X1 U6900 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N309 ) );
  OR2_X1 U6901 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N303 ) );
  OR2_X1 U6902 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N297 ) );
  OR2_X1 U6903 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N285 ) );
  OR2_X1 U6904 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/Nextpc_decoding/N291 ) );
  INV_X1 U6905 ( .A(\Mcontrol/st_logic/branch_uses_main_mem_result ), .ZN(
        \Mcontrol/st_logic/N25 ) );
  INV_X1 U6906 ( .A(\Mcontrol/st_logic/branch_uses_rega ), .ZN(
        \Mcontrol/st_logic/N51 ) );
  OR2_X1 U6907 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N60 ) );
  OR2_X1 U6908 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N67 ) );
  OR2_X1 U6909 ( .A1(\Mcontrol/st_logic/N103 ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N105 ) );
  OR2_X1 U6910 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N98 ) );
  OR2_X1 U6911 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N92 ) );
  OR2_X1 U6912 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N85 ) );
  OR2_X1 U6913 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N73 ) );
  OR2_X1 U6914 ( .A1(\Mcontrol/d_jump_type[3] ), .A2(net58101), .ZN(
        \Mcontrol/st_logic/N79 ) );
  NAND2_X1 U6915 ( .A1(n371), .A2(\Mcontrol/f_currpc[23] ), .ZN(n7654) );
  INV_X1 U6916 ( .A(n373), .ZN(n7655) );
  INV_X1 U6917 ( .A(net56319), .ZN(n5743) );
  NOR2_X1 U6918 ( .A1(n7544), .A2(n6068), .ZN(n1844) );
  INV_X1 U6919 ( .A(n7667), .ZN(n7656) );
  OR2_X1 U6920 ( .A1(branch_rega[4]), .A2(branch_rega[3]), .ZN(n7657) );
  INV_X1 U6921 ( .A(branch_rega[15]), .ZN(n7684) );
  OR2_X4 U6922 ( .A1(\Mcontrol/bp_logicA/memory_main ), .A2(
        \Mcontrol/bp_logicA/exec_main ), .ZN(byp_controlA[2]) );
  INV_X4 U6923 ( .A(n292), .ZN(n294) );
  INV_X1 U6924 ( .A(branch_rega[25]), .ZN(n7667) );
  INV_X1 U6925 ( .A(n7670), .ZN(n7664) );
  NAND2_X1 U6926 ( .A1(n5637), .A2(\regfile/reg_out[25][31] ), .ZN(n7665) );
  NAND2_X1 U6927 ( .A1(n5638), .A2(\regfile/reg_out[24][31] ), .ZN(n7666) );
  AND2_X2 U6928 ( .A1(n7665), .A2(n7666), .ZN(n6423) );
  OR2_X1 U6929 ( .A1(n7063), .A2(\Mcontrol/Operation_decoding32/N1889 ), .ZN(
        \Mcontrol/Operation_decoding32/N1890 ) );
  OR2_X1 U6930 ( .A1(n7054), .A2(n7455), .ZN(
        \Mcontrol/Operation_decoding32/N1984 ) );
  NOR2_X1 U6931 ( .A1(branch_rega[0]), .A2(\Mcontrol/Nextpc_decoding/N249 ), 
        .ZN(n7669) );
  INV_X4 U6932 ( .A(n7074), .ZN(n313) );
  INV_X4 U6933 ( .A(n308), .ZN(n310) );
  INV_X4 U6934 ( .A(n7112), .ZN(n307) );
  NOR2_X1 U6935 ( .A1(n7421), .A2(n7397), .ZN(n6096) );
  INV_X4 U6936 ( .A(n237), .ZN(n239) );
  INV_X4 U6937 ( .A(n7115), .ZN(n262) );
  INV_X4 U6938 ( .A(n255), .ZN(n257) );
  INV_X4 U6939 ( .A(n7119), .ZN(n287) );
  INV_X4 U6940 ( .A(n282), .ZN(n284) );
  INV_X4 U6941 ( .A(n7122), .ZN(n281) );
  NAND2_X2 U6942 ( .A1(n1221), .A2(n1222), .ZN(n1108) );
  INV_X4 U6943 ( .A(n270), .ZN(n271) );
  INV_X4 U6944 ( .A(n298), .ZN(n300) );
  INV_X4 U6945 ( .A(n295), .ZN(n297) );
  INV_X4 U6946 ( .A(n290), .ZN(n291) );
  OR2_X1 U6947 ( .A1(n7152), .A2(n7039), .ZN(
        \Mcontrol/Operation_decoding32/N1923 ) );
  NAND3_X2 U6948 ( .A1(n7328), .A2(rs1_addr[1]), .A3(n6433), .ZN(n5654) );
  INV_X4 U6949 ( .A(n288), .ZN(n289) );
  INV_X4 U6950 ( .A(n246), .ZN(n248) );
  INV_X1 U6951 ( .A(rs1_addr[4]), .ZN(n6422) );
  INV_X2 U6952 ( .A(n7686), .ZN(rs1_addr[3]) );
  OAI222_X1 U6953 ( .A1(n5549), .A2(n5621), .B1(n5507), .B2(n7485), .C1(n5551), 
        .C2(n5623), .ZN(branch_rega[30]) );
  OR2_X1 U6954 ( .A1(\Mpath/out_regA[6] ), .A2(\Mpath/out_regB[6] ), .ZN(
        \Mpath/the_alu/N151 ) );
  AND2_X1 U6955 ( .A1(\Mpath/out_regA[6] ), .A2(\Mpath/out_regB[6] ), .ZN(
        \Mpath/the_alu/N119 ) );
  AND2_X4 U6956 ( .A1(n6414), .A2(n6422), .ZN(n6431) );
  AND3_X4 U6957 ( .A1(rs1_addr[3]), .A2(rs1_addr[4]), .A3(n6420), .ZN(n5643)
         );
  INV_X4 U6958 ( .A(n5645), .ZN(n2323) );
  OR2_X1 U6959 ( .A1(\Mpath/out_regA[7] ), .A2(\Mpath/out_regB[7] ), .ZN(
        \Mpath/the_alu/N150 ) );
  AND2_X1 U6960 ( .A1(\Mpath/out_regA[7] ), .A2(\Mpath/out_regB[7] ), .ZN(
        \Mpath/the_alu/N118 ) );
  XNOR2_X1 U6961 ( .A(\Mcontrol/m_sampled_xrd[3] ), .B(rs1_addr[3]), .ZN(n7678) );
  XNOR2_X1 U6962 ( .A(\Mcontrol/m_sampled_xrd[4] ), .B(rs1_addr[4]), .ZN(n7679) );
  AND3_X1 U6963 ( .A1(n7681), .A2(n7682), .A3(n7683), .ZN(
        \Mcontrol/bp_logicA/N2 ) );
  XNOR2_X1 U6964 ( .A(\Mcontrol/x_rd[3] ), .B(rs1_addr[3]), .ZN(n7682) );
  XNOR2_X1 U6965 ( .A(\Mcontrol/x_rd[4] ), .B(rs1_addr[4]), .ZN(n7683) );
  OR2_X1 U6966 ( .A1(\Mpath/out_regA[5] ), .A2(\Mpath/out_regB[5] ), .ZN(
        \Mpath/the_alu/N152 ) );
  AND2_X1 U6967 ( .A1(\Mpath/out_regA[5] ), .A2(\Mpath/out_regB[5] ), .ZN(
        \Mpath/the_alu/N120 ) );
  AND2_X4 U6968 ( .A1(n6424), .A2(n6425), .ZN(n5637) );
  AND3_X1 U6969 ( .A1(rs1_addr[1]), .A2(rs1_addr[2]), .A3(n6429), .ZN(n7688)
         );
  OAI222_X4 U6970 ( .A1(n5623), .A2(n5554), .B1(n7487), .B2(n2632), .C1(n5621), 
        .C2(n5552), .ZN(branch_rega[2]) );
  INV_X1 U6971 ( .A(byp_controlA[2]), .ZN(\Mcontrol/st_logic/N55 ) );
  OAI222_X4 U6972 ( .A1(n5623), .A2(n5581), .B1(n7486), .B2(n2683), .C1(n5621), 
        .C2(n5579), .ZN(branch_rega[21]) );
  AND2_X4 U6973 ( .A1(n6426), .A2(n6416), .ZN(n6424) );
  AND3_X4 U6974 ( .A1(rs1_addr[4]), .A2(n7687), .A3(n6424), .ZN(n5638) );
  NOR4_X2 U6975 ( .A1(n2427), .A2(n2429), .A3(n2430), .A4(n2428), .ZN(n2426)
         );
  NAND3_X4 U6976 ( .A1(rs1_addr[1]), .A2(n6428), .A3(n6433), .ZN(n5652) );
  NAND3_X4 U6977 ( .A1(rs1_addr[2]), .A2(n7686), .A3(n6431), .ZN(n5647) );
  OR2_X4 U6978 ( .A1(n5892), .A2(n6434), .ZN(n7686) );
  OR2_X1 U6979 ( .A1(n7463), .A2(n7065), .ZN(
        \Mcontrol/Operation_decoding32/N1889 ) );
  OR2_X1 U6980 ( .A1(rs1_addr[1]), .A2(\regfile/N261 ), .ZN(\regfile/N262 ) );
  NAND2_X4 U6981 ( .A1(\Mcontrol/st_logic/N47 ), .A2(byp_controlA[2]), .ZN(
        n5621) );
  AND2_X1 U6982 ( .A1(\Mpath/out_regA[19] ), .A2(n7332), .ZN(
        \Mpath/the_alu/N106 ) );
  OR2_X1 U6983 ( .A1(\Mpath/out_regA[19] ), .A2(n7333), .ZN(
        \Mpath/the_alu/N138 ) );
  NAND3_X4 U6984 ( .A1(rs1_addr[0]), .A2(n6416), .A3(n6413), .ZN(n5624) );
  NAND2_X4 U6985 ( .A1(byp_controlA[0]), .A2(byp_controlA[2]), .ZN(n5623) );
  NAND2_X4 U6986 ( .A1(n6424), .A2(n6433), .ZN(n2327) );
  AND2_X1 U6987 ( .A1(\Mpath/out_regA[18] ), .A2(n7360), .ZN(
        \Mpath/the_alu/N107 ) );
  OR2_X1 U6988 ( .A1(\Mpath/out_regA[18] ), .A2(n7361), .ZN(
        \Mpath/the_alu/N139 ) );
  OR2_X1 U6989 ( .A1(branch_rega[23]), .A2(branch_rega[22]), .ZN(n7690) );
  OR2_X1 U6990 ( .A1(branch_rega[9]), .A2(branch_rega[8]), .ZN(n7692) );
  NAND2_X1 U6991 ( .A1(n7696), .A2(n7695), .ZN(\Mcontrol/Nextpc_decoding/N198 ) );
  INV_X32 U6992 ( .A(n7694), .ZN(n7695) );
  CLKBUF_X1 U6993 ( .A(n7880), .Z(I_ADDR_OUTBUS[11]) );
  AND2_X1 U6994 ( .A1(n6102), .A2(n6517), .ZN(n7700) );
  AND2_X1 U6995 ( .A1(jar_in[11]), .A2(n1561), .ZN(n7702) );
  NOR3_X2 U6996 ( .A1(n7700), .A2(n7701), .A3(n7702), .ZN(n2859) );
  OAI222_X4 U6997 ( .A1(n5623), .A2(n5590), .B1(n7487), .B2(n2720), .C1(n5621), 
        .C2(n5588), .ZN(branch_rega[19]) );
  OR2_X1 U6998 ( .A1(\Mpath/out_regA[16] ), .A2(n7388), .ZN(
        \Mpath/the_alu/N141 ) );
  AND2_X1 U6999 ( .A1(\Mpath/out_regA[16] ), .A2(n7387), .ZN(
        \Mpath/the_alu/N109 ) );
  NAND3_X4 U7000 ( .A1(n7687), .A2(n2896), .A3(n6424), .ZN(n2329) );
  AND2_X1 U7001 ( .A1(\Mpath/out_regA[13] ), .A2(n7106), .ZN(
        \Mpath/the_alu/N112 ) );
  OR2_X1 U7002 ( .A1(\Mpath/out_regA[13] ), .A2(n7106), .ZN(
        \Mpath/the_alu/N144 ) );
  AND2_X4 U7003 ( .A1(n7703), .A2(n7326), .ZN(rs1_addr[1]) );
  OAI222_X4 U7004 ( .A1(n5623), .A2(n5587), .B1(n7487), .B2(n2464), .C1(n5621), 
        .C2(n5585), .ZN(branch_rega[1]) );
  AND2_X1 U7005 ( .A1(\Mpath/out_regA[17] ), .A2(n7344), .ZN(
        \Mpath/the_alu/N108 ) );
  OR2_X1 U7006 ( .A1(\Mpath/out_regA[17] ), .A2(n7344), .ZN(
        \Mpath/the_alu/N140 ) );
  AND2_X1 U7007 ( .A1(\Mpath/out_regA[15] ), .A2(n7323), .ZN(
        \Mpath/the_alu/N110 ) );
  OR2_X1 U7008 ( .A1(\Mpath/out_regA[15] ), .A2(n7323), .ZN(
        \Mpath/the_alu/N142 ) );
  AND2_X1 U7009 ( .A1(\Mpath/out_regA[14] ), .A2(n7394), .ZN(
        \Mpath/the_alu/N111 ) );
  OR2_X1 U7010 ( .A1(\Mpath/out_regA[14] ), .A2(n7395), .ZN(
        \Mpath/the_alu/N143 ) );
  AND2_X1 U7011 ( .A1(\Mpath/out_regA[20] ), .A2(n7476), .ZN(
        \Mpath/the_alu/N105 ) );
  OR2_X1 U7012 ( .A1(\Mpath/out_regA[20] ), .A2(n7476), .ZN(
        \Mpath/the_alu/N137 ) );
  AND2_X1 U7013 ( .A1(n7182), .A2(\Mpath/out_regB[12] ), .ZN(
        \Mpath/the_alu/N113 ) );
  OR2_X1 U7014 ( .A1(n7182), .A2(\Mpath/out_regB[12] ), .ZN(
        \Mpath/the_alu/N145 ) );
  OR2_X1 U7015 ( .A1(\Mpath/out_regA[9] ), .A2(\Mpath/out_regB[9] ), .ZN(
        \Mpath/the_alu/N148 ) );
  AND2_X1 U7016 ( .A1(\Mpath/out_regA[9] ), .A2(\Mpath/out_regB[9] ), .ZN(
        \Mpath/the_alu/N116 ) );
  AND2_X1 U7017 ( .A1(\Mpath/out_regA[11] ), .A2(\Mpath/out_regB[11] ), .ZN(
        \Mpath/the_alu/N114 ) );
  OR2_X1 U7018 ( .A1(\Mpath/out_regA[11] ), .A2(\Mpath/out_regB[11] ), .ZN(
        \Mpath/the_alu/N146 ) );
  NAND3_X4 U7019 ( .A1(n6416), .A2(n7173), .A3(n6429), .ZN(n2328) );
  OR2_X1 U7020 ( .A1(rs1_addr[3]), .A2(rs1_addr[4]), .ZN(\regfile/N260 ) );
  AND2_X1 U7021 ( .A1(n7185), .A2(n7615), .ZN(\Mpath/the_alu/N117 ) );
  OR2_X1 U7022 ( .A1(n7185), .A2(n7616), .ZN(\Mpath/the_alu/N149 ) );
  AND2_X1 U7023 ( .A1(\Mpath/out_regA[10] ), .A2(n7192), .ZN(
        \Mpath/the_alu/N115 ) );
  OR2_X1 U7024 ( .A1(\Mpath/out_regA[10] ), .A2(n7192), .ZN(
        \Mpath/the_alu/N147 ) );
  NOR2_X4 U7025 ( .A1(n7634), .A2(n2456), .ZN(n1698) );
  INV_X1 U7026 ( .A(n7267), .ZN(\Mcontrol/Nextpc_decoding/N219 ) );
  INV_X1 U7027 ( .A(net55870), .ZN(net55822) );
  INV_X1 U7028 ( .A(net55868), .ZN(net55824) );
  INV_X1 U7029 ( .A(net55868), .ZN(net55826) );
  INV_X1 U7030 ( .A(net55868), .ZN(net55828) );
  INV_X1 U7031 ( .A(net55868), .ZN(net55830) );
  INV_X1 U7032 ( .A(net55868), .ZN(net55832) );
  INV_X1 U7033 ( .A(net55870), .ZN(net55834) );
  INV_X1 U7034 ( .A(net55868), .ZN(net55836) );
  INV_X1 U7035 ( .A(net55866), .ZN(net55838) );
  INV_X1 U7036 ( .A(net55866), .ZN(net55840) );
  INV_X1 U7037 ( .A(net55866), .ZN(net55842) );
  INV_X1 U7038 ( .A(net55866), .ZN(net55844) );
  INV_X1 U7039 ( .A(net55866), .ZN(net55846) );
  INV_X1 U7040 ( .A(net55866), .ZN(net55848) );
  INV_X1 U7041 ( .A(net55866), .ZN(net55850) );
  INV_X1 U7042 ( .A(net55864), .ZN(net55852) );
  INV_X1 U7043 ( .A(net55868), .ZN(net55854) );
  INV_X1 U7044 ( .A(net55864), .ZN(net55856) );
  INV_X1 U7045 ( .A(net55864), .ZN(net55858) );
  INV_X1 U7046 ( .A(net55864), .ZN(net55860) );
  INV_X1 U7047 ( .A(net55864), .ZN(net55862) );
  CLKBUF_X3 U7048 ( .A(n220), .Z(net55864) );
  CLKBUF_X3 U7049 ( .A(n220), .Z(net55866) );
  CLKBUF_X3 U7050 ( .A(n220), .Z(net55868) );
  CLKBUF_X3 U7051 ( .A(n220), .Z(net55870) );
  CLKBUF_X3 U7052 ( .A(n220), .Z(net55872) );
  CLKBUF_X3 U7053 ( .A(n220), .Z(net55874) );
  CLKBUF_X3 U7054 ( .A(n220), .Z(net55876) );
  CLKBUF_X3 U7055 ( .A(n220), .Z(net55878) );
  CLKBUF_X3 U7056 ( .A(n220), .Z(net55880) );
  CLKBUF_X3 U7057 ( .A(n220), .Z(net55882) );
  CLKBUF_X3 U7058 ( .A(n220), .Z(net55884) );
  CLKBUF_X3 U7059 ( .A(n220), .Z(net55886) );
  CLKBUF_X3 U7060 ( .A(n220), .Z(net55888) );
  CLKBUF_X3 U7061 ( .A(n220), .Z(net55890) );
  CLKBUF_X3 U7062 ( .A(n220), .Z(net55892) );
  CLKBUF_X3 U7063 ( .A(n220), .Z(net55894) );
  CLKBUF_X3 U7064 ( .A(n220), .Z(net55898) );
  CLKBUF_X3 U7065 ( .A(n220), .Z(net55900) );
  CLKBUF_X3 U7066 ( .A(n220), .Z(net55902) );
  CLKBUF_X3 U7067 ( .A(n220), .Z(net55904) );
  CLKBUF_X3 U7068 ( .A(n220), .Z(net55906) );
  CLKBUF_X3 U7069 ( .A(n220), .Z(net55908) );
  CLKBUF_X3 U7070 ( .A(n220), .Z(net55910) );
  CLKBUF_X3 U7071 ( .A(n220), .Z(net55912) );
  CLKBUF_X3 U7072 ( .A(n220), .Z(net55914) );
  CLKBUF_X3 U7073 ( .A(n220), .Z(net55916) );
  CLKBUF_X3 U7074 ( .A(n220), .Z(net55918) );
  CLKBUF_X3 U7075 ( .A(\Mpath/out_regB[4] ), .Z(n7706) );
  CLKBUF_X3 U7076 ( .A(\Mpath/out_regB[4] ), .Z(n7707) );
  CLKBUF_X1 U7077 ( .A(\Mpath/out_regB[2] ), .Z(n7710) );
  CLKBUF_X3 U7078 ( .A(\Mpath/out_regB[1] ), .Z(n7712) );
  CLKBUF_X3 U7079 ( .A(\Mpath/out_regB[1] ), .Z(n7713) );
  CLKBUF_X3 U7080 ( .A(\Mpath/out_regB[0] ), .Z(n7714) );
  CLKBUF_X3 U7081 ( .A(\Mpath/out_regB[0] ), .Z(n7715) );
  CLKBUF_X1 U7082 ( .A(n7844), .Z(n7716) );
  CLKBUF_X1 U7083 ( .A(n7844), .Z(n7717) );
  CLKBUF_X1 U7084 ( .A(n7843), .Z(n7718) );
  CLKBUF_X1 U7085 ( .A(n7843), .Z(n7719) );
  CLKBUF_X1 U7086 ( .A(n7843), .Z(n7720) );
  CLKBUF_X1 U7087 ( .A(n7843), .Z(n7721) );
  CLKBUF_X1 U7088 ( .A(n7843), .Z(n7722) );
  CLKBUF_X1 U7089 ( .A(n7843), .Z(n7723) );
  CLKBUF_X1 U7090 ( .A(n7842), .Z(n7724) );
  CLKBUF_X1 U7091 ( .A(n7842), .Z(n7725) );
  CLKBUF_X1 U7092 ( .A(n7842), .Z(n7726) );
  CLKBUF_X1 U7093 ( .A(n7842), .Z(n7727) );
  CLKBUF_X1 U7094 ( .A(n7842), .Z(n7728) );
  CLKBUF_X1 U7095 ( .A(n7842), .Z(n7729) );
  CLKBUF_X1 U7096 ( .A(n7841), .Z(n7730) );
  CLKBUF_X1 U7097 ( .A(n7841), .Z(n7731) );
  CLKBUF_X1 U7098 ( .A(n7841), .Z(n7732) );
  CLKBUF_X1 U7099 ( .A(n7841), .Z(n7733) );
  CLKBUF_X1 U7100 ( .A(n7841), .Z(n7734) );
  CLKBUF_X1 U7101 ( .A(n7841), .Z(n7735) );
  CLKBUF_X1 U7102 ( .A(n7840), .Z(n7736) );
  CLKBUF_X1 U7103 ( .A(n7840), .Z(n7737) );
  CLKBUF_X1 U7104 ( .A(n7840), .Z(n7738) );
  CLKBUF_X1 U7105 ( .A(n7840), .Z(n7739) );
  CLKBUF_X1 U7106 ( .A(n7840), .Z(n7740) );
  CLKBUF_X1 U7107 ( .A(n7840), .Z(n7741) );
  CLKBUF_X1 U7108 ( .A(n7839), .Z(n7742) );
  CLKBUF_X1 U7109 ( .A(n7839), .Z(n7743) );
  CLKBUF_X1 U7110 ( .A(n7839), .Z(n7744) );
  CLKBUF_X1 U7111 ( .A(n7839), .Z(n7745) );
  CLKBUF_X1 U7112 ( .A(n7839), .Z(n7746) );
  CLKBUF_X1 U7113 ( .A(n7839), .Z(n7747) );
  CLKBUF_X1 U7114 ( .A(n7838), .Z(n7748) );
  CLKBUF_X1 U7115 ( .A(n7838), .Z(n7749) );
  CLKBUF_X1 U7116 ( .A(n7838), .Z(n7750) );
  CLKBUF_X1 U7117 ( .A(n7838), .Z(n7751) );
  CLKBUF_X1 U7118 ( .A(n7838), .Z(n7752) );
  CLKBUF_X1 U7119 ( .A(n7838), .Z(n7753) );
  CLKBUF_X1 U7120 ( .A(n7837), .Z(n7754) );
  CLKBUF_X1 U7121 ( .A(n7837), .Z(n7755) );
  CLKBUF_X1 U7122 ( .A(n7837), .Z(n7756) );
  CLKBUF_X1 U7123 ( .A(n7837), .Z(n7757) );
  CLKBUF_X1 U7124 ( .A(n7837), .Z(n7758) );
  CLKBUF_X1 U7125 ( .A(n7837), .Z(n7759) );
  CLKBUF_X1 U7126 ( .A(n7836), .Z(n7760) );
  CLKBUF_X1 U7127 ( .A(n7836), .Z(n7761) );
  CLKBUF_X1 U7128 ( .A(n7836), .Z(n7762) );
  CLKBUF_X1 U7129 ( .A(n7836), .Z(n7763) );
  CLKBUF_X1 U7130 ( .A(n7836), .Z(n7764) );
  CLKBUF_X1 U7131 ( .A(n7836), .Z(n7765) );
  CLKBUF_X1 U7132 ( .A(n7835), .Z(n7766) );
  CLKBUF_X1 U7133 ( .A(n7835), .Z(n7767) );
  CLKBUF_X1 U7134 ( .A(n7835), .Z(n7768) );
  CLKBUF_X1 U7135 ( .A(n7835), .Z(n7769) );
  CLKBUF_X1 U7136 ( .A(n7835), .Z(n7770) );
  CLKBUF_X1 U7137 ( .A(n7835), .Z(n7771) );
  CLKBUF_X1 U7138 ( .A(n7834), .Z(n7772) );
  CLKBUF_X1 U7139 ( .A(n7834), .Z(n7773) );
  CLKBUF_X1 U7140 ( .A(n7834), .Z(n7774) );
  CLKBUF_X1 U7141 ( .A(n7834), .Z(n7775) );
  CLKBUF_X1 U7142 ( .A(n7834), .Z(n7776) );
  CLKBUF_X1 U7143 ( .A(n7834), .Z(n7777) );
  CLKBUF_X1 U7144 ( .A(n7833), .Z(n7778) );
  CLKBUF_X1 U7145 ( .A(n7833), .Z(n7779) );
  CLKBUF_X1 U7146 ( .A(n7833), .Z(n7780) );
  CLKBUF_X1 U7147 ( .A(n7833), .Z(n7781) );
  CLKBUF_X1 U7148 ( .A(n7833), .Z(n7782) );
  CLKBUF_X1 U7149 ( .A(n7833), .Z(n7783) );
  CLKBUF_X1 U7150 ( .A(n7832), .Z(n7784) );
  CLKBUF_X1 U7151 ( .A(n7832), .Z(n7785) );
  CLKBUF_X1 U7152 ( .A(n7832), .Z(n7786) );
  CLKBUF_X1 U7153 ( .A(n7832), .Z(n7787) );
  CLKBUF_X1 U7154 ( .A(n7832), .Z(n7788) );
  CLKBUF_X1 U7155 ( .A(n7832), .Z(n7789) );
  CLKBUF_X1 U7156 ( .A(n7831), .Z(n7790) );
  CLKBUF_X1 U7157 ( .A(n7831), .Z(n7791) );
  CLKBUF_X1 U7158 ( .A(n7831), .Z(n7792) );
  CLKBUF_X1 U7159 ( .A(n7831), .Z(n7793) );
  CLKBUF_X1 U7160 ( .A(n7831), .Z(n7794) );
  CLKBUF_X1 U7161 ( .A(n7831), .Z(n7795) );
  CLKBUF_X1 U7162 ( .A(n7830), .Z(n7796) );
  CLKBUF_X1 U7163 ( .A(n7830), .Z(n7797) );
  CLKBUF_X1 U7164 ( .A(n7830), .Z(n7798) );
  CLKBUF_X1 U7165 ( .A(n7830), .Z(n7799) );
  CLKBUF_X1 U7166 ( .A(n7830), .Z(n7800) );
  CLKBUF_X1 U7167 ( .A(n7830), .Z(n7801) );
  CLKBUF_X1 U7168 ( .A(n7829), .Z(n7802) );
  CLKBUF_X1 U7169 ( .A(n7829), .Z(n7803) );
  CLKBUF_X1 U7170 ( .A(n7829), .Z(n7804) );
  CLKBUF_X1 U7171 ( .A(n7829), .Z(n7805) );
  CLKBUF_X1 U7172 ( .A(n7829), .Z(n7806) );
  CLKBUF_X1 U7173 ( .A(n7829), .Z(n7807) );
  CLKBUF_X1 U7174 ( .A(n7828), .Z(n7808) );
  CLKBUF_X1 U7175 ( .A(n7828), .Z(n7809) );
  CLKBUF_X1 U7176 ( .A(n7828), .Z(n7810) );
  CLKBUF_X1 U7177 ( .A(n7828), .Z(n7811) );
  CLKBUF_X1 U7178 ( .A(n7828), .Z(n7812) );
  CLKBUF_X1 U7179 ( .A(n7828), .Z(n7813) );
  CLKBUF_X1 U7180 ( .A(n7827), .Z(n7814) );
  CLKBUF_X1 U7181 ( .A(n7827), .Z(n7815) );
  CLKBUF_X1 U7182 ( .A(n7827), .Z(n7816) );
  CLKBUF_X1 U7183 ( .A(n7827), .Z(n7817) );
  CLKBUF_X1 U7184 ( .A(n7827), .Z(n7818) );
  CLKBUF_X1 U7185 ( .A(n7827), .Z(n7819) );
  CLKBUF_X1 U7186 ( .A(n7826), .Z(n7820) );
  CLKBUF_X1 U7187 ( .A(n7826), .Z(n7821) );
  CLKBUF_X1 U7188 ( .A(n7826), .Z(n7822) );
  CLKBUF_X1 U7189 ( .A(n7826), .Z(n7823) );
  CLKBUF_X1 U7190 ( .A(n7826), .Z(n7824) );
  CLKBUF_X1 U7191 ( .A(n7826), .Z(n7825) );
  CLKBUF_X3 U7192 ( .A(n7851), .Z(n7826) );
  CLKBUF_X3 U7193 ( .A(n7850), .Z(n7827) );
  CLKBUF_X3 U7194 ( .A(n7850), .Z(n7828) );
  CLKBUF_X3 U7195 ( .A(n7850), .Z(n7829) );
  CLKBUF_X3 U7196 ( .A(n7849), .Z(n7830) );
  CLKBUF_X3 U7197 ( .A(n7849), .Z(n7831) );
  CLKBUF_X3 U7198 ( .A(n7849), .Z(n7832) );
  CLKBUF_X3 U7199 ( .A(n7848), .Z(n7833) );
  CLKBUF_X3 U7200 ( .A(n7848), .Z(n7834) );
  CLKBUF_X3 U7201 ( .A(n7848), .Z(n7835) );
  CLKBUF_X3 U7202 ( .A(n7847), .Z(n7836) );
  CLKBUF_X3 U7203 ( .A(n7847), .Z(n7837) );
  CLKBUF_X3 U7204 ( .A(n7847), .Z(n7838) );
  CLKBUF_X3 U7205 ( .A(n7846), .Z(n7839) );
  CLKBUF_X3 U7206 ( .A(n7846), .Z(n7840) );
  CLKBUF_X3 U7207 ( .A(n7846), .Z(n7841) );
  CLKBUF_X3 U7208 ( .A(n7845), .Z(n7842) );
  CLKBUF_X3 U7209 ( .A(n7845), .Z(n7843) );
  CLKBUF_X3 U7210 ( .A(n7852), .Z(n7845) );
  CLKBUF_X3 U7211 ( .A(n7852), .Z(n7846) );
  CLKBUF_X3 U7212 ( .A(n7852), .Z(n7847) );
  CLKBUF_X3 U7213 ( .A(n7852), .Z(n7848) );
  CLKBUF_X3 U7214 ( .A(n7852), .Z(n7849) );
  CLKBUF_X3 U7215 ( .A(n7852), .Z(n7850) );
  XNOR2_X1 U7216 ( .A(\Mcontrol/x_rd[0] ), .B(rs2_addr[0]), .ZN(n7855) );
  XNOR2_X1 U7217 ( .A(\Mcontrol/x_rd[2] ), .B(rs2_addr[2]), .ZN(n7854) );
  XNOR2_X1 U7218 ( .A(\Mcontrol/x_rd[1] ), .B(rs2_addr[1]), .ZN(n7853) );
  NAND3_X1 U7219 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(n7858) );
  XOR2_X1 U7220 ( .A(\Mcontrol/x_rd[3] ), .B(rs2_addr[3]), .Z(n7857) );
  XOR2_X1 U7221 ( .A(\Mcontrol/x_rd[4] ), .B(rs2_addr[4]), .Z(n7856) );
  NOR3_X1 U7222 ( .A1(n7858), .A2(n7857), .A3(n7856), .ZN(
        \Mcontrol/bp_logicB/N2 ) );
  XNOR2_X1 U7223 ( .A(\Mcontrol/m_sampled_xrd[0] ), .B(rs2_addr[0]), .ZN(n7861) );
  XNOR2_X1 U7224 ( .A(\Mcontrol/m_sampled_xrd[2] ), .B(rs2_addr[2]), .ZN(n7860) );
  XNOR2_X1 U7225 ( .A(\Mcontrol/m_sampled_xrd[1] ), .B(rs2_addr[1]), .ZN(n7859) );
  NAND3_X1 U7226 ( .A1(n7861), .A2(n7860), .A3(n7859), .ZN(n7864) );
  XOR2_X1 U7227 ( .A(\Mcontrol/m_sampled_xrd[3] ), .B(rs2_addr[3]), .Z(n7863)
         );
  XOR2_X1 U7228 ( .A(\Mcontrol/m_sampled_xrd[4] ), .B(rs2_addr[4]), .Z(n7862)
         );
  NOR3_X1 U7229 ( .A1(n7864), .A2(n7863), .A3(n7862), .ZN(
        \Mcontrol/bp_logicB/N3 ) );
  XNOR2_X1 U7230 ( .A(\Mcontrol/x_rd[0] ), .B(rs1_addr[0]), .ZN(n7867) );
  XNOR2_X1 U7231 ( .A(\Mcontrol/x_rd[2] ), .B(rs1_addr[2]), .ZN(n7866) );
  XNOR2_X1 U7232 ( .A(\Mcontrol/x_rd[1] ), .B(rs1_addr[1]), .ZN(n7865) );
  XNOR2_X1 U7233 ( .A(\Mcontrol/m_sampled_xrd[0] ), .B(rs1_addr[0]), .ZN(n7870) );
  XNOR2_X1 U7234 ( .A(\Mcontrol/m_sampled_xrd[2] ), .B(rs1_addr[2]), .ZN(n7869) );
  XNOR2_X1 U7235 ( .A(\Mcontrol/m_sampled_xrd[1] ), .B(rs1_addr[1]), .ZN(n7868) );
  OAI21_X1 U7236 ( .B1(n5720), .B2(n6305), .A(n6306), .ZN(n6303) );
  OAI21_X1 U7237 ( .B1(n5720), .B2(n6317), .A(n6318), .ZN(n6315) );
  OAI21_X1 U7238 ( .B1(n5720), .B2(n6291), .A(n6292), .ZN(n6289) );
  OAI21_X1 U7239 ( .B1(n5720), .B2(n6276), .A(n6277), .ZN(n6274) );
  OAI21_X1 U7240 ( .B1(n5720), .B2(n6247), .A(n6248), .ZN(n6245) );
  OAI21_X1 U7241 ( .B1(n5720), .B2(n6263), .A(n6264), .ZN(n6261) );
  OAI21_X1 U7242 ( .B1(n5720), .B2(n6235), .A(n6236), .ZN(n6233) );
  OAI21_X1 U7243 ( .B1(n5720), .B2(n6223), .A(n6224), .ZN(n6220) );
  OAI21_X1 U7244 ( .B1(n5720), .B2(n6341), .A(n6343), .ZN(n6340) );
  OAI21_X1 U7245 ( .B1(n5720), .B2(n6329), .A(n6331), .ZN(n6328) );
  OAI21_X1 U7246 ( .B1(n5720), .B2(n6365), .A(n6367), .ZN(n6364) );
  OAI21_X1 U7247 ( .B1(n5720), .B2(n6377), .A(n6379), .ZN(n6376) );
  OAI21_X1 U7248 ( .B1(n5720), .B2(n6139), .A(n6141), .ZN(n6138) );
  OAI21_X1 U7249 ( .B1(n5720), .B2(n6151), .A(n6153), .ZN(n6150) );
  OAI21_X1 U7250 ( .B1(n5720), .B2(n6114), .A(n6116), .ZN(n6113) );
  OAI21_X1 U7251 ( .B1(n5720), .B2(n6127), .A(n6129), .ZN(n6126) );
  OAI21_X1 U7252 ( .B1(n5720), .B2(n6353), .A(n6355), .ZN(n6352) );
  OAI21_X1 U7253 ( .B1(n5720), .B2(n6163), .A(n6165), .ZN(n6162) );
  OAI21_X1 U7254 ( .B1(n5720), .B2(n6194), .A(n6196), .ZN(n6193) );
  OAI21_X1 U7255 ( .B1(n5720), .B2(n6180), .A(n6182), .ZN(n6179) );
  OAI21_X1 U7256 ( .B1(n5720), .B2(n6209), .A(n6211), .ZN(n6208) );
  OAI21_X1 U7257 ( .B1(n5720), .B2(n6087), .A(n6090), .ZN(n6086) );
  NAND2_X1 U7258 ( .A1(\Mpath/out_jar[0] ), .A2(n5717), .ZN(n5716) );
  OAI21_X1 U7259 ( .B1(n5720), .B2(n6391), .A(n6393), .ZN(n6390) );
endmodule

