module up_island_DW_cmp_1 (
	A, 
	B, 
	TC, 
	GE_LT, 
	GE_GT_EQ, 
	GE_LT_GT_LE, 
	EQ_NE);
   input [31:0] A;
   input [31:0] B;
   input TC;
   input GE_LT;
   input GE_GT_EQ;
   output GE_LT_GT_LE;
   output EQ_NE;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;

   OAI21_X1 U1 (.ZN(GE_LT_GT_LE), 
	.B2(n6), 
	.B1(n1), 
	.A(n7));
   NAND2_X1 U2 (.ZN(n6), 
	.A2(n8), 
	.A1(n3));
   AOI21_X1 U3 (.ZN(n7), 
	.B2(n8), 
	.B1(n2), 
	.A(n9));
   NOR2_X1 U4 (.ZN(n8), 
	.A2(n10), 
	.A1(n5));
   OAI21_X1 U5 (.ZN(n9), 
	.B2(n10), 
	.B1(n4), 
	.A(n11));
   NAND2_X1 U6 (.ZN(n10), 
	.A2(n12), 
	.A1(n18));
   AOI21_X1 U7 (.ZN(n11), 
	.B2(n19), 
	.B1(n12), 
	.A(n13));
   NOR2_X1 U8 (.ZN(n12), 
	.A2(n14), 
	.A1(n16));
   OAI21_X1 U9 (.ZN(n13), 
	.B2(n17), 
	.B1(n14), 
	.A(n15));
   NOR2_X1 U10 (.ZN(n14), 
	.A2(B[31]), 
	.A1(n151));
   NAND2_X1 U11 (.ZN(n15), 
	.A2(B[31]), 
	.A1(n151));
   NOR2_X1 U12 (.ZN(n16), 
	.A2(B[30]), 
	.A1(n150));
   NAND2_X1 U13 (.ZN(n17), 
	.A2(B[30]), 
	.A1(n150));
   NOR2_X1 U14 (.ZN(n18), 
	.A2(n20), 
	.A1(n22));
   OAI21_X1 U15 (.ZN(n19), 
	.B2(n23), 
	.B1(n20), 
	.A(n21));
   NOR2_X1 U16 (.ZN(n20), 
	.A2(B[29]), 
	.A1(n149));
   NAND2_X1 U17 (.ZN(n21), 
	.A2(B[29]), 
	.A1(n149));
   NOR2_X1 U18 (.ZN(n22), 
	.A2(B[28]), 
	.A1(n148));
   NAND2_X1 U19 (.ZN(n23), 
	.A2(B[28]), 
	.A1(n148));
   NAND2_X1 U20 (.ZN(n5), 
	.A2(n24), 
	.A1(n30));
   AOI21_X1 U21 (.ZN(n4), 
	.B2(n31), 
	.B1(n24), 
	.A(n25));
   NOR2_X1 U22 (.ZN(n24), 
	.A2(n26), 
	.A1(n28));
   OAI21_X1 U23 (.ZN(n25), 
	.B2(n29), 
	.B1(n26), 
	.A(n27));
   NOR2_X1 U24 (.ZN(n26), 
	.A2(B[27]), 
	.A1(n147));
   NAND2_X1 U25 (.ZN(n27), 
	.A2(B[27]), 
	.A1(n147));
   NOR2_X1 U26 (.ZN(n28), 
	.A2(B[26]), 
	.A1(n146));
   NAND2_X1 U27 (.ZN(n29), 
	.A2(B[26]), 
	.A1(n146));
   NOR2_X1 U28 (.ZN(n30), 
	.A2(n32), 
	.A1(n34));
   OAI21_X1 U29 (.ZN(n31), 
	.B2(n35), 
	.B1(n32), 
	.A(n33));
   NOR2_X1 U30 (.ZN(n32), 
	.A2(B[25]), 
	.A1(n145));
   NAND2_X1 U31 (.ZN(n33), 
	.A2(B[25]), 
	.A1(n145));
   NOR2_X1 U32 (.ZN(n34), 
	.A2(B[24]), 
	.A1(n144));
   NAND2_X1 U33 (.ZN(n35), 
	.A2(B[24]), 
	.A1(n144));
   NOR2_X1 U34 (.ZN(n3), 
	.A2(n36), 
	.A1(n50));
   OAI21_X1 U35 (.ZN(n2), 
	.B2(n36), 
	.B1(n51), 
	.A(n37));
   NAND2_X1 U36 (.ZN(n36), 
	.A2(n38), 
	.A1(n44));
   AOI21_X1 U37 (.ZN(n37), 
	.B2(n45), 
	.B1(n38), 
	.A(n39));
   NOR2_X1 U38 (.ZN(n38), 
	.A2(n40), 
	.A1(n42));
   OAI21_X1 U39 (.ZN(n39), 
	.B2(n43), 
	.B1(n40), 
	.A(n41));
   NOR2_X1 U40 (.ZN(n40), 
	.A2(B[23]), 
	.A1(n143));
   NAND2_X1 U41 (.ZN(n41), 
	.A2(B[23]), 
	.A1(n143));
   NOR2_X1 U42 (.ZN(n42), 
	.A2(B[22]), 
	.A1(n142));
   NAND2_X1 U43 (.ZN(n43), 
	.A2(B[22]), 
	.A1(n142));
   NOR2_X1 U44 (.ZN(n44), 
	.A2(n46), 
	.A1(n48));
   OAI21_X1 U45 (.ZN(n45), 
	.B2(n49), 
	.B1(n46), 
	.A(n47));
   NOR2_X1 U46 (.ZN(n46), 
	.A2(B[21]), 
	.A1(n141));
   NAND2_X1 U47 (.ZN(n47), 
	.A2(B[21]), 
	.A1(n141));
   NOR2_X1 U48 (.ZN(n48), 
	.A2(B[20]), 
	.A1(n140));
   NAND2_X1 U49 (.ZN(n49), 
	.A2(B[20]), 
	.A1(n140));
   NAND2_X1 U50 (.ZN(n50), 
	.A2(n52), 
	.A1(n58));
   AOI21_X1 U51 (.ZN(n51), 
	.B2(n59), 
	.B1(n52), 
	.A(n53));
   NOR2_X1 U52 (.ZN(n52), 
	.A2(n54), 
	.A1(n56));
   OAI21_X1 U53 (.ZN(n53), 
	.B2(n57), 
	.B1(n54), 
	.A(n55));
   NOR2_X1 U54 (.ZN(n54), 
	.A2(B[19]), 
	.A1(n139));
   NAND2_X1 U55 (.ZN(n55), 
	.A2(B[19]), 
	.A1(n139));
   NOR2_X1 U56 (.ZN(n56), 
	.A2(B[18]), 
	.A1(n138));
   NAND2_X1 U57 (.ZN(n57), 
	.A2(B[18]), 
	.A1(n138));
   NOR2_X1 U58 (.ZN(n58), 
	.A2(n60), 
	.A1(n62));
   OAI21_X1 U59 (.ZN(n59), 
	.B2(n63), 
	.B1(n60), 
	.A(n61));
   NOR2_X1 U60 (.ZN(n60), 
	.A2(B[17]), 
	.A1(n137));
   NAND2_X1 U61 (.ZN(n61), 
	.A2(B[17]), 
	.A1(n137));
   NOR2_X1 U62 (.ZN(n62), 
	.A2(B[16]), 
	.A1(n136));
   NAND2_X1 U63 (.ZN(n63), 
	.A2(B[16]), 
	.A1(n136));
   AOI21_X1 U64 (.ZN(n1), 
	.B2(n64), 
	.B1(n94), 
	.A(n65));
   NOR2_X1 U65 (.ZN(n64), 
	.A2(n66), 
	.A1(n80));
   OAI21_X1 U66 (.ZN(n65), 
	.B2(n66), 
	.B1(n81), 
	.A(n67));
   NAND2_X1 U67 (.ZN(n66), 
	.A2(n68), 
	.A1(n74));
   AOI21_X1 U68 (.ZN(n67), 
	.B2(n75), 
	.B1(n68), 
	.A(n69));
   NOR2_X1 U69 (.ZN(n68), 
	.A2(n70), 
	.A1(n72));
   OAI21_X1 U70 (.ZN(n69), 
	.B2(n73), 
	.B1(n70), 
	.A(n71));
   NOR2_X1 U71 (.ZN(n70), 
	.A2(B[15]), 
	.A1(n135));
   NAND2_X1 U72 (.ZN(n71), 
	.A2(B[15]), 
	.A1(n135));
   NOR2_X1 U73 (.ZN(n72), 
	.A2(B[14]), 
	.A1(n134));
   NAND2_X1 U74 (.ZN(n73), 
	.A2(B[14]), 
	.A1(n134));
   NOR2_X1 U75 (.ZN(n74), 
	.A2(n76), 
	.A1(n78));
   OAI21_X1 U76 (.ZN(n75), 
	.B2(n79), 
	.B1(n76), 
	.A(n77));
   NOR2_X1 U77 (.ZN(n76), 
	.A2(B[13]), 
	.A1(n133));
   NAND2_X1 U78 (.ZN(n77), 
	.A2(B[13]), 
	.A1(n133));
   NOR2_X1 U79 (.ZN(n78), 
	.A2(B[12]), 
	.A1(n132));
   NAND2_X1 U80 (.ZN(n79), 
	.A2(B[12]), 
	.A1(n132));
   NAND2_X1 U81 (.ZN(n80), 
	.A2(n82), 
	.A1(n88));
   AOI21_X1 U82 (.ZN(n81), 
	.B2(n89), 
	.B1(n82), 
	.A(n83));
   NOR2_X1 U83 (.ZN(n82), 
	.A2(n84), 
	.A1(n86));
   OAI21_X1 U84 (.ZN(n83), 
	.B2(n87), 
	.B1(n84), 
	.A(n85));
   NOR2_X1 U85 (.ZN(n84), 
	.A2(B[11]), 
	.A1(n131));
   NAND2_X1 U86 (.ZN(n85), 
	.A2(B[11]), 
	.A1(n131));
   NOR2_X1 U87 (.ZN(n86), 
	.A2(B[10]), 
	.A1(n130));
   NAND2_X1 U88 (.ZN(n87), 
	.A2(B[10]), 
	.A1(n130));
   NOR2_X1 U89 (.ZN(n88), 
	.A2(n90), 
	.A1(n92));
   OAI21_X1 U90 (.ZN(n89), 
	.B2(n93), 
	.B1(n90), 
	.A(n91));
   NOR2_X1 U91 (.ZN(n90), 
	.A2(B[9]), 
	.A1(n129));
   NAND2_X1 U92 (.ZN(n91), 
	.A2(B[9]), 
	.A1(n129));
   NOR2_X1 U93 (.ZN(n92), 
	.A2(B[8]), 
	.A1(n128));
   NAND2_X1 U94 (.ZN(n93), 
	.A2(B[8]), 
	.A1(n128));
   OAI21_X1 U95 (.ZN(n94), 
	.B2(n95), 
	.B1(n109), 
	.A(n96));
   NAND2_X1 U96 (.ZN(n95), 
	.A2(n97), 
	.A1(n103));
   AOI21_X1 U97 (.ZN(n96), 
	.B2(n104), 
	.B1(n97), 
	.A(n98));
   NOR2_X1 U98 (.ZN(n97), 
	.A2(n99), 
	.A1(n101));
   OAI21_X1 U99 (.ZN(n98), 
	.B2(n102), 
	.B1(n99), 
	.A(n100));
   NOR2_X1 U100 (.ZN(n99), 
	.A2(B[7]), 
	.A1(n127));
   NAND2_X1 U101 (.ZN(n100), 
	.A2(B[7]), 
	.A1(n127));
   NOR2_X1 U102 (.ZN(n101), 
	.A2(B[6]), 
	.A1(n126));
   NAND2_X1 U103 (.ZN(n102), 
	.A2(B[6]), 
	.A1(n126));
   NOR2_X1 U104 (.ZN(n103), 
	.A2(n105), 
	.A1(n107));
   OAI21_X1 U105 (.ZN(n104), 
	.B2(n108), 
	.B1(n105), 
	.A(n106));
   NOR2_X1 U106 (.ZN(n105), 
	.A2(B[5]), 
	.A1(n125));
   NAND2_X1 U107 (.ZN(n106), 
	.A2(B[5]), 
	.A1(n125));
   NOR2_X1 U108 (.ZN(n107), 
	.A2(B[4]), 
	.A1(n124));
   NAND2_X1 U109 (.ZN(n108), 
	.A2(B[4]), 
	.A1(n124));
   AOI21_X1 U110 (.ZN(n109), 
	.B2(n116), 
	.B1(n110), 
	.A(n111));
   NOR2_X1 U111 (.ZN(n110), 
	.A2(n112), 
	.A1(n114));
   OAI21_X1 U112 (.ZN(n111), 
	.B2(n115), 
	.B1(n112), 
	.A(n113));
   NOR2_X1 U113 (.ZN(n112), 
	.A2(B[3]), 
	.A1(n123));
   NAND2_X1 U114 (.ZN(n113), 
	.A2(B[3]), 
	.A1(n123));
   NOR2_X1 U115 (.ZN(n114), 
	.A2(B[2]), 
	.A1(n122));
   NAND2_X1 U116 (.ZN(n115), 
	.A2(B[2]), 
	.A1(n122));
   OAI21_X1 U117 (.ZN(n116), 
	.B2(n119), 
	.B1(n117), 
	.A(n118));
   INV_X1 U121 (.ZN(n151), 
	.A(A[31]));
   INV_X1 U157 (.ZN(n138), 
	.A(A[18]));
   INV_X1 U158 (.ZN(n135), 
	.A(A[15]));
   INV_X1 U159 (.ZN(n139), 
	.A(A[19]));
   INV_X1 U160 (.ZN(n140), 
	.A(A[20]));
   INV_X1 U161 (.ZN(n141), 
	.A(A[21]));
   INV_X1 U162 (.ZN(n129), 
	.A(A[9]));
   INV_X1 U163 (.ZN(n130), 
	.A(A[10]));
   INV_X1 U164 (.ZN(n142), 
	.A(A[22]));
   INV_X1 U165 (.ZN(n143), 
	.A(A[23]));
   INV_X1 U166 (.ZN(n128), 
	.A(A[8]));
   INV_X1 U167 (.ZN(n136), 
	.A(A[16]));
   INV_X1 U168 (.ZN(n137), 
	.A(A[17]));
   INV_X1 U169 (.ZN(n148), 
	.A(A[28]));
   INV_X1 U170 (.ZN(n147), 
	.A(A[27]));
   INV_X1 U171 (.ZN(n145), 
	.A(A[25]));
   INV_X1 U172 (.ZN(n150), 
	.A(A[30]));
   INV_X1 U173 (.ZN(n127), 
	.A(A[7]));
   INV_X1 U174 (.ZN(n134), 
	.A(A[14]));
   INV_X1 U175 (.ZN(n133), 
	.A(A[13]));
   INV_X1 U176 (.ZN(n131), 
	.A(A[11]));
   INV_X1 U177 (.ZN(n132), 
	.A(A[12]));
   INV_X1 U178 (.ZN(n149), 
	.A(A[29]));
   INV_X1 U179 (.ZN(n125), 
	.A(A[5]));
   INV_X1 U180 (.ZN(n146), 
	.A(A[26]));
   INV_X1 U181 (.ZN(n144), 
	.A(A[24]));
   INV_X1 U182 (.ZN(n126), 
	.A(A[6]));
   INV_X1 U183 (.ZN(n124), 
	.A(A[4]));
   INV_X1 U184 (.ZN(n121), 
	.A(A[1]));
   INV_X1 U185 (.ZN(n123), 
	.A(A[3]));
   INV_X1 U186 (.ZN(n122), 
	.A(A[2]));
   NAND2_X1 U187 (.ZN(n118), 
	.A2(B[1]), 
	.A1(n121));
   NOR2_X1 U188 (.ZN(n117), 
	.A2(B[1]), 
	.A1(n121));
   NAND2_X1 U189 (.ZN(n119), 
	.A2(B[0]), 
	.A1(n120));
   INV_X1 U190 (.ZN(n120), 
	.A(A[0]));
endmodule

module up_island_DW_cmp_0 (
	A, 
	B, 
	TC, 
	GE_LT, 
	GE_GT_EQ, 
	GE_LT_GT_LE, 
	EQ_NE);
   input [31:0] A;
   input [31:0] B;
   input TC;
   input GE_LT;
   input GE_GT_EQ;
   output GE_LT_GT_LE;
   output EQ_NE;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;

   OAI21_X1 U1 (.ZN(GE_LT_GT_LE), 
	.B2(n6), 
	.B1(n1), 
	.A(n7));
   NAND2_X1 U2 (.ZN(n6), 
	.A2(n8), 
	.A1(n3));
   AOI21_X1 U3 (.ZN(n7), 
	.B2(n8), 
	.B1(n2), 
	.A(n9));
   NOR2_X1 U4 (.ZN(n8), 
	.A2(n10), 
	.A1(n5));
   OAI21_X1 U5 (.ZN(n9), 
	.B2(n10), 
	.B1(n4), 
	.A(n11));
   NAND2_X1 U6 (.ZN(n10), 
	.A2(n12), 
	.A1(n18));
   AOI21_X1 U7 (.ZN(n11), 
	.B2(n19), 
	.B1(n12), 
	.A(n13));
   NOR2_X1 U8 (.ZN(n12), 
	.A2(n14), 
	.A1(n16));
   OAI21_X1 U9 (.ZN(n13), 
	.B2(n17), 
	.B1(n14), 
	.A(n15));
   NOR2_X1 U10 (.ZN(n14), 
	.A2(A[31]), 
	.A1(n151));
   NAND2_X1 U11 (.ZN(n15), 
	.A2(A[31]), 
	.A1(n151));
   NOR2_X1 U12 (.ZN(n16), 
	.A2(B[30]), 
	.A1(n150));
   NAND2_X1 U13 (.ZN(n17), 
	.A2(B[30]), 
	.A1(n150));
   NOR2_X1 U14 (.ZN(n18), 
	.A2(n20), 
	.A1(n22));
   OAI21_X1 U15 (.ZN(n19), 
	.B2(n23), 
	.B1(n20), 
	.A(n21));
   NOR2_X1 U16 (.ZN(n20), 
	.A2(B[29]), 
	.A1(n149));
   NAND2_X1 U17 (.ZN(n21), 
	.A2(B[29]), 
	.A1(n149));
   NOR2_X1 U18 (.ZN(n22), 
	.A2(B[28]), 
	.A1(n148));
   NAND2_X1 U19 (.ZN(n23), 
	.A2(B[28]), 
	.A1(n148));
   NAND2_X1 U20 (.ZN(n5), 
	.A2(n24), 
	.A1(n30));
   AOI21_X1 U21 (.ZN(n4), 
	.B2(n31), 
	.B1(n24), 
	.A(n25));
   NOR2_X1 U22 (.ZN(n24), 
	.A2(n26), 
	.A1(n28));
   OAI21_X1 U23 (.ZN(n25), 
	.B2(n29), 
	.B1(n26), 
	.A(n27));
   NOR2_X1 U24 (.ZN(n26), 
	.A2(B[27]), 
	.A1(n147));
   NAND2_X1 U25 (.ZN(n27), 
	.A2(B[27]), 
	.A1(n147));
   NOR2_X1 U26 (.ZN(n28), 
	.A2(B[26]), 
	.A1(n146));
   NAND2_X1 U27 (.ZN(n29), 
	.A2(B[26]), 
	.A1(n146));
   NOR2_X1 U28 (.ZN(n30), 
	.A2(n32), 
	.A1(n34));
   OAI21_X1 U29 (.ZN(n31), 
	.B2(n35), 
	.B1(n32), 
	.A(n33));
   NOR2_X1 U30 (.ZN(n32), 
	.A2(B[25]), 
	.A1(n145));
   NAND2_X1 U31 (.ZN(n33), 
	.A2(B[25]), 
	.A1(n145));
   NOR2_X1 U32 (.ZN(n34), 
	.A2(B[24]), 
	.A1(n144));
   NAND2_X1 U33 (.ZN(n35), 
	.A2(B[24]), 
	.A1(n144));
   NOR2_X1 U34 (.ZN(n3), 
	.A2(n36), 
	.A1(n50));
   OAI21_X1 U35 (.ZN(n2), 
	.B2(n36), 
	.B1(n51), 
	.A(n37));
   NAND2_X1 U36 (.ZN(n36), 
	.A2(n38), 
	.A1(n44));
   AOI21_X1 U37 (.ZN(n37), 
	.B2(n45), 
	.B1(n38), 
	.A(n39));
   NOR2_X1 U38 (.ZN(n38), 
	.A2(n40), 
	.A1(n42));
   OAI21_X1 U39 (.ZN(n39), 
	.B2(n43), 
	.B1(n40), 
	.A(n41));
   NOR2_X1 U40 (.ZN(n40), 
	.A2(B[23]), 
	.A1(n143));
   NAND2_X1 U41 (.ZN(n41), 
	.A2(B[23]), 
	.A1(n143));
   NOR2_X1 U42 (.ZN(n42), 
	.A2(B[22]), 
	.A1(n142));
   NAND2_X1 U43 (.ZN(n43), 
	.A2(B[22]), 
	.A1(n142));
   NOR2_X1 U44 (.ZN(n44), 
	.A2(n46), 
	.A1(n48));
   OAI21_X1 U45 (.ZN(n45), 
	.B2(n49), 
	.B1(n46), 
	.A(n47));
   NOR2_X1 U46 (.ZN(n46), 
	.A2(B[21]), 
	.A1(n141));
   NAND2_X1 U47 (.ZN(n47), 
	.A2(B[21]), 
	.A1(n141));
   NOR2_X1 U48 (.ZN(n48), 
	.A2(B[20]), 
	.A1(n140));
   NAND2_X1 U49 (.ZN(n49), 
	.A2(B[20]), 
	.A1(n140));
   NAND2_X1 U50 (.ZN(n50), 
	.A2(n52), 
	.A1(n58));
   AOI21_X1 U51 (.ZN(n51), 
	.B2(n59), 
	.B1(n52), 
	.A(n53));
   NOR2_X1 U52 (.ZN(n52), 
	.A2(n54), 
	.A1(n56));
   OAI21_X1 U53 (.ZN(n53), 
	.B2(n57), 
	.B1(n54), 
	.A(n55));
   NOR2_X1 U54 (.ZN(n54), 
	.A2(B[19]), 
	.A1(n139));
   NAND2_X1 U55 (.ZN(n55), 
	.A2(B[19]), 
	.A1(n139));
   NOR2_X1 U56 (.ZN(n56), 
	.A2(B[18]), 
	.A1(n138));
   NAND2_X1 U57 (.ZN(n57), 
	.A2(B[18]), 
	.A1(n138));
   NOR2_X1 U58 (.ZN(n58), 
	.A2(n60), 
	.A1(n62));
   OAI21_X1 U59 (.ZN(n59), 
	.B2(n63), 
	.B1(n60), 
	.A(n61));
   NOR2_X1 U60 (.ZN(n60), 
	.A2(B[17]), 
	.A1(n137));
   NAND2_X1 U61 (.ZN(n61), 
	.A2(B[17]), 
	.A1(n137));
   NOR2_X1 U62 (.ZN(n62), 
	.A2(B[16]), 
	.A1(n136));
   NAND2_X1 U63 (.ZN(n63), 
	.A2(B[16]), 
	.A1(n136));
   AOI21_X1 U64 (.ZN(n1), 
	.B2(n64), 
	.B1(n94), 
	.A(n65));
   NOR2_X1 U65 (.ZN(n64), 
	.A2(n66), 
	.A1(n80));
   OAI21_X1 U66 (.ZN(n65), 
	.B2(n66), 
	.B1(n81), 
	.A(n67));
   NAND2_X1 U67 (.ZN(n66), 
	.A2(n68), 
	.A1(n74));
   AOI21_X1 U68 (.ZN(n67), 
	.B2(n75), 
	.B1(n68), 
	.A(n69));
   NOR2_X1 U69 (.ZN(n68), 
	.A2(n70), 
	.A1(n72));
   OAI21_X1 U70 (.ZN(n69), 
	.B2(n73), 
	.B1(n70), 
	.A(n71));
   NOR2_X1 U71 (.ZN(n70), 
	.A2(B[15]), 
	.A1(n135));
   NAND2_X1 U72 (.ZN(n71), 
	.A2(B[15]), 
	.A1(n135));
   NOR2_X1 U73 (.ZN(n72), 
	.A2(B[14]), 
	.A1(n134));
   NAND2_X1 U74 (.ZN(n73), 
	.A2(B[14]), 
	.A1(n134));
   NOR2_X1 U75 (.ZN(n74), 
	.A2(n76), 
	.A1(n78));
   OAI21_X1 U76 (.ZN(n75), 
	.B2(n79), 
	.B1(n76), 
	.A(n77));
   NOR2_X1 U77 (.ZN(n76), 
	.A2(B[13]), 
	.A1(n133));
   NAND2_X1 U78 (.ZN(n77), 
	.A2(B[13]), 
	.A1(n133));
   NOR2_X1 U79 (.ZN(n78), 
	.A2(B[12]), 
	.A1(n132));
   NAND2_X1 U80 (.ZN(n79), 
	.A2(B[12]), 
	.A1(n132));
   NAND2_X1 U81 (.ZN(n80), 
	.A2(n82), 
	.A1(n88));
   AOI21_X1 U82 (.ZN(n81), 
	.B2(n89), 
	.B1(n82), 
	.A(n83));
   NOR2_X1 U83 (.ZN(n82), 
	.A2(n84), 
	.A1(n86));
   OAI21_X1 U84 (.ZN(n83), 
	.B2(n87), 
	.B1(n84), 
	.A(n85));
   NOR2_X1 U85 (.ZN(n84), 
	.A2(B[11]), 
	.A1(n131));
   NAND2_X1 U86 (.ZN(n85), 
	.A2(B[11]), 
	.A1(n131));
   NOR2_X1 U87 (.ZN(n86), 
	.A2(B[10]), 
	.A1(n130));
   NAND2_X1 U88 (.ZN(n87), 
	.A2(B[10]), 
	.A1(n130));
   NOR2_X1 U89 (.ZN(n88), 
	.A2(n90), 
	.A1(n92));
   OAI21_X1 U90 (.ZN(n89), 
	.B2(n93), 
	.B1(n90), 
	.A(n91));
   NOR2_X1 U91 (.ZN(n90), 
	.A2(B[9]), 
	.A1(n129));
   NAND2_X1 U92 (.ZN(n91), 
	.A2(B[9]), 
	.A1(n129));
   NOR2_X1 U93 (.ZN(n92), 
	.A2(B[8]), 
	.A1(n128));
   NAND2_X1 U94 (.ZN(n93), 
	.A2(B[8]), 
	.A1(n128));
   OAI21_X1 U95 (.ZN(n94), 
	.B2(n95), 
	.B1(n109), 
	.A(n96));
   NAND2_X1 U96 (.ZN(n95), 
	.A2(n97), 
	.A1(n103));
   AOI21_X1 U97 (.ZN(n96), 
	.B2(n104), 
	.B1(n97), 
	.A(n98));
   NOR2_X1 U98 (.ZN(n97), 
	.A2(n99), 
	.A1(n101));
   OAI21_X1 U99 (.ZN(n98), 
	.B2(n102), 
	.B1(n99), 
	.A(n100));
   NOR2_X1 U100 (.ZN(n99), 
	.A2(B[7]), 
	.A1(n127));
   NAND2_X1 U101 (.ZN(n100), 
	.A2(B[7]), 
	.A1(n127));
   NOR2_X1 U102 (.ZN(n101), 
	.A2(B[6]), 
	.A1(n126));
   NAND2_X1 U103 (.ZN(n102), 
	.A2(B[6]), 
	.A1(n126));
   NOR2_X1 U104 (.ZN(n103), 
	.A2(n105), 
	.A1(n107));
   OAI21_X1 U105 (.ZN(n104), 
	.B2(n108), 
	.B1(n105), 
	.A(n106));
   NOR2_X1 U106 (.ZN(n105), 
	.A2(B[5]), 
	.A1(n125));
   NAND2_X1 U107 (.ZN(n106), 
	.A2(B[5]), 
	.A1(n125));
   NOR2_X1 U108 (.ZN(n107), 
	.A2(B[4]), 
	.A1(n124));
   NAND2_X1 U109 (.ZN(n108), 
	.A2(B[4]), 
	.A1(n124));
   AOI21_X1 U110 (.ZN(n109), 
	.B2(n116), 
	.B1(n110), 
	.A(n111));
   NOR2_X1 U111 (.ZN(n110), 
	.A2(n112), 
	.A1(n114));
   OAI21_X1 U112 (.ZN(n111), 
	.B2(n115), 
	.B1(n112), 
	.A(n113));
   NOR2_X1 U113 (.ZN(n112), 
	.A2(B[3]), 
	.A1(n123));
   NAND2_X1 U114 (.ZN(n113), 
	.A2(B[3]), 
	.A1(n123));
   NOR2_X1 U115 (.ZN(n114), 
	.A2(B[2]), 
	.A1(n122));
   NAND2_X1 U116 (.ZN(n115), 
	.A2(B[2]), 
	.A1(n122));
   OAI21_X1 U117 (.ZN(n116), 
	.B2(n119), 
	.B1(n117), 
	.A(n118));
   INV_X1 U152 (.ZN(n151), 
	.A(B[31]));
   INV_X1 U157 (.ZN(n138), 
	.A(A[18]));
   INV_X1 U158 (.ZN(n135), 
	.A(A[15]));
   INV_X1 U159 (.ZN(n139), 
	.A(A[19]));
   INV_X1 U160 (.ZN(n140), 
	.A(A[20]));
   INV_X1 U161 (.ZN(n141), 
	.A(A[21]));
   INV_X1 U162 (.ZN(n129), 
	.A(A[9]));
   INV_X1 U163 (.ZN(n130), 
	.A(A[10]));
   INV_X1 U164 (.ZN(n142), 
	.A(A[22]));
   INV_X1 U165 (.ZN(n143), 
	.A(A[23]));
   INV_X1 U166 (.ZN(n128), 
	.A(A[8]));
   INV_X1 U167 (.ZN(n136), 
	.A(A[16]));
   INV_X1 U168 (.ZN(n137), 
	.A(A[17]));
   INV_X1 U169 (.ZN(n148), 
	.A(A[28]));
   INV_X1 U170 (.ZN(n147), 
	.A(A[27]));
   INV_X1 U171 (.ZN(n145), 
	.A(A[25]));
   INV_X1 U172 (.ZN(n150), 
	.A(A[30]));
   INV_X1 U173 (.ZN(n127), 
	.A(A[7]));
   INV_X1 U174 (.ZN(n134), 
	.A(A[14]));
   INV_X1 U175 (.ZN(n133), 
	.A(A[13]));
   INV_X1 U176 (.ZN(n131), 
	.A(A[11]));
   INV_X1 U177 (.ZN(n132), 
	.A(A[12]));
   INV_X1 U178 (.ZN(n149), 
	.A(A[29]));
   INV_X1 U179 (.ZN(n125), 
	.A(A[5]));
   INV_X1 U180 (.ZN(n146), 
	.A(A[26]));
   INV_X1 U181 (.ZN(n144), 
	.A(A[24]));
   INV_X1 U182 (.ZN(n126), 
	.A(A[6]));
   INV_X1 U183 (.ZN(n124), 
	.A(A[4]));
   INV_X1 U184 (.ZN(n121), 
	.A(A[1]));
   INV_X1 U185 (.ZN(n123), 
	.A(A[3]));
   INV_X1 U186 (.ZN(n122), 
	.A(A[2]));
   NAND2_X1 U187 (.ZN(n118), 
	.A2(B[1]), 
	.A1(n121));
   NOR2_X1 U188 (.ZN(n117), 
	.A2(B[1]), 
	.A1(n121));
   NAND2_X1 U189 (.ZN(n119), 
	.A2(B[0]), 
	.A1(n120));
   INV_X1 U190 (.ZN(n120), 
	.A(A[0]));
endmodule

module up_island_DW_leftsh_1 (
	A, 
	SH, 
	B, 
	FE_OFN163_UUT_Mpath_out_regB_3_, 
	FE_OFN180_UUT_Mpath_out_regB_0_, 
	FE_OFN184_UUT_Mpath_out_regB_0_);
   input [31:0] A;
   input [4:0] SH;
   output [31:0] B;
   input FE_OFN163_UUT_Mpath_out_regB_3_;
   input FE_OFN180_UUT_Mpath_out_regB_0_;
   input FE_OFN184_UUT_Mpath_out_regB_0_;

   // Internal wires
   wire n377;
   wire n378;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n389;
   wire n390;
   wire n395;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;

   INV_X1 U173 (.ZN(n549), 
	.A(A[18]));
   NAND2_X1 U174 (.ZN(n555), 
	.A2(n378), 
	.A1(A[15]));
   INV_X1 U175 (.ZN(n542), 
	.A(A[19]));
   INV_X1 U176 (.ZN(n529), 
	.A(A[20]));
   INV_X1 U177 (.ZN(n522), 
	.A(A[21]));
   INV_X1 U178 (.ZN(n494), 
	.A(A[9]));
   NAND2_X1 U179 (.ZN(n595), 
	.A2(n377), 
	.A1(A[9]));
   INV_X1 U180 (.ZN(n486), 
	.A(A[10]));
   NAND2_X1 U181 (.ZN(n587), 
	.A2(n377), 
	.A1(A[10]));
   INV_X1 U182 (.ZN(n515), 
	.A(A[22]));
   INV_X1 U183 (.ZN(n508), 
	.A(A[23]));
   INV_X1 U184 (.ZN(n502), 
	.A(A[8]));
   NAND2_X1 U185 (.ZN(n583), 
	.A2(n377), 
	.A1(A[8]));
   INV_X1 U186 (.ZN(n563), 
	.A(A[16]));
   INV_X1 U187 (.ZN(n556), 
	.A(A[17]));
   INV_X1 U188 (.ZN(n469), 
	.A(A[28]));
   INV_X1 U189 (.ZN(n477), 
	.A(A[27]));
   INV_X1 U190 (.ZN(n493), 
	.A(A[25]));
   INV_X1 U191 (.ZN(n446), 
	.A(A[30]));
   INV_X1 U192 (.ZN(n509), 
	.A(A[7]));
   NAND2_X1 U193 (.ZN(n591), 
	.A2(n377), 
	.A1(A[7]));
   INV_X1 U194 (.ZN(n447), 
	.A(A[14]));
   NAND2_X1 U195 (.ZN(n562), 
	.A2(n378), 
	.A1(A[14]));
   INV_X1 U196 (.ZN(n461), 
	.A(A[13]));
   NAND2_X1 U197 (.ZN(n569), 
	.A2(n378), 
	.A1(A[13]));
   INV_X1 U198 (.ZN(n478), 
	.A(A[11]));
   NAND2_X1 U199 (.ZN(n579), 
	.A2(n377), 
	.A1(A[11]));
   INV_X1 U200 (.ZN(n470), 
	.A(A[12]));
   NAND2_X1 U201 (.ZN(n574), 
	.A2(n378), 
	.A1(A[12]));
   INV_X1 U202 (.ZN(n460), 
	.A(A[29]));
   INV_X1 U203 (.ZN(n523), 
	.A(A[5]));
   NAND2_X1 U204 (.ZN(n592), 
	.A2(n377), 
	.A1(A[5]));
   INV_X1 U205 (.ZN(n485), 
	.A(A[26]));
   INV_X1 U206 (.ZN(n501), 
	.A(A[24]));
   INV_X1 U207 (.ZN(n516), 
	.A(A[6]));
   NAND2_X1 U208 (.ZN(n584), 
	.A2(n377), 
	.A1(A[6]));
   INV_X1 U209 (.ZN(n530), 
	.A(A[4]));
   NAND2_X1 U210 (.ZN(n585), 
	.A2(n377), 
	.A1(A[4]));
   NAND2_X1 U211 (.ZN(n593), 
	.A2(n377), 
	.A1(A[3]));
   INV_X1 U212 (.ZN(n543), 
	.A(A[3]));
   INV_X1 U213 (.ZN(n550), 
	.A(A[2]));
   NAND2_X1 U214 (.ZN(n586), 
	.A2(n377), 
	.A1(A[2]));
   INV_X1 U215 (.ZN(n564), 
	.A(A[0]));
   NAND2_X1 U216 (.ZN(n601), 
	.A2(n377), 
	.A1(A[0]));
   NAND2_X1 U217 (.ZN(n594), 
	.A2(n377), 
	.A1(A[1]));
   INV_X1 U218 (.ZN(n557), 
	.A(A[1]));
   INV_X1 U219 (.ZN(n377), 
	.A(SH[4]));
   INV_X1 U220 (.ZN(n378), 
	.A(SH[4]));
   INV_X1 U223 (.ZN(n381), 
	.A(SH[3]));
   INV_X1 U224 (.ZN(n382), 
	.A(SH[3]));
   INV_X1 U225 (.ZN(n383), 
	.A(SH[3]));
   INV_X1 U226 (.ZN(n384), 
	.A(SH[3]));
   INV_X1 U231 (.ZN(n389), 
	.A(SH[2]));
   INV_X1 U232 (.ZN(n390), 
	.A(SH[2]));
   INV_X1 U237 (.ZN(n395), 
	.A(SH[1]));
   MUX2_X1 U241 (.Z(B[9]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n400), 
	.A(n399));
   MUX2_X1 U242 (.Z(B[8]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n401), 
	.A(n400));
   INV_X1 U243 (.ZN(n400), 
	.A(n402));
   MUX2_X1 U244 (.Z(n402), 
	.S(SH[2]), 
	.B(n404), 
	.A(n403));
   MUX2_X1 U245 (.Z(B[7]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n405), 
	.A(n401));
   INV_X1 U246 (.ZN(n401), 
	.A(n406));
   MUX2_X1 U247 (.Z(n406), 
	.S(SH[2]), 
	.B(n408), 
	.A(n407));
   MUX2_X1 U248 (.Z(B[6]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n409), 
	.A(n405));
   INV_X1 U249 (.ZN(n405), 
	.A(n410));
   MUX2_X1 U250 (.Z(n410), 
	.S(SH[2]), 
	.B(n412), 
	.A(n411));
   MUX2_X1 U251 (.Z(B[5]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n413), 
	.A(n409));
   INV_X1 U252 (.ZN(n409), 
	.A(n414));
   MUX2_X1 U253 (.Z(n414), 
	.S(SH[2]), 
	.B(n416), 
	.A(n415));
   MUX2_X1 U254 (.Z(B[4]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n417), 
	.A(n413));
   INV_X1 U255 (.ZN(n413), 
	.A(n418));
   MUX2_X1 U256 (.Z(n418), 
	.S(SH[2]), 
	.B(n419), 
	.A(n404));
   NAND2_X1 U257 (.ZN(n404), 
	.A2(n381), 
	.A1(n420));
   INV_X1 U258 (.ZN(n420), 
	.A(n421));
   MUX2_X1 U259 (.Z(B[3]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n422), 
	.A(n417));
   INV_X1 U260 (.ZN(n417), 
	.A(n423));
   NAND2_X1 U261 (.ZN(n423), 
	.A2(n389), 
	.A1(n424));
   INV_X1 U262 (.ZN(n424), 
	.A(n408));
   NAND2_X1 U263 (.ZN(n408), 
	.A2(n381), 
	.A1(n425));
   INV_X1 U264 (.ZN(n425), 
	.A(n426));
   MUX2_X1 U265 (.Z(B[31]), 
	.S(SH[0]), 
	.B(n428), 
	.A(n427));
   MUX2_X1 U266 (.Z(n427), 
	.S(SH[2]), 
	.B(n430), 
	.A(n429));
   INV_X1 U267 (.ZN(n430), 
	.A(n431));
   MUX2_X1 U268 (.Z(n429), 
	.S(SH[3]), 
	.B(n433), 
	.A(n432));
   INV_X1 U269 (.ZN(n433), 
	.A(n434));
   MUX2_X1 U270 (.Z(n432), 
	.S(SH[1]), 
	.B(n436), 
	.A(n435));
   INV_X1 U271 (.ZN(n436), 
	.A(n437));
   MUX2_X1 U272 (.Z(n435), 
	.S(SH[4]), 
	.B(A[15]), 
	.A(A[31]));
   MUX2_X1 U273 (.Z(B[30]), 
	.S(SH[0]), 
	.B(n438), 
	.A(n428));
   INV_X1 U274 (.ZN(n428), 
	.A(n439));
   MUX2_X1 U275 (.Z(n439), 
	.S(SH[2]), 
	.B(n441), 
	.A(n440));
   MUX2_X1 U276 (.Z(n440), 
	.S(SH[3]), 
	.B(n443), 
	.A(n442));
   MUX2_X1 U277 (.Z(n442), 
	.S(SH[1]), 
	.B(n445), 
	.A(n444));
   MUX2_X1 U278 (.Z(n444), 
	.S(SH[4]), 
	.B(n447), 
	.A(n446));
   MUX2_X1 U279 (.Z(B[2]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n448), 
	.A(n422));
   INV_X1 U280 (.ZN(n422), 
	.A(n449));
   NAND2_X1 U281 (.ZN(n449), 
	.A2(n389), 
	.A1(n450));
   INV_X1 U282 (.ZN(n450), 
	.A(n412));
   NAND2_X1 U283 (.ZN(n412), 
	.A2(n382), 
	.A1(n451));
   INV_X1 U284 (.ZN(n451), 
	.A(n452));
   MUX2_X1 U285 (.Z(B[29]), 
	.S(SH[0]), 
	.B(n453), 
	.A(n438));
   INV_X1 U286 (.ZN(n438), 
	.A(n454));
   MUX2_X1 U287 (.Z(n454), 
	.S(SH[2]), 
	.B(n456), 
	.A(n455));
   MUX2_X1 U288 (.Z(n455), 
	.S(SH[3]), 
	.B(n458), 
	.A(n457));
   MUX2_X1 U289 (.Z(n457), 
	.S(SH[1]), 
	.B(n459), 
	.A(n437));
   MUX2_X1 U290 (.Z(n437), 
	.S(SH[4]), 
	.B(n461), 
	.A(n460));
   MUX2_X1 U291 (.Z(B[28]), 
	.S(SH[0]), 
	.B(n462), 
	.A(n453));
   INV_X1 U292 (.ZN(n453), 
	.A(n463));
   MUX2_X1 U293 (.Z(n463), 
	.S(SH[2]), 
	.B(n465), 
	.A(n464));
   MUX2_X1 U294 (.Z(n464), 
	.S(SH[3]), 
	.B(n467), 
	.A(n466));
   MUX2_X1 U295 (.Z(n466), 
	.S(SH[1]), 
	.B(n468), 
	.A(n445));
   MUX2_X1 U296 (.Z(n445), 
	.S(SH[4]), 
	.B(n470), 
	.A(n469));
   MUX2_X1 U297 (.Z(B[27]), 
	.S(SH[0]), 
	.B(n471), 
	.A(n462));
   INV_X1 U298 (.ZN(n462), 
	.A(n472));
   MUX2_X1 U299 (.Z(n472), 
	.S(SH[2]), 
	.B(n473), 
	.A(n431));
   MUX2_X1 U300 (.Z(n431), 
	.S(SH[3]), 
	.B(n475), 
	.A(n474));
   MUX2_X1 U301 (.Z(n474), 
	.S(SH[1]), 
	.B(n476), 
	.A(n459));
   MUX2_X1 U302 (.Z(n459), 
	.S(SH[4]), 
	.B(n478), 
	.A(n477));
   MUX2_X1 U303 (.Z(B[26]), 
	.S(SH[0]), 
	.B(n479), 
	.A(n471));
   INV_X1 U304 (.ZN(n471), 
	.A(n480));
   MUX2_X1 U305 (.Z(n480), 
	.S(SH[2]), 
	.B(n481), 
	.A(n441));
   MUX2_X1 U306 (.Z(n441), 
	.S(SH[3]), 
	.B(n483), 
	.A(n482));
   MUX2_X1 U307 (.Z(n482), 
	.S(SH[1]), 
	.B(n484), 
	.A(n468));
   MUX2_X1 U308 (.Z(n468), 
	.S(SH[4]), 
	.B(n486), 
	.A(n485));
   MUX2_X1 U309 (.Z(B[25]), 
	.S(SH[0]), 
	.B(n487), 
	.A(n479));
   INV_X1 U310 (.ZN(n479), 
	.A(n488));
   MUX2_X1 U311 (.Z(n488), 
	.S(SH[2]), 
	.B(n489), 
	.A(n456));
   MUX2_X1 U312 (.Z(n456), 
	.S(SH[3]), 
	.B(n491), 
	.A(n490));
   MUX2_X1 U313 (.Z(n490), 
	.S(SH[1]), 
	.B(n492), 
	.A(n476));
   MUX2_X1 U314 (.Z(n476), 
	.S(SH[4]), 
	.B(n494), 
	.A(n493));
   MUX2_X1 U315 (.Z(B[24]), 
	.S(SH[0]), 
	.B(n495), 
	.A(n487));
   INV_X1 U316 (.ZN(n487), 
	.A(n496));
   MUX2_X1 U317 (.Z(n496), 
	.S(SH[2]), 
	.B(n497), 
	.A(n465));
   MUX2_X1 U318 (.Z(n465), 
	.S(SH[3]), 
	.B(n499), 
	.A(n498));
   MUX2_X1 U319 (.Z(n498), 
	.S(SH[1]), 
	.B(n500), 
	.A(n484));
   MUX2_X1 U320 (.Z(n484), 
	.S(SH[4]), 
	.B(n502), 
	.A(n501));
   MUX2_X1 U321 (.Z(B[23]), 
	.S(SH[0]), 
	.B(n503), 
	.A(n495));
   INV_X1 U322 (.ZN(n495), 
	.A(n504));
   MUX2_X1 U323 (.Z(n504), 
	.S(SH[2]), 
	.B(n505), 
	.A(n473));
   MUX2_X1 U324 (.Z(n473), 
	.S(SH[3]), 
	.B(n506), 
	.A(n434));
   MUX2_X1 U325 (.Z(n434), 
	.S(SH[1]), 
	.B(n507), 
	.A(n492));
   MUX2_X1 U326 (.Z(n492), 
	.S(SH[4]), 
	.B(n509), 
	.A(n508));
   MUX2_X1 U327 (.Z(B[22]), 
	.S(SH[0]), 
	.B(n510), 
	.A(n503));
   INV_X1 U328 (.ZN(n503), 
	.A(n511));
   MUX2_X1 U329 (.Z(n511), 
	.S(SH[2]), 
	.B(n512), 
	.A(n481));
   MUX2_X1 U330 (.Z(n481), 
	.S(SH[3]), 
	.B(n513), 
	.A(n443));
   MUX2_X1 U331 (.Z(n443), 
	.S(SH[1]), 
	.B(n514), 
	.A(n500));
   MUX2_X1 U332 (.Z(n500), 
	.S(SH[4]), 
	.B(n516), 
	.A(n515));
   MUX2_X1 U333 (.Z(B[21]), 
	.S(SH[0]), 
	.B(n517), 
	.A(n510));
   INV_X1 U334 (.ZN(n510), 
	.A(n518));
   MUX2_X1 U335 (.Z(n518), 
	.S(SH[2]), 
	.B(n519), 
	.A(n489));
   MUX2_X1 U336 (.Z(n489), 
	.S(SH[3]), 
	.B(n520), 
	.A(n458));
   MUX2_X1 U337 (.Z(n458), 
	.S(SH[1]), 
	.B(n521), 
	.A(n507));
   MUX2_X1 U338 (.Z(n507), 
	.S(SH[4]), 
	.B(n523), 
	.A(n522));
   MUX2_X1 U339 (.Z(B[20]), 
	.S(SH[0]), 
	.B(n524), 
	.A(n517));
   INV_X1 U340 (.ZN(n517), 
	.A(n525));
   MUX2_X1 U341 (.Z(n525), 
	.S(SH[2]), 
	.B(n526), 
	.A(n497));
   MUX2_X1 U342 (.Z(n497), 
	.S(SH[3]), 
	.B(n527), 
	.A(n467));
   MUX2_X1 U343 (.Z(n467), 
	.S(SH[1]), 
	.B(n528), 
	.A(n514));
   MUX2_X1 U344 (.Z(n514), 
	.S(SH[4]), 
	.B(n530), 
	.A(n529));
   MUX2_X1 U345 (.Z(B[1]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n531), 
	.A(n448));
   INV_X1 U346 (.ZN(n531), 
	.A(n532));
   INV_X1 U347 (.ZN(n448), 
	.A(n533));
   NAND2_X1 U348 (.ZN(n533), 
	.A2(n390), 
	.A1(n534));
   INV_X1 U349 (.ZN(n534), 
	.A(n416));
   NAND2_X1 U350 (.ZN(n416), 
	.A2(n382), 
	.A1(n535));
   INV_X1 U351 (.ZN(n535), 
	.A(n536));
   MUX2_X1 U352 (.Z(B[19]), 
	.S(SH[0]), 
	.B(n537), 
	.A(n524));
   INV_X1 U353 (.ZN(n524), 
	.A(n538));
   MUX2_X1 U354 (.Z(n538), 
	.S(SH[2]), 
	.B(n539), 
	.A(n505));
   MUX2_X1 U355 (.Z(n505), 
	.S(SH[3]), 
	.B(n540), 
	.A(n475));
   MUX2_X1 U356 (.Z(n475), 
	.S(SH[1]), 
	.B(n541), 
	.A(n521));
   MUX2_X1 U357 (.Z(n521), 
	.S(SH[4]), 
	.B(n543), 
	.A(n542));
   MUX2_X1 U358 (.Z(B[18]), 
	.S(SH[0]), 
	.B(n544), 
	.A(n537));
   INV_X1 U359 (.ZN(n537), 
	.A(n545));
   MUX2_X1 U360 (.Z(n545), 
	.S(SH[2]), 
	.B(n546), 
	.A(n512));
   MUX2_X1 U361 (.Z(n512), 
	.S(SH[3]), 
	.B(n547), 
	.A(n483));
   MUX2_X1 U362 (.Z(n483), 
	.S(SH[1]), 
	.B(n548), 
	.A(n528));
   MUX2_X1 U363 (.Z(n528), 
	.S(SH[4]), 
	.B(n550), 
	.A(n549));
   MUX2_X1 U364 (.Z(B[17]), 
	.S(SH[0]), 
	.B(n551), 
	.A(n544));
   INV_X1 U365 (.ZN(n544), 
	.A(n552));
   MUX2_X1 U366 (.Z(n552), 
	.S(SH[2]), 
	.B(n553), 
	.A(n519));
   MUX2_X1 U367 (.Z(n519), 
	.S(SH[3]), 
	.B(n554), 
	.A(n491));
   MUX2_X1 U368 (.Z(n491), 
	.S(SH[1]), 
	.B(n555), 
	.A(n541));
   MUX2_X1 U369 (.Z(n541), 
	.S(SH[4]), 
	.B(n557), 
	.A(n556));
   MUX2_X1 U370 (.Z(B[16]), 
	.S(SH[0]), 
	.B(n558), 
	.A(n551));
   INV_X1 U371 (.ZN(n551), 
	.A(n559));
   MUX2_X1 U372 (.Z(n559), 
	.S(SH[2]), 
	.B(n560), 
	.A(n526));
   MUX2_X1 U373 (.Z(n526), 
	.S(SH[3]), 
	.B(n561), 
	.A(n499));
   MUX2_X1 U374 (.Z(n499), 
	.S(SH[1]), 
	.B(n562), 
	.A(n548));
   MUX2_X1 U375 (.Z(n548), 
	.S(SH[4]), 
	.B(n564), 
	.A(n563));
   MUX2_X1 U376 (.Z(B[15]), 
	.S(SH[0]), 
	.B(n565), 
	.A(n558));
   INV_X1 U377 (.ZN(n558), 
	.A(n566));
   MUX2_X1 U378 (.Z(n566), 
	.S(SH[2]), 
	.B(n567), 
	.A(n539));
   MUX2_X1 U379 (.Z(n539), 
	.S(SH[3]), 
	.B(n568), 
	.A(n506));
   MUX2_X1 U380 (.Z(n506), 
	.S(SH[1]), 
	.B(n569), 
	.A(n555));
   MUX2_X1 U381 (.Z(B[14]), 
	.S(FE_OFN180_UUT_Mpath_out_regB_0_), 
	.B(n570), 
	.A(n565));
   INV_X1 U382 (.ZN(n565), 
	.A(n571));
   MUX2_X1 U383 (.Z(n571), 
	.S(SH[2]), 
	.B(n572), 
	.A(n546));
   MUX2_X1 U384 (.Z(n546), 
	.S(SH[3]), 
	.B(n573), 
	.A(n513));
   MUX2_X1 U385 (.Z(n513), 
	.S(SH[1]), 
	.B(n574), 
	.A(n562));
   MUX2_X1 U386 (.Z(B[13]), 
	.S(FE_OFN180_UUT_Mpath_out_regB_0_), 
	.B(n575), 
	.A(n570));
   INV_X1 U387 (.ZN(n570), 
	.A(n576));
   MUX2_X1 U388 (.Z(n576), 
	.S(SH[2]), 
	.B(n577), 
	.A(n553));
   MUX2_X1 U389 (.Z(n553), 
	.S(SH[3]), 
	.B(n578), 
	.A(n520));
   MUX2_X1 U390 (.Z(n520), 
	.S(SH[1]), 
	.B(n579), 
	.A(n569));
   MUX2_X1 U391 (.Z(B[12]), 
	.S(FE_OFN180_UUT_Mpath_out_regB_0_), 
	.B(n580), 
	.A(n575));
   INV_X1 U392 (.ZN(n575), 
	.A(n581));
   MUX2_X1 U393 (.Z(n581), 
	.S(SH[2]), 
	.B(n403), 
	.A(n560));
   MUX2_X1 U394 (.Z(n403), 
	.S(FE_OFN163_UUT_Mpath_out_regB_3_), 
	.B(n582), 
	.A(n561));
   MUX2_X1 U395 (.Z(n561), 
	.S(SH[1]), 
	.B(n584), 
	.A(n583));
   MUX2_X1 U396 (.Z(n560), 
	.S(SH[3]), 
	.B(n421), 
	.A(n527));
   MUX2_X1 U397 (.Z(n421), 
	.S(SH[1]), 
	.B(n586), 
	.A(n585));
   MUX2_X1 U398 (.Z(n527), 
	.S(SH[1]), 
	.B(n587), 
	.A(n574));
   MUX2_X1 U399 (.Z(B[11]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n588), 
	.A(n580));
   INV_X1 U400 (.ZN(n580), 
	.A(n589));
   MUX2_X1 U401 (.Z(n589), 
	.S(SH[2]), 
	.B(n407), 
	.A(n567));
   NAND2_X1 U402 (.ZN(n407), 
	.A2(n383), 
	.A1(n590));
   INV_X1 U403 (.ZN(n590), 
	.A(n568));
   MUX2_X1 U404 (.Z(n568), 
	.S(SH[1]), 
	.B(n592), 
	.A(n591));
   MUX2_X1 U405 (.Z(n567), 
	.S(SH[3]), 
	.B(n426), 
	.A(n540));
   MUX2_X1 U406 (.Z(n426), 
	.S(SH[1]), 
	.B(n594), 
	.A(n593));
   MUX2_X1 U407 (.Z(n540), 
	.S(SH[1]), 
	.B(n595), 
	.A(n579));
   MUX2_X1 U408 (.Z(B[10]), 
	.S(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.B(n399), 
	.A(n588));
   INV_X1 U409 (.ZN(n399), 
	.A(n596));
   MUX2_X1 U410 (.Z(n596), 
	.S(SH[2]), 
	.B(n415), 
	.A(n577));
   NAND2_X1 U411 (.ZN(n415), 
	.A2(n383), 
	.A1(n597));
   INV_X1 U412 (.ZN(n597), 
	.A(n578));
   MUX2_X1 U413 (.Z(n578), 
	.S(SH[1]), 
	.B(n593), 
	.A(n592));
   MUX2_X1 U414 (.Z(n577), 
	.S(SH[3]), 
	.B(n536), 
	.A(n554));
   NAND2_X1 U415 (.ZN(n536), 
	.A2(n395), 
	.A1(n598));
   INV_X1 U416 (.ZN(n598), 
	.A(n594));
   MUX2_X1 U417 (.Z(n554), 
	.S(SH[1]), 
	.B(n591), 
	.A(n595));
   INV_X1 U418 (.ZN(n588), 
	.A(n599));
   MUX2_X1 U419 (.Z(n599), 
	.S(SH[2]), 
	.B(n411), 
	.A(n572));
   NAND2_X1 U420 (.ZN(n411), 
	.A2(n384), 
	.A1(n600));
   INV_X1 U421 (.ZN(n600), 
	.A(n573));
   MUX2_X1 U422 (.Z(n573), 
	.S(SH[1]), 
	.B(n585), 
	.A(n584));
   MUX2_X1 U423 (.Z(n572), 
	.S(SH[3]), 
	.B(n452), 
	.A(n547));
   MUX2_X1 U424 (.Z(n452), 
	.S(SH[1]), 
	.B(n601), 
	.A(n586));
   MUX2_X1 U425 (.Z(n547), 
	.S(SH[1]), 
	.B(n583), 
	.A(n587));
   NOR2_X1 U426 (.ZN(B[0]), 
	.A2(n532), 
	.A1(FE_OFN184_UUT_Mpath_out_regB_0_));
   NAND2_X1 U427 (.ZN(n532), 
	.A2(n390), 
	.A1(n602));
   INV_X1 U428 (.ZN(n602), 
	.A(n419));
   NAND2_X1 U429 (.ZN(n419), 
	.A2(n384), 
	.A1(n603));
   INV_X1 U430 (.ZN(n603), 
	.A(n582));
   NAND2_X1 U431 (.ZN(n582), 
	.A2(n395), 
	.A1(n604));
   INV_X1 U432 (.ZN(n604), 
	.A(n601));
endmodule

module up_island_DW01_bsh_1 (
	A, 
	SH, 
	B, 
	FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_);
   input [31:0] A;
   input [4:0] SH;
   output [31:0] B;
   input FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_;

   // Internal wires
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;

   INV_X1 U163 (.ZN(n402), 
	.A(A[18]));
   INV_X1 U164 (.ZN(n343), 
	.A(A[15]));
   INV_X1 U165 (.ZN(n383), 
	.A(A[19]));
   INV_X1 U166 (.ZN(n397), 
	.A(A[20]));
   INV_X1 U167 (.ZN(n385), 
	.A(A[21]));
   INV_X1 U168 (.ZN(n391), 
	.A(A[9]));
   INV_X1 U169 (.ZN(n405), 
	.A(A[10]));
   INV_X1 U170 (.ZN(n399), 
	.A(A[22]));
   INV_X1 U171 (.ZN(n390), 
	.A(A[23]));
   INV_X1 U172 (.ZN(n403), 
	.A(A[8]));
   INV_X1 U173 (.ZN(n336), 
	.A(A[16]));
   INV_X1 U174 (.ZN(n388), 
	.A(A[17]));
   INV_X1 U175 (.ZN(n368), 
	.A(A[28]));
   INV_X1 U176 (.ZN(n378), 
	.A(A[27]));
   INV_X1 U177 (.ZN(n392), 
	.A(A[25]));
   INV_X1 U178 (.ZN(n351), 
	.A(A[30]));
   INV_X1 U179 (.ZN(n389), 
	.A(A[7]));
   INV_X1 U180 (.ZN(n350), 
	.A(A[14]));
   INV_X1 U181 (.ZN(n357), 
	.A(A[13]));
   INV_X1 U182 (.ZN(n377), 
	.A(A[11]));
   INV_X1 U183 (.ZN(n367), 
	.A(A[12]));
   INV_X1 U184 (.ZN(n358), 
	.A(A[29]));
   INV_X1 U185 (.ZN(n384), 
	.A(A[5]));
   INV_X1 U186 (.ZN(n406), 
	.A(A[26]));
   INV_X1 U187 (.ZN(n404), 
	.A(A[24]));
   INV_X1 U188 (.ZN(n398), 
	.A(A[6]));
   INV_X1 U189 (.ZN(n396), 
	.A(A[4]));
   INV_X1 U190 (.ZN(n382), 
	.A(A[3]));
   INV_X1 U191 (.ZN(n401), 
	.A(A[2]));
   INV_X1 U192 (.ZN(n337), 
	.A(A[0]));
   INV_X1 U193 (.ZN(n387), 
	.A(A[1]));
   MUX2_X1 U209 (.Z(B[9]), 
	.S(SH[0]), 
	.B(n218), 
	.A(n217));
   MUX2_X1 U210 (.Z(B[8]), 
	.S(SH[0]), 
	.B(n219), 
	.A(n218));
   INV_X1 U211 (.ZN(n218), 
	.A(n220));
   MUX2_X1 U212 (.Z(n220), 
	.S(SH[2]), 
	.B(n222), 
	.A(n221));
   MUX2_X1 U213 (.Z(B[7]), 
	.S(SH[0]), 
	.B(n223), 
	.A(n219));
   INV_X1 U214 (.ZN(n219), 
	.A(n224));
   MUX2_X1 U215 (.Z(n224), 
	.S(SH[2]), 
	.B(n226), 
	.A(n225));
   MUX2_X1 U216 (.Z(B[6]), 
	.S(SH[0]), 
	.B(n227), 
	.A(n223));
   INV_X1 U217 (.ZN(n223), 
	.A(n228));
   MUX2_X1 U218 (.Z(n228), 
	.S(SH[2]), 
	.B(n230), 
	.A(n229));
   MUX2_X1 U219 (.Z(B[5]), 
	.S(SH[0]), 
	.B(n231), 
	.A(n227));
   INV_X1 U220 (.ZN(n227), 
	.A(n232));
   MUX2_X1 U221 (.Z(n232), 
	.S(SH[2]), 
	.B(n234), 
	.A(n233));
   MUX2_X1 U222 (.Z(B[4]), 
	.S(SH[0]), 
	.B(n235), 
	.A(n231));
   INV_X1 U223 (.ZN(n231), 
	.A(n236));
   MUX2_X1 U224 (.Z(n236), 
	.S(SH[2]), 
	.B(n237), 
	.A(n222));
   MUX2_X1 U225 (.Z(n222), 
	.S(SH[3]), 
	.B(n239), 
	.A(n238));
   MUX2_X1 U226 (.Z(B[3]), 
	.S(SH[0]), 
	.B(n240), 
	.A(n235));
   INV_X1 U227 (.ZN(n235), 
	.A(n241));
   MUX2_X1 U228 (.Z(n241), 
	.S(SH[2]), 
	.B(n242), 
	.A(n226));
   MUX2_X1 U229 (.Z(n226), 
	.S(SH[3]), 
	.B(n244), 
	.A(n243));
   MUX2_X1 U230 (.Z(B[31]), 
	.S(SH[0]), 
	.B(n246), 
	.A(n245));
   MUX2_X1 U231 (.Z(B[30]), 
	.S(SH[0]), 
	.B(n247), 
	.A(n246));
   INV_X1 U232 (.ZN(n246), 
	.A(n248));
   MUX2_X1 U233 (.Z(n248), 
	.S(SH[2]), 
	.B(n250), 
	.A(n249));
   MUX2_X1 U234 (.Z(B[2]), 
	.S(SH[0]), 
	.B(n251), 
	.A(n240));
   INV_X1 U235 (.ZN(n240), 
	.A(n252));
   MUX2_X1 U236 (.Z(n252), 
	.S(SH[2]), 
	.B(n249), 
	.A(n230));
   MUX2_X1 U237 (.Z(n249), 
	.S(SH[3]), 
	.B(n254), 
	.A(n253));
   MUX2_X1 U238 (.Z(n230), 
	.S(SH[3]), 
	.B(n256), 
	.A(n255));
   MUX2_X1 U239 (.Z(B[29]), 
	.S(SH[0]), 
	.B(n257), 
	.A(n247));
   INV_X1 U240 (.ZN(n247), 
	.A(n258));
   MUX2_X1 U241 (.Z(n258), 
	.S(SH[2]), 
	.B(n260), 
	.A(n259));
   MUX2_X1 U242 (.Z(B[28]), 
	.S(SH[0]), 
	.B(n261), 
	.A(n257));
   INV_X1 U243 (.ZN(n257), 
	.A(n262));
   MUX2_X1 U244 (.Z(n262), 
	.S(SH[2]), 
	.B(n264), 
	.A(n263));
   MUX2_X1 U245 (.Z(B[27]), 
	.S(SH[0]), 
	.B(n265), 
	.A(n261));
   INV_X1 U246 (.ZN(n261), 
	.A(n266));
   MUX2_X1 U247 (.Z(n266), 
	.S(SH[2]), 
	.B(n268), 
	.A(n267));
   MUX2_X1 U248 (.Z(B[26]), 
	.S(SH[0]), 
	.B(n269), 
	.A(n265));
   INV_X1 U249 (.ZN(n265), 
	.A(n270));
   MUX2_X1 U250 (.Z(n270), 
	.S(SH[2]), 
	.B(n271), 
	.A(n250));
   MUX2_X1 U251 (.Z(n250), 
	.S(SH[3]), 
	.B(n272), 
	.A(n256));
   MUX2_X1 U252 (.Z(n256), 
	.S(SH[1]), 
	.B(n274), 
	.A(n273));
   MUX2_X1 U253 (.Z(B[25]), 
	.S(SH[0]), 
	.B(n275), 
	.A(n269));
   INV_X1 U254 (.ZN(n269), 
	.A(n276));
   MUX2_X1 U255 (.Z(n276), 
	.S(SH[2]), 
	.B(n277), 
	.A(n260));
   MUX2_X1 U256 (.Z(n260), 
	.S(SH[3]), 
	.B(n279), 
	.A(n278));
   MUX2_X1 U257 (.Z(B[24]), 
	.S(SH[0]), 
	.B(n280), 
	.A(n275));
   INV_X1 U258 (.ZN(n275), 
	.A(n281));
   MUX2_X1 U259 (.Z(n281), 
	.S(SH[2]), 
	.B(n282), 
	.A(n264));
   MUX2_X1 U260 (.Z(n264), 
	.S(SH[3]), 
	.B(n284), 
	.A(n283));
   MUX2_X1 U261 (.Z(B[23]), 
	.S(SH[0]), 
	.B(n285), 
	.A(n280));
   INV_X1 U262 (.ZN(n280), 
	.A(n286));
   MUX2_X1 U263 (.Z(n286), 
	.S(SH[2]), 
	.B(n287), 
	.A(n268));
   MUX2_X1 U264 (.Z(n268), 
	.S(SH[3]), 
	.B(n289), 
	.A(n288));
   MUX2_X1 U265 (.Z(B[22]), 
	.S(SH[0]), 
	.B(n290), 
	.A(n285));
   INV_X1 U266 (.ZN(n285), 
	.A(n291));
   MUX2_X1 U267 (.Z(n291), 
	.S(SH[2]), 
	.B(n292), 
	.A(n271));
   MUX2_X1 U268 (.Z(n271), 
	.S(SH[3]), 
	.B(n293), 
	.A(n254));
   MUX2_X1 U269 (.Z(n254), 
	.S(SH[1]), 
	.B(n295), 
	.A(n294));
   MUX2_X1 U270 (.Z(B[21]), 
	.S(SH[0]), 
	.B(n296), 
	.A(n290));
   INV_X1 U271 (.ZN(n290), 
	.A(n297));
   MUX2_X1 U272 (.Z(n297), 
	.S(SH[2]), 
	.B(n298), 
	.A(n277));
   MUX2_X1 U273 (.Z(n277), 
	.S(SH[3]), 
	.B(n300), 
	.A(n299));
   MUX2_X1 U274 (.Z(B[20]), 
	.S(SH[0]), 
	.B(n301), 
	.A(n296));
   INV_X1 U275 (.ZN(n296), 
	.A(n302));
   MUX2_X1 U276 (.Z(n302), 
	.S(SH[2]), 
	.B(n303), 
	.A(n282));
   MUX2_X1 U277 (.Z(n282), 
	.S(SH[3]), 
	.B(n305), 
	.A(n304));
   MUX2_X1 U278 (.Z(B[1]), 
	.S(SH[0]), 
	.B(n306), 
	.A(n251));
   INV_X1 U279 (.ZN(n251), 
	.A(n307));
   MUX2_X1 U280 (.Z(n307), 
	.S(SH[2]), 
	.B(n259), 
	.A(n234));
   MUX2_X1 U281 (.Z(n259), 
	.S(SH[3]), 
	.B(n299), 
	.A(n308));
   MUX2_X1 U282 (.Z(n299), 
	.S(SH[1]), 
	.B(n310), 
	.A(n309));
   MUX2_X1 U283 (.Z(n234), 
	.S(SH[3]), 
	.B(n278), 
	.A(n311));
   MUX2_X1 U284 (.Z(n278), 
	.S(SH[1]), 
	.B(n313), 
	.A(n312));
   MUX2_X1 U285 (.Z(B[19]), 
	.S(SH[0]), 
	.B(n314), 
	.A(n301));
   INV_X1 U286 (.ZN(n301), 
	.A(n315));
   MUX2_X1 U287 (.Z(n315), 
	.S(SH[2]), 
	.B(n316), 
	.A(n287));
   MUX2_X1 U288 (.Z(n287), 
	.S(SH[3]), 
	.B(n318), 
	.A(n317));
   MUX2_X1 U289 (.Z(B[18]), 
	.S(SH[0]), 
	.B(n319), 
	.A(n314));
   INV_X1 U290 (.ZN(n314), 
	.A(n320));
   MUX2_X1 U291 (.Z(n320), 
	.S(SH[2]), 
	.B(n321), 
	.A(n292));
   MUX2_X1 U292 (.Z(n292), 
	.S(SH[3]), 
	.B(n322), 
	.A(n272));
   MUX2_X1 U293 (.Z(n272), 
	.S(SH[1]), 
	.B(n324), 
	.A(n323));
   MUX2_X1 U294 (.Z(B[17]), 
	.S(SH[0]), 
	.B(n325), 
	.A(n319));
   INV_X1 U295 (.ZN(n319), 
	.A(n326));
   MUX2_X1 U296 (.Z(n326), 
	.S(SH[2]), 
	.B(n327), 
	.A(n298));
   MUX2_X1 U297 (.Z(n298), 
	.S(SH[3]), 
	.B(n328), 
	.A(n279));
   MUX2_X1 U298 (.Z(n279), 
	.S(SH[1]), 
	.B(n330), 
	.A(n329));
   MUX2_X1 U299 (.Z(B[16]), 
	.S(SH[0]), 
	.B(n331), 
	.A(n325));
   INV_X1 U300 (.ZN(n325), 
	.A(n332));
   MUX2_X1 U301 (.Z(n332), 
	.S(SH[2]), 
	.B(n333), 
	.A(n303));
   MUX2_X1 U302 (.Z(n303), 
	.S(SH[3]), 
	.B(n334), 
	.A(n284));
   MUX2_X1 U303 (.Z(n284), 
	.S(SH[1]), 
	.B(n335), 
	.A(n324));
   MUX2_X1 U304 (.Z(n324), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n337), 
	.A(n336));
   MUX2_X1 U305 (.Z(B[15]), 
	.S(SH[0]), 
	.B(n338), 
	.A(n331));
   INV_X1 U306 (.ZN(n331), 
	.A(n339));
   MUX2_X1 U307 (.Z(n339), 
	.S(SH[2]), 
	.B(n340), 
	.A(n316));
   MUX2_X1 U308 (.Z(n316), 
	.S(SH[3]), 
	.B(n341), 
	.A(n289));
   MUX2_X1 U309 (.Z(n289), 
	.S(SH[1]), 
	.B(n342), 
	.A(n330));
   MUX2_X1 U310 (.Z(n330), 
	.S(SH[4]), 
	.B(n344), 
	.A(n343));
   MUX2_X1 U311 (.Z(B[14]), 
	.S(SH[0]), 
	.B(n345), 
	.A(n338));
   INV_X1 U312 (.ZN(n338), 
	.A(n346));
   MUX2_X1 U313 (.Z(n346), 
	.S(SH[2]), 
	.B(n347), 
	.A(n321));
   MUX2_X1 U314 (.Z(n321), 
	.S(SH[3]), 
	.B(n348), 
	.A(n293));
   MUX2_X1 U315 (.Z(n293), 
	.S(SH[1]), 
	.B(n349), 
	.A(n335));
   MUX2_X1 U316 (.Z(n335), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n351), 
	.A(n350));
   MUX2_X1 U317 (.Z(B[13]), 
	.S(SH[0]), 
	.B(n352), 
	.A(n345));
   INV_X1 U318 (.ZN(n345), 
	.A(n353));
   MUX2_X1 U319 (.Z(n353), 
	.S(SH[2]), 
	.B(n354), 
	.A(n327));
   MUX2_X1 U320 (.Z(n327), 
	.S(SH[3]), 
	.B(n355), 
	.A(n300));
   MUX2_X1 U321 (.Z(n300), 
	.S(SH[1]), 
	.B(n356), 
	.A(n342));
   MUX2_X1 U322 (.Z(n342), 
	.S(SH[4]), 
	.B(n358), 
	.A(n357));
   MUX2_X1 U323 (.Z(B[12]), 
	.S(SH[0]), 
	.B(n359), 
	.A(n352));
   INV_X1 U324 (.ZN(n352), 
	.A(n360));
   MUX2_X1 U325 (.Z(n360), 
	.S(SH[2]), 
	.B(n221), 
	.A(n333));
   MUX2_X1 U326 (.Z(n221), 
	.S(SH[3]), 
	.B(n361), 
	.A(n334));
   MUX2_X1 U327 (.Z(n334), 
	.S(SH[1]), 
	.B(n363), 
	.A(n362));
   MUX2_X1 U328 (.Z(n333), 
	.S(SH[3]), 
	.B(n238), 
	.A(n305));
   MUX2_X1 U329 (.Z(n238), 
	.S(SH[1]), 
	.B(n365), 
	.A(n364));
   MUX2_X1 U330 (.Z(n305), 
	.S(SH[1]), 
	.B(n366), 
	.A(n349));
   MUX2_X1 U331 (.Z(n349), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n368), 
	.A(n367));
   MUX2_X1 U332 (.Z(B[11]), 
	.S(SH[0]), 
	.B(n369), 
	.A(n359));
   INV_X1 U333 (.ZN(n359), 
	.A(n370));
   MUX2_X1 U334 (.Z(n370), 
	.S(SH[2]), 
	.B(n225), 
	.A(n340));
   MUX2_X1 U335 (.Z(n225), 
	.S(SH[3]), 
	.B(n371), 
	.A(n341));
   MUX2_X1 U336 (.Z(n341), 
	.S(SH[1]), 
	.B(n373), 
	.A(n372));
   MUX2_X1 U337 (.Z(n340), 
	.S(SH[3]), 
	.B(n243), 
	.A(n318));
   MUX2_X1 U338 (.Z(n243), 
	.S(SH[1]), 
	.B(n375), 
	.A(n374));
   MUX2_X1 U339 (.Z(n318), 
	.S(SH[1]), 
	.B(n376), 
	.A(n356));
   MUX2_X1 U340 (.Z(n356), 
	.S(SH[4]), 
	.B(n378), 
	.A(n377));
   MUX2_X1 U341 (.Z(B[10]), 
	.S(SH[0]), 
	.B(n217), 
	.A(n369));
   INV_X1 U342 (.ZN(n217), 
	.A(n379));
   MUX2_X1 U343 (.Z(n379), 
	.S(SH[2]), 
	.B(n233), 
	.A(n354));
   MUX2_X1 U344 (.Z(n233), 
	.S(SH[3]), 
	.B(n308), 
	.A(n355));
   MUX2_X1 U345 (.Z(n308), 
	.S(SH[1]), 
	.B(n381), 
	.A(n380));
   MUX2_X1 U346 (.Z(n355), 
	.S(SH[1]), 
	.B(n374), 
	.A(n373));
   MUX2_X1 U347 (.Z(n374), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n383), 
	.A(n382));
   MUX2_X1 U348 (.Z(n373), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n385), 
	.A(n384));
   MUX2_X1 U349 (.Z(n354), 
	.S(SH[3]), 
	.B(n311), 
	.A(n328));
   MUX2_X1 U350 (.Z(n311), 
	.S(SH[1]), 
	.B(n386), 
	.A(n375));
   MUX2_X1 U351 (.Z(n375), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n388), 
	.A(n387));
   MUX2_X1 U352 (.Z(n328), 
	.S(SH[1]), 
	.B(n372), 
	.A(n376));
   MUX2_X1 U353 (.Z(n372), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n390), 
	.A(n389));
   MUX2_X1 U354 (.Z(n376), 
	.S(SH[4]), 
	.B(n392), 
	.A(n391));
   INV_X1 U355 (.ZN(n369), 
	.A(n393));
   MUX2_X1 U356 (.Z(n393), 
	.S(SH[2]), 
	.B(n229), 
	.A(n347));
   MUX2_X1 U357 (.Z(n229), 
	.S(SH[3]), 
	.B(n253), 
	.A(n348));
   MUX2_X1 U358 (.Z(n253), 
	.S(SH[1]), 
	.B(n395), 
	.A(n394));
   MUX2_X1 U359 (.Z(n348), 
	.S(SH[1]), 
	.B(n364), 
	.A(n363));
   MUX2_X1 U360 (.Z(n364), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n397), 
	.A(n396));
   MUX2_X1 U361 (.Z(n363), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n399), 
	.A(n398));
   MUX2_X1 U362 (.Z(n347), 
	.S(SH[3]), 
	.B(n255), 
	.A(n322));
   MUX2_X1 U363 (.Z(n255), 
	.S(SH[1]), 
	.B(n400), 
	.A(n365));
   MUX2_X1 U364 (.Z(n365), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n402), 
	.A(n401));
   MUX2_X1 U365 (.Z(n322), 
	.S(SH[1]), 
	.B(n362), 
	.A(n366));
   MUX2_X1 U366 (.Z(n362), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n404), 
	.A(n403));
   MUX2_X1 U367 (.Z(n366), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n406), 
	.A(n405));
   MUX2_X1 U368 (.Z(B[0]), 
	.S(SH[0]), 
	.B(n245), 
	.A(n306));
   INV_X1 U369 (.ZN(n245), 
	.A(n407));
   MUX2_X1 U370 (.Z(n407), 
	.S(SH[2]), 
	.B(n267), 
	.A(n242));
   MUX2_X1 U371 (.Z(n267), 
	.S(SH[3]), 
	.B(n317), 
	.A(n244));
   MUX2_X1 U372 (.Z(n317), 
	.S(SH[1]), 
	.B(n329), 
	.A(n310));
   MUX2_X1 U373 (.Z(n329), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n387), 
	.A(n388));
   MUX2_X1 U374 (.Z(n310), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n382), 
	.A(n383));
   MUX2_X1 U375 (.Z(n244), 
	.S(SH[1]), 
	.B(n312), 
	.A(n381));
   MUX2_X1 U376 (.Z(n312), 
	.S(SH[4]), 
	.B(n391), 
	.A(n392));
   MUX2_X1 U377 (.Z(n381), 
	.S(SH[4]), 
	.B(n377), 
	.A(n378));
   MUX2_X1 U378 (.Z(n242), 
	.S(SH[3]), 
	.B(n288), 
	.A(n371));
   MUX2_X1 U379 (.Z(n288), 
	.S(SH[1]), 
	.B(n309), 
	.A(n313));
   MUX2_X1 U380 (.Z(n309), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n384), 
	.A(n385));
   MUX2_X1 U381 (.Z(n313), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n389), 
	.A(n390));
   MUX2_X1 U382 (.Z(n371), 
	.S(SH[1]), 
	.B(n380), 
	.A(n386));
   MUX2_X1 U383 (.Z(n380), 
	.S(SH[4]), 
	.B(n357), 
	.A(n358));
   MUX2_X1 U384 (.Z(n386), 
	.S(SH[4]), 
	.B(n343), 
	.A(n344));
   INV_X1 U385 (.ZN(n344), 
	.A(A[31]));
   INV_X1 U386 (.ZN(n306), 
	.A(n408));
   MUX2_X1 U387 (.Z(n408), 
	.S(SH[2]), 
	.B(n263), 
	.A(n237));
   MUX2_X1 U388 (.Z(n263), 
	.S(SH[3]), 
	.B(n304), 
	.A(n239));
   MUX2_X1 U389 (.Z(n304), 
	.S(SH[1]), 
	.B(n323), 
	.A(n295));
   MUX2_X1 U390 (.Z(n323), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n401), 
	.A(n402));
   MUX2_X1 U391 (.Z(n295), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n396), 
	.A(n397));
   MUX2_X1 U392 (.Z(n239), 
	.S(SH[1]), 
	.B(n273), 
	.A(n395));
   MUX2_X1 U393 (.Z(n273), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n405), 
	.A(n406));
   MUX2_X1 U394 (.Z(n395), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n367), 
	.A(n368));
   MUX2_X1 U395 (.Z(n237), 
	.S(SH[3]), 
	.B(n283), 
	.A(n361));
   MUX2_X1 U396 (.Z(n283), 
	.S(SH[1]), 
	.B(n294), 
	.A(n274));
   MUX2_X1 U397 (.Z(n294), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n398), 
	.A(n399));
   MUX2_X1 U398 (.Z(n274), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n403), 
	.A(n404));
   MUX2_X1 U399 (.Z(n361), 
	.S(SH[1]), 
	.B(n394), 
	.A(n400));
   MUX2_X1 U400 (.Z(n394), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n350), 
	.A(n351));
   MUX2_X1 U401 (.Z(n400), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n336), 
	.A(n337));
endmodule

module up_island_DW_rbsh_1 (
	A, 
	SH, 
	B, 
	SH_TC, 
	FE_OFN176_UUT_Mpath_out_regB_1_, 
	FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_, 
	FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_);
   input [31:0] A;
   input [4:0] SH;
   output [31:0] B;
   input SH_TC;
   input FE_OFN176_UUT_Mpath_out_regB_1_;
   input FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_;
   input FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_;

   // Internal wires
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;

   INV_X1 U164 (.ZN(n404), 
	.A(A[18]));
   INV_X1 U165 (.ZN(n338), 
	.A(A[15]));
   INV_X1 U166 (.ZN(n390), 
	.A(A[19]));
   INV_X1 U167 (.ZN(n402), 
	.A(A[20]));
   INV_X1 U168 (.ZN(n388), 
	.A(A[21]));
   INV_X1 U169 (.ZN(n382), 
	.A(A[9]));
   INV_X1 U170 (.ZN(n374), 
	.A(A[10]));
   INV_X1 U171 (.ZN(n397), 
	.A(A[22]));
   INV_X1 U172 (.ZN(n383), 
	.A(A[23]));
   INV_X1 U173 (.ZN(n396), 
	.A(A[8]));
   INV_X1 U174 (.ZN(n400), 
	.A(A[16]));
   INV_X1 U175 (.ZN(n386), 
	.A(A[17]));
   INV_X1 U176 (.ZN(n358), 
	.A(A[28]));
   INV_X1 U177 (.ZN(n363), 
	.A(A[27]));
   INV_X1 U178 (.ZN(n381), 
	.A(A[25]));
   INV_X1 U179 (.ZN(n344), 
	.A(A[30]));
   INV_X1 U180 (.ZN(n384), 
	.A(A[7]));
   INV_X1 U181 (.ZN(n345), 
	.A(A[14]));
   INV_X1 U182 (.ZN(n352), 
	.A(A[13]));
   INV_X1 U183 (.ZN(n364), 
	.A(A[11]));
   INV_X1 U184 (.ZN(n359), 
	.A(A[12]));
   INV_X1 U185 (.ZN(n351), 
	.A(A[29]));
   INV_X1 U186 (.ZN(n389), 
	.A(A[5]));
   INV_X1 U187 (.ZN(n373), 
	.A(A[26]));
   INV_X1 U188 (.ZN(n395), 
	.A(A[24]));
   INV_X1 U189 (.ZN(n398), 
	.A(A[6]));
   INV_X1 U190 (.ZN(n403), 
	.A(A[4]));
   INV_X1 U191 (.ZN(n391), 
	.A(A[3]));
   INV_X1 U192 (.ZN(n405), 
	.A(A[2]));
   INV_X1 U193 (.ZN(n401), 
	.A(A[0]));
   INV_X1 U194 (.ZN(n387), 
	.A(A[1]));
   MUX2_X1 U210 (.Z(B[9]), 
	.S(SH[0]), 
	.B(n219), 
	.A(n218));
   MUX2_X1 U211 (.Z(B[8]), 
	.S(SH[0]), 
	.B(n218), 
	.A(n220));
   INV_X1 U212 (.ZN(n218), 
	.A(n221));
   MUX2_X1 U213 (.Z(n221), 
	.S(SH[2]), 
	.B(n223), 
	.A(n222));
   MUX2_X1 U214 (.Z(B[7]), 
	.S(SH[0]), 
	.B(n220), 
	.A(n224));
   INV_X1 U215 (.ZN(n220), 
	.A(n225));
   MUX2_X1 U216 (.Z(n225), 
	.S(SH[2]), 
	.B(n227), 
	.A(n226));
   MUX2_X1 U217 (.Z(B[6]), 
	.S(SH[0]), 
	.B(n224), 
	.A(n228));
   INV_X1 U218 (.ZN(n224), 
	.A(n229));
   MUX2_X1 U219 (.Z(n229), 
	.S(SH[2]), 
	.B(n231), 
	.A(n230));
   MUX2_X1 U220 (.Z(B[5]), 
	.S(SH[0]), 
	.B(n228), 
	.A(n232));
   INV_X1 U221 (.ZN(n228), 
	.A(n233));
   MUX2_X1 U222 (.Z(n233), 
	.S(SH[2]), 
	.B(n235), 
	.A(n234));
   MUX2_X1 U223 (.Z(B[4]), 
	.S(SH[0]), 
	.B(n232), 
	.A(n236));
   INV_X1 U224 (.ZN(n232), 
	.A(n237));
   MUX2_X1 U225 (.Z(n237), 
	.S(SH[2]), 
	.B(n222), 
	.A(n238));
   MUX2_X1 U226 (.Z(n222), 
	.S(SH[3]), 
	.B(n240), 
	.A(n239));
   MUX2_X1 U227 (.Z(B[3]), 
	.S(SH[0]), 
	.B(n236), 
	.A(n241));
   INV_X1 U228 (.ZN(n236), 
	.A(n242));
   MUX2_X1 U229 (.Z(n242), 
	.S(SH[2]), 
	.B(n226), 
	.A(n243));
   MUX2_X1 U230 (.Z(n226), 
	.S(SH[3]), 
	.B(n245), 
	.A(n244));
   MUX2_X1 U231 (.Z(B[31]), 
	.S(SH[0]), 
	.B(n247), 
	.A(n246));
   MUX2_X1 U232 (.Z(B[30]), 
	.S(SH[0]), 
	.B(n246), 
	.A(n248));
   INV_X1 U233 (.ZN(n246), 
	.A(n249));
   MUX2_X1 U234 (.Z(n249), 
	.S(SH[2]), 
	.B(n251), 
	.A(n250));
   MUX2_X1 U235 (.Z(B[2]), 
	.S(SH[0]), 
	.B(n241), 
	.A(n252));
   INV_X1 U236 (.ZN(n241), 
	.A(n253));
   MUX2_X1 U237 (.Z(n253), 
	.S(SH[2]), 
	.B(n230), 
	.A(n251));
   MUX2_X1 U238 (.Z(n230), 
	.S(SH[3]), 
	.B(n255), 
	.A(n254));
   MUX2_X1 U239 (.Z(n251), 
	.S(SH[3]), 
	.B(n257), 
	.A(n256));
   MUX2_X1 U240 (.Z(B[29]), 
	.S(SH[0]), 
	.B(n248), 
	.A(n258));
   INV_X1 U241 (.ZN(n248), 
	.A(n259));
   MUX2_X1 U242 (.Z(n259), 
	.S(SH[2]), 
	.B(n261), 
	.A(n260));
   MUX2_X1 U243 (.Z(B[28]), 
	.S(SH[0]), 
	.B(n258), 
	.A(n262));
   INV_X1 U244 (.ZN(n258), 
	.A(n263));
   MUX2_X1 U245 (.Z(n263), 
	.S(SH[2]), 
	.B(n265), 
	.A(n264));
   MUX2_X1 U246 (.Z(B[27]), 
	.S(SH[0]), 
	.B(n262), 
	.A(n266));
   INV_X1 U247 (.ZN(n262), 
	.A(n267));
   MUX2_X1 U248 (.Z(n267), 
	.S(SH[2]), 
	.B(n269), 
	.A(n268));
   MUX2_X1 U249 (.Z(B[26]), 
	.S(SH[0]), 
	.B(n266), 
	.A(n270));
   INV_X1 U250 (.ZN(n266), 
	.A(n271));
   MUX2_X1 U251 (.Z(n271), 
	.S(SH[2]), 
	.B(n250), 
	.A(n272));
   MUX2_X1 U252 (.Z(n250), 
	.S(SH[3]), 
	.B(n254), 
	.A(n273));
   MUX2_X1 U253 (.Z(n254), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n275), 
	.A(n274));
   MUX2_X1 U254 (.Z(B[25]), 
	.S(SH[0]), 
	.B(n270), 
	.A(n276));
   INV_X1 U255 (.ZN(n270), 
	.A(n277));
   MUX2_X1 U256 (.Z(n277), 
	.S(SH[2]), 
	.B(n260), 
	.A(n278));
   MUX2_X1 U257 (.Z(n260), 
	.S(SH[3]), 
	.B(n280), 
	.A(n279));
   MUX2_X1 U258 (.Z(B[24]), 
	.S(SH[0]), 
	.B(n276), 
	.A(n281));
   INV_X1 U259 (.ZN(n276), 
	.A(n282));
   MUX2_X1 U260 (.Z(n282), 
	.S(SH[2]), 
	.B(n264), 
	.A(n283));
   MUX2_X1 U261 (.Z(n264), 
	.S(SH[3]), 
	.B(n285), 
	.A(n284));
   MUX2_X1 U262 (.Z(B[23]), 
	.S(SH[0]), 
	.B(n281), 
	.A(n286));
   INV_X1 U263 (.ZN(n281), 
	.A(n287));
   MUX2_X1 U264 (.Z(n287), 
	.S(SH[2]), 
	.B(n268), 
	.A(n288));
   MUX2_X1 U265 (.Z(n268), 
	.S(SH[3]), 
	.B(n290), 
	.A(n289));
   MUX2_X1 U266 (.Z(B[22]), 
	.S(SH[0]), 
	.B(n286), 
	.A(n291));
   INV_X1 U267 (.ZN(n286), 
	.A(n292));
   MUX2_X1 U268 (.Z(n292), 
	.S(SH[2]), 
	.B(n272), 
	.A(n293));
   MUX2_X1 U269 (.Z(n272), 
	.S(SH[3]), 
	.B(n256), 
	.A(n294));
   MUX2_X1 U270 (.Z(n256), 
	.S(FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n296), 
	.A(n295));
   MUX2_X1 U271 (.Z(B[21]), 
	.S(SH[0]), 
	.B(n291), 
	.A(n297));
   INV_X1 U272 (.ZN(n291), 
	.A(n298));
   MUX2_X1 U273 (.Z(n298), 
	.S(SH[2]), 
	.B(n278), 
	.A(n299));
   MUX2_X1 U274 (.Z(n278), 
	.S(SH[3]), 
	.B(n301), 
	.A(n300));
   MUX2_X1 U275 (.Z(B[20]), 
	.S(SH[0]), 
	.B(n297), 
	.A(n302));
   INV_X1 U276 (.ZN(n297), 
	.A(n303));
   MUX2_X1 U277 (.Z(n303), 
	.S(SH[2]), 
	.B(n283), 
	.A(n304));
   MUX2_X1 U278 (.Z(n283), 
	.S(SH[3]), 
	.B(n306), 
	.A(n305));
   MUX2_X1 U279 (.Z(B[1]), 
	.S(SH[0]), 
	.B(n252), 
	.A(n307));
   INV_X1 U280 (.ZN(n252), 
	.A(n308));
   MUX2_X1 U281 (.Z(n308), 
	.S(SH[2]), 
	.B(n234), 
	.A(n261));
   MUX2_X1 U282 (.Z(n234), 
	.S(SH[3]), 
	.B(n309), 
	.A(n280));
   MUX2_X1 U283 (.Z(n280), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n311), 
	.A(n310));
   MUX2_X1 U284 (.Z(n261), 
	.S(SH[3]), 
	.B(n312), 
	.A(n301));
   MUX2_X1 U285 (.Z(n301), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n314), 
	.A(n313));
   MUX2_X1 U286 (.Z(B[19]), 
	.S(SH[0]), 
	.B(n302), 
	.A(n315));
   INV_X1 U287 (.ZN(n302), 
	.A(n316));
   MUX2_X1 U288 (.Z(n316), 
	.S(SH[2]), 
	.B(n288), 
	.A(n317));
   MUX2_X1 U289 (.Z(n288), 
	.S(SH[3]), 
	.B(n319), 
	.A(n318));
   MUX2_X1 U290 (.Z(B[18]), 
	.S(SH[0]), 
	.B(n315), 
	.A(n320));
   INV_X1 U291 (.ZN(n315), 
	.A(n321));
   MUX2_X1 U292 (.Z(n321), 
	.S(SH[2]), 
	.B(n293), 
	.A(n322));
   MUX2_X1 U293 (.Z(n293), 
	.S(SH[3]), 
	.B(n273), 
	.A(n323));
   MUX2_X1 U294 (.Z(n273), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n325), 
	.A(n324));
   MUX2_X1 U295 (.Z(B[17]), 
	.S(SH[0]), 
	.B(n320), 
	.A(n326));
   INV_X1 U296 (.ZN(n320), 
	.A(n327));
   MUX2_X1 U297 (.Z(n327), 
	.S(SH[2]), 
	.B(n299), 
	.A(n328));
   MUX2_X1 U298 (.Z(n299), 
	.S(SH[3]), 
	.B(n279), 
	.A(n329));
   MUX2_X1 U299 (.Z(n279), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n331), 
	.A(n330));
   MUX2_X1 U300 (.Z(B[16]), 
	.S(SH[0]), 
	.B(n326), 
	.A(n332));
   INV_X1 U301 (.ZN(n326), 
	.A(n333));
   MUX2_X1 U302 (.Z(n333), 
	.S(SH[2]), 
	.B(n304), 
	.A(n334));
   MUX2_X1 U303 (.Z(n304), 
	.S(SH[3]), 
	.B(n284), 
	.A(n335));
   MUX2_X1 U304 (.Z(n284), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n324), 
	.A(n336));
   MUX2_X1 U305 (.Z(n324), 
	.S(SH[4]), 
	.B(n338), 
	.A(n337));
   MUX2_X1 U306 (.Z(B[15]), 
	.S(SH[0]), 
	.B(n332), 
	.A(n339));
   INV_X1 U307 (.ZN(n332), 
	.A(n340));
   MUX2_X1 U308 (.Z(n340), 
	.S(SH[2]), 
	.B(n317), 
	.A(n341));
   MUX2_X1 U309 (.Z(n317), 
	.S(SH[3]), 
	.B(n289), 
	.A(n342));
   MUX2_X1 U310 (.Z(n289), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n330), 
	.A(n343));
   MUX2_X1 U311 (.Z(n330), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n345), 
	.A(n344));
   MUX2_X1 U312 (.Z(B[14]), 
	.S(SH[0]), 
	.B(n339), 
	.A(n346));
   INV_X1 U313 (.ZN(n339), 
	.A(n347));
   MUX2_X1 U314 (.Z(n347), 
	.S(SH[2]), 
	.B(n322), 
	.A(n348));
   MUX2_X1 U315 (.Z(n322), 
	.S(SH[3]), 
	.B(n294), 
	.A(n349));
   MUX2_X1 U316 (.Z(n294), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n336), 
	.A(n350));
   MUX2_X1 U317 (.Z(n336), 
	.S(SH[4]), 
	.B(n352), 
	.A(n351));
   MUX2_X1 U318 (.Z(B[13]), 
	.S(SH[0]), 
	.B(n346), 
	.A(n353));
   INV_X1 U319 (.ZN(n346), 
	.A(n354));
   MUX2_X1 U320 (.Z(n354), 
	.S(SH[2]), 
	.B(n328), 
	.A(n355));
   MUX2_X1 U321 (.Z(n328), 
	.S(SH[3]), 
	.B(n300), 
	.A(n356));
   MUX2_X1 U322 (.Z(n300), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n343), 
	.A(n357));
   MUX2_X1 U323 (.Z(n343), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n359), 
	.A(n358));
   MUX2_X1 U324 (.Z(B[12]), 
	.S(SH[0]), 
	.B(n353), 
	.A(n360));
   INV_X1 U325 (.ZN(n353), 
	.A(n361));
   MUX2_X1 U326 (.Z(n361), 
	.S(SH[2]), 
	.B(n334), 
	.A(n223));
   MUX2_X1 U327 (.Z(n334), 
	.S(SH[3]), 
	.B(n305), 
	.A(n240));
   MUX2_X1 U328 (.Z(n305), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n350), 
	.A(n362));
   MUX2_X1 U329 (.Z(n350), 
	.S(SH[4]), 
	.B(n364), 
	.A(n363));
   MUX2_X1 U330 (.Z(n240), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n366), 
	.A(n365));
   MUX2_X1 U331 (.Z(n223), 
	.S(SH[3]), 
	.B(n335), 
	.A(n367));
   MUX2_X1 U332 (.Z(n335), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n369), 
	.A(n368));
   MUX2_X1 U333 (.Z(B[11]), 
	.S(SH[0]), 
	.B(n360), 
	.A(n370));
   INV_X1 U334 (.ZN(n360), 
	.A(n371));
   MUX2_X1 U335 (.Z(n371), 
	.S(SH[2]), 
	.B(n341), 
	.A(n227));
   MUX2_X1 U336 (.Z(n341), 
	.S(SH[3]), 
	.B(n318), 
	.A(n245));
   MUX2_X1 U337 (.Z(n318), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n357), 
	.A(n372));
   MUX2_X1 U338 (.Z(n357), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n374), 
	.A(n373));
   MUX2_X1 U339 (.Z(n245), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n376), 
	.A(n375));
   MUX2_X1 U340 (.Z(n227), 
	.S(SH[3]), 
	.B(n342), 
	.A(n377));
   MUX2_X1 U341 (.Z(n342), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n379), 
	.A(n378));
   MUX2_X1 U342 (.Z(B[10]), 
	.S(SH[0]), 
	.B(n370), 
	.A(n219));
   INV_X1 U343 (.ZN(n370), 
	.A(n380));
   MUX2_X1 U344 (.Z(n380), 
	.S(SH[2]), 
	.B(n348), 
	.A(n231));
   MUX2_X1 U345 (.Z(n348), 
	.S(SH[3]), 
	.B(n323), 
	.A(n255));
   MUX2_X1 U346 (.Z(n323), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n362), 
	.A(n369));
   MUX2_X1 U347 (.Z(n362), 
	.S(SH[4]), 
	.B(n382), 
	.A(n381));
   MUX2_X1 U348 (.Z(n369), 
	.S(SH[4]), 
	.B(n384), 
	.A(n383));
   MUX2_X1 U349 (.Z(n255), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n365), 
	.A(n385));
   MUX2_X1 U350 (.Z(n365), 
	.S(SH[4]), 
	.B(n387), 
	.A(n386));
   MUX2_X1 U351 (.Z(n231), 
	.S(SH[3]), 
	.B(n349), 
	.A(n257));
   MUX2_X1 U352 (.Z(n349), 
	.S(SH[1]), 
	.B(n368), 
	.A(n366));
   MUX2_X1 U353 (.Z(n368), 
	.S(SH[4]), 
	.B(n389), 
	.A(n388));
   MUX2_X1 U354 (.Z(n366), 
	.S(SH[4]), 
	.B(n391), 
	.A(n390));
   MUX2_X1 U355 (.Z(n257), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n393), 
	.A(n392));
   INV_X1 U356 (.ZN(n219), 
	.A(n394));
   MUX2_X1 U357 (.Z(n394), 
	.S(SH[2]), 
	.B(n355), 
	.A(n235));
   MUX2_X1 U358 (.Z(n355), 
	.S(SH[3]), 
	.B(n329), 
	.A(n309));
   MUX2_X1 U359 (.Z(n329), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n372), 
	.A(n379));
   MUX2_X1 U360 (.Z(n372), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n396), 
	.A(n395));
   MUX2_X1 U361 (.Z(n379), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n398), 
	.A(n397));
   MUX2_X1 U362 (.Z(n309), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n375), 
	.A(n399));
   MUX2_X1 U363 (.Z(n375), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n401), 
	.A(n400));
   MUX2_X1 U364 (.Z(n235), 
	.S(SH[3]), 
	.B(n356), 
	.A(n312));
   MUX2_X1 U365 (.Z(n356), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n378), 
	.A(n376));
   MUX2_X1 U366 (.Z(n378), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n403), 
	.A(n402));
   MUX2_X1 U367 (.Z(n376), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n405), 
	.A(n404));
   MUX2_X1 U368 (.Z(n312), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n407), 
	.A(n406));
   MUX2_X1 U369 (.Z(B[0]), 
	.S(SH[0]), 
	.B(n307), 
	.A(n247));
   INV_X1 U370 (.ZN(n307), 
	.A(n408));
   MUX2_X1 U371 (.Z(n408), 
	.S(SH[2]), 
	.B(n238), 
	.A(n265));
   MUX2_X1 U372 (.Z(n238), 
	.S(SH[3]), 
	.B(n367), 
	.A(n285));
   MUX2_X1 U373 (.Z(n367), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n385), 
	.A(n393));
   MUX2_X1 U374 (.Z(n385), 
	.S(SH[4]), 
	.B(n337), 
	.A(n338));
   INV_X1 U375 (.ZN(n337), 
	.A(A[31]));
   MUX2_X1 U376 (.Z(n393), 
	.S(SH[4]), 
	.B(n351), 
	.A(n352));
   MUX2_X1 U377 (.Z(n285), 
	.S(FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n274), 
	.A(n296));
   MUX2_X1 U378 (.Z(n274), 
	.S(SH[4]), 
	.B(n383), 
	.A(n384));
   MUX2_X1 U379 (.Z(n296), 
	.S(SH[4]), 
	.B(n388), 
	.A(n389));
   MUX2_X1 U380 (.Z(n265), 
	.S(SH[3]), 
	.B(n239), 
	.A(n306));
   MUX2_X1 U381 (.Z(n239), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n392), 
	.A(n275));
   MUX2_X1 U382 (.Z(n392), 
	.S(SH[4]), 
	.B(n363), 
	.A(n364));
   MUX2_X1 U383 (.Z(n275), 
	.S(SH[4]), 
	.B(n381), 
	.A(n382));
   MUX2_X1 U384 (.Z(n306), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n295), 
	.A(n325));
   MUX2_X1 U385 (.Z(n295), 
	.S(SH[4]), 
	.B(n390), 
	.A(n391));
   MUX2_X1 U386 (.Z(n325), 
	.S(SH[4]), 
	.B(n386), 
	.A(n387));
   INV_X1 U387 (.ZN(n247), 
	.A(n409));
   MUX2_X1 U388 (.Z(n409), 
	.S(SH[2]), 
	.B(n243), 
	.A(n269));
   MUX2_X1 U389 (.Z(n243), 
	.S(SH[3]), 
	.B(n377), 
	.A(n290));
   MUX2_X1 U390 (.Z(n377), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n399), 
	.A(n407));
   MUX2_X1 U391 (.Z(n399), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n344), 
	.A(n345));
   MUX2_X1 U392 (.Z(n407), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n358), 
	.A(n359));
   MUX2_X1 U393 (.Z(n290), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n310), 
	.A(n314));
   MUX2_X1 U394 (.Z(n310), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n397), 
	.A(n398));
   MUX2_X1 U395 (.Z(n314), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n402), 
	.A(n403));
   MUX2_X1 U396 (.Z(n269), 
	.S(SH[3]), 
	.B(n244), 
	.A(n319));
   MUX2_X1 U397 (.Z(n244), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n406), 
	.A(n311));
   MUX2_X1 U398 (.Z(n406), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n373), 
	.A(n374));
   MUX2_X1 U399 (.Z(n311), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n395), 
	.A(n396));
   MUX2_X1 U400 (.Z(n319), 
	.S(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.B(n313), 
	.A(n331));
   MUX2_X1 U401 (.Z(n313), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n404), 
	.A(n405));
   MUX2_X1 U402 (.Z(n331), 
	.S(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n400), 
	.A(n401));
endmodule

module up_island_DW_sra_1 (
	A, 
	SH, 
	B, 
	SH_TC, 
	FE_OFN160_UUT_Mpath_out_regB_4_, 
	FE_OFN164_UUT_Mpath_out_regB_3_, 
	FE_OFN180_UUT_Mpath_out_regB_0_, 
	FE_OFN181_UUT_Mpath_out_regB_0_, 
	FE_OFN184_UUT_Mpath_out_regB_0_, 
	FE_OFN185_UUT_Mpath_out_regB_0_, 
	FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_);
   input [31:0] A;
   input [4:0] SH;
   output [31:0] B;
   input SH_TC;
   input FE_OFN160_UUT_Mpath_out_regB_4_;
   input FE_OFN164_UUT_Mpath_out_regB_3_;
   input FE_OFN180_UUT_Mpath_out_regB_0_;
   input FE_OFN181_UUT_Mpath_out_regB_0_;
   input FE_OFN184_UUT_Mpath_out_regB_0_;
   input FE_OFN185_UUT_Mpath_out_regB_0_;
   input FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_;

   // Internal wires
   wire FE_OFN183_UUT_Mpath_out_regB_0_;
   wire \A[31] ;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1491;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;

   assign B[31] = \A[31]  ;
   assign \A[31]  = A[31] ;

   CLKBUF_X1 FE_OFC183_UUT_Mpath_out_regB_0_ (.Z(FE_OFN183_UUT_Mpath_out_regB_0_), 
	.A(SH[0]));
   INV_X1 U170 (.ZN(n1580), 
	.A(A[18]));
   INV_X1 U171 (.ZN(n1592), 
	.A(A[15]));
   INV_X1 U172 (.ZN(n1556), 
	.A(A[19]));
   INV_X1 U173 (.ZN(n1578), 
	.A(A[20]));
   INV_X1 U174 (.ZN(n1554), 
	.A(A[21]));
   INV_X1 U175 (.ZN(n1608), 
	.A(A[9]));
   INV_X1 U176 (.ZN(n1640), 
	.A(A[10]));
   INV_X1 U177 (.ZN(n1568), 
	.A(A[22]));
   INV_X1 U178 (.ZN(n1544), 
	.A(A[23]));
   INV_X1 U179 (.ZN(n1642), 
	.A(A[8]));
   INV_X1 U180 (.ZN(n1572), 
	.A(A[16]));
   INV_X1 U181 (.ZN(n1548), 
	.A(A[17]));
   INV_X1 U182 (.ZN(n1488), 
	.A(A[28]));
   INV_X1 U183 (.ZN(n1502), 
	.A(A[27]));
   INV_X1 U184 (.ZN(n1542), 
	.A(A[25]));
   INV_X1 U185 (.ZN(n1458), 
	.A(A[30]));
   INV_X1 U186 (.ZN(n1598), 
	.A(A[7]));
   INV_X1 U187 (.ZN(n1621), 
	.A(A[14]));
   INV_X1 U188 (.ZN(n1594), 
	.A(A[13]));
   INV_X1 U189 (.ZN(n1606), 
	.A(A[11]));
   INV_X1 U190 (.ZN(n1623), 
	.A(A[12]));
   INV_X1 U191 (.ZN(n1474), 
	.A(A[29]));
   INV_X1 U192 (.ZN(n1600), 
	.A(A[5]));
   INV_X1 U193 (.ZN(n1522), 
	.A(A[26]));
   INV_X1 U194 (.ZN(n1566), 
	.A(A[24]));
   INV_X1 U195 (.ZN(n1627), 
	.A(A[6]));
   INV_X1 U196 (.ZN(n1629), 
	.A(A[4]));
   INV_X1 U197 (.ZN(n1612), 
	.A(A[3]));
   INV_X1 U198 (.ZN(n1635), 
	.A(A[2]));
   INV_X1 U199 (.ZN(n1150), 
	.A(SH[1]));
   INV_X1 U200 (.ZN(n1152), 
	.A(SH[1]));
   INV_X1 U201 (.ZN(n1151), 
	.A(SH[1]));
   INV_X1 U205 (.ZN(n1109), 
	.A(FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_));
   INV_X1 U206 (.ZN(n1110), 
	.A(SH[3]));
   INV_X1 U207 (.ZN(n1111), 
	.A(SH[3]));
   INV_X1 U208 (.ZN(n1112), 
	.A(SH[3]));
   INV_X1 U209 (.ZN(n1113), 
	.A(SH[3]));
   INV_X2 U237 (.ZN(n1141), 
	.A(n1145));
   INV_X1 U238 (.ZN(n1142), 
	.A(n1145));
   INV_X1 U239 (.ZN(n1143), 
	.A(n1145));
   INV_X1 U241 (.ZN(n1145), 
	.A(SH[2]));
   INV_X1 U242 (.ZN(n1146), 
	.A(n1151));
   INV_X1 U243 (.ZN(n1147), 
	.A(n1151));
   INV_X1 U244 (.ZN(n1148), 
	.A(n1151));
   INV_X1 U246 (.ZN(n1153), 
	.A(FE_OFN180_UUT_Mpath_out_regB_0_));
   INV_X1 U247 (.ZN(n1154), 
	.A(FE_OFN183_UUT_Mpath_out_regB_0_));
   INV_X1 U248 (.ZN(n1155), 
	.A(FE_OFN183_UUT_Mpath_out_regB_0_));
   INV_X1 U249 (.ZN(n1156), 
	.A(FE_OFN183_UUT_Mpath_out_regB_0_));
   INV_X1 U250 (.ZN(n1157), 
	.A(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U282 (.ZN(B[9]), 
	.A2(n1190), 
	.A1(n1189));
   MUX2_X1 U283 (.Z(n1190), 
	.S(n1141), 
	.B(n1192), 
	.A(n1191));
   NAND2_X1 U284 (.ZN(n1192), 
	.A2(n1193), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U285 (.ZN(n1191), 
	.A2(n1194), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U286 (.Z(n1189), 
	.S(n1141), 
	.B(n1196), 
	.A(n1195));
   NAND2_X1 U287 (.ZN(n1196), 
	.A2(n1155), 
	.A1(n1197));
   NAND2_X1 U288 (.ZN(n1195), 
	.A2(n1153), 
	.A1(n1198));
   NAND2_X1 U289 (.ZN(B[8]), 
	.A2(n1200), 
	.A1(n1199));
   MUX2_X1 U290 (.Z(n1200), 
	.S(n1141), 
	.B(n1202), 
	.A(n1201));
   NAND2_X1 U291 (.ZN(n1202), 
	.A2(n1197), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U292 (.ZN(n1201), 
	.A2(n1198), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U293 (.Z(n1199), 
	.S(n1141), 
	.B(n1204), 
	.A(n1203));
   NAND2_X1 U294 (.ZN(n1204), 
	.A2(n1153), 
	.A1(n1205));
   NAND2_X1 U295 (.ZN(n1203), 
	.A2(n1153), 
	.A1(n1206));
   NAND2_X1 U296 (.ZN(B[7]), 
	.A2(n1208), 
	.A1(n1207));
   MUX2_X1 U297 (.Z(n1208), 
	.S(n1141), 
	.B(n1210), 
	.A(n1209));
   NAND2_X1 U298 (.ZN(n1210), 
	.A2(n1205), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U299 (.ZN(n1209), 
	.A2(n1206), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U300 (.Z(n1207), 
	.S(n1141), 
	.B(n1212), 
	.A(n1211));
   NAND2_X1 U301 (.ZN(n1212), 
	.A2(n1153), 
	.A1(n1213));
   NAND2_X1 U302 (.ZN(n1211), 
	.A2(n1153), 
	.A1(n1214));
   NAND2_X1 U303 (.ZN(B[6]), 
	.A2(n1216), 
	.A1(n1215));
   MUX2_X1 U304 (.Z(n1216), 
	.S(n1141), 
	.B(n1218), 
	.A(n1217));
   NAND2_X1 U305 (.ZN(n1218), 
	.A2(n1213), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U306 (.ZN(n1217), 
	.A2(n1214), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U307 (.Z(n1215), 
	.S(n1141), 
	.B(n1220), 
	.A(n1219));
   NAND2_X1 U308 (.ZN(n1220), 
	.A2(n1153), 
	.A1(n1194));
   NAND2_X1 U309 (.ZN(n1219), 
	.A2(n1153), 
	.A1(n1221));
   NAND2_X1 U310 (.ZN(B[5]), 
	.A2(n1223), 
	.A1(n1222));
   MUX2_X1 U311 (.Z(n1223), 
	.S(n1141), 
	.B(n1225), 
	.A(n1224));
   NAND2_X1 U312 (.ZN(n1225), 
	.A2(n1194), 
	.A1(FE_OFN181_UUT_Mpath_out_regB_0_));
   NAND2_X1 U313 (.ZN(n1224), 
	.A2(n1221), 
	.A1(FE_OFN185_UUT_Mpath_out_regB_0_));
   MUX2_X1 U314 (.Z(n1222), 
	.S(n1143), 
	.B(n1195), 
	.A(n1226));
   NAND2_X1 U316 (.ZN(n1226), 
	.A2(n1153), 
	.A1(n1228));
   NAND2_X1 U317 (.ZN(B[4]), 
	.A2(n1230), 
	.A1(n1229));
   MUX2_X1 U318 (.Z(n1230), 
	.S(n1143), 
	.B(n1232), 
	.A(n1231));
   NAND2_X1 U319 (.ZN(n1232), 
	.A2(n1198), 
	.A1(FE_OFN184_UUT_Mpath_out_regB_0_));
   NAND2_X1 U320 (.ZN(n1198), 
	.A2(n1234), 
	.A1(n1233));
   MUX2_X1 U321 (.Z(n1234), 
	.S(n1146), 
	.B(n1236), 
	.A(n1235));
   NAND2_X1 U322 (.ZN(n1236), 
	.A2(n1237), 
	.A1(SH[3]));
   NAND2_X1 U323 (.ZN(n1235), 
	.A2(n1238), 
	.A1(SH[3]));
   MUX2_X1 U324 (.Z(n1233), 
	.S(n1146), 
	.B(n1240), 
	.A(n1239));
   NAND2_X1 U325 (.ZN(n1240), 
	.A2(n1110), 
	.A1(n1241));
   NAND2_X1 U326 (.ZN(n1239), 
	.A2(n1109), 
	.A1(n1242));
   NAND2_X1 U327 (.ZN(n1231), 
	.A2(n1228), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U328 (.Z(n1229), 
	.S(n1143), 
	.B(n1203), 
	.A(n1243));
   NAND2_X1 U330 (.ZN(n1243), 
	.A2(n1153), 
	.A1(n1245));
   NAND2_X1 U331 (.ZN(B[3]), 
	.A2(n1247), 
	.A1(n1246));
   MUX2_X1 U332 (.Z(n1247), 
	.S(n1143), 
	.B(n1249), 
	.A(n1248));
   NAND2_X1 U333 (.ZN(n1249), 
	.A2(n1206), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U334 (.ZN(n1206), 
	.A2(n1251), 
	.A1(n1250));
   MUX2_X1 U335 (.Z(n1251), 
	.S(n1146), 
	.B(n1253), 
	.A(n1252));
   NAND2_X1 U336 (.ZN(n1253), 
	.A2(n1254), 
	.A1(SH[3]));
   NAND2_X1 U337 (.ZN(n1252), 
	.A2(n1255), 
	.A1(SH[3]));
   MUX2_X1 U338 (.Z(n1250), 
	.S(n1146), 
	.B(n1257), 
	.A(n1256));
   NAND2_X1 U339 (.ZN(n1257), 
	.A2(n1109), 
	.A1(n1258));
   NAND2_X1 U340 (.ZN(n1256), 
	.A2(n1109), 
	.A1(n1259));
   NAND2_X1 U341 (.ZN(n1248), 
	.A2(n1245), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U342 (.Z(n1246), 
	.S(n1143), 
	.B(n1211), 
	.A(n1260));
   NAND2_X1 U344 (.ZN(n1260), 
	.A2(n1154), 
	.A1(n1262));
   NAND2_X1 U345 (.ZN(B[30]), 
	.A2(n1264), 
	.A1(n1263));
   NAND2_X1 U346 (.ZN(n1264), 
	.A2(\A[31] ), 
	.A1(n1141));
   MUX2_X1 U347 (.Z(n1263), 
	.S(FE_OFN180_UUT_Mpath_out_regB_0_), 
	.B(n1266), 
	.A(n1265));
   NAND2_X1 U348 (.ZN(n1265), 
	.A2(n1145), 
	.A1(n1267));
   NAND2_X1 U349 (.ZN(B[2]), 
	.A2(n1269), 
	.A1(n1268));
   MUX2_X1 U350 (.Z(n1269), 
	.S(n1143), 
	.B(n1271), 
	.A(n1270));
   NAND2_X1 U351 (.ZN(n1271), 
	.A2(n1214), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U352 (.ZN(n1214), 
	.A2(n1273), 
	.A1(n1272));
   MUX2_X1 U353 (.Z(n1273), 
	.S(n1146), 
	.B(n1275), 
	.A(n1274));
   NAND2_X1 U354 (.ZN(n1275), 
	.A2(n1238), 
	.A1(SH[3]));
   NAND2_X1 U355 (.ZN(n1274), 
	.A2(n1276), 
	.A1(SH[3]));
   MUX2_X1 U356 (.Z(n1272), 
	.S(n1148), 
	.B(n1239), 
	.A(n1277));
   NAND2_X1 U358 (.ZN(n1277), 
	.A2(n1109), 
	.A1(n1279));
   NAND2_X1 U359 (.ZN(n1270), 
	.A2(n1262), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U360 (.ZN(n1262), 
	.A2(n1281), 
	.A1(n1280));
   MUX2_X1 U361 (.Z(n1281), 
	.S(n1148), 
	.B(n1283), 
	.A(n1282));
   NAND2_X1 U362 (.ZN(n1283), 
	.A2(n1284), 
	.A1(FE_OFN164_UUT_Mpath_out_regB_3_));
   NAND2_X1 U363 (.ZN(n1282), 
	.A2(n1241), 
	.A1(FE_OFN164_UUT_Mpath_out_regB_3_));
   MUX2_X1 U364 (.Z(n1280), 
	.S(n1148), 
	.B(n1286), 
	.A(n1285));
   NAND2_X1 U365 (.ZN(n1286), 
	.A2(n1109), 
	.A1(n1287));
   NAND2_X1 U366 (.ZN(n1285), 
	.A2(n1109), 
	.A1(n1288));
   MUX2_X1 U367 (.Z(n1268), 
	.S(n1143), 
	.B(n1290), 
	.A(n1289));
   NAND2_X1 U368 (.ZN(n1290), 
	.A2(n1154), 
	.A1(n1221));
   NAND2_X1 U369 (.ZN(n1289), 
	.A2(n1154), 
	.A1(n1291));
   NAND2_X1 U370 (.ZN(B[29]), 
	.A2(n1293), 
	.A1(n1292));
   NAND3_X1 U371 (.ZN(n1293), 
	.A3(n1294), 
	.A2(n1145), 
	.A1(n1157));
   MUX2_X1 U372 (.Z(n1292), 
	.S(n1143), 
	.B(n1266), 
	.A(n1295));
   NAND2_X1 U373 (.ZN(n1295), 
	.A2(n1267), 
	.A1(FE_OFN184_UUT_Mpath_out_regB_0_));
   NAND2_X1 U374 (.ZN(B[28]), 
	.A2(n1297), 
	.A1(n1296));
   NAND3_X1 U375 (.ZN(n1297), 
	.A3(n1298), 
	.A2(n1145), 
	.A1(n1157));
   MUX2_X1 U376 (.Z(n1296), 
	.S(n1143), 
	.B(n1266), 
	.A(n1299));
   NAND2_X1 U377 (.ZN(n1299), 
	.A2(n1294), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U378 (.ZN(B[27]), 
	.A2(n1301), 
	.A1(n1300));
   NAND3_X1 U379 (.ZN(n1301), 
	.A3(n1302), 
	.A2(n1145), 
	.A1(n1157));
   MUX2_X1 U380 (.Z(n1300), 
	.S(n1143), 
	.B(n1266), 
	.A(n1303));
   NAND2_X1 U381 (.ZN(n1303), 
	.A2(n1298), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U382 (.ZN(B[26]), 
	.A2(n1305), 
	.A1(n1304));
   MUX2_X1 U383 (.Z(n1305), 
	.S(n1143), 
	.B(n1307), 
	.A(n1306));
   NAND2_X1 U384 (.ZN(n1307), 
	.A2(\A[31] ), 
	.A1(FE_OFN184_UUT_Mpath_out_regB_0_));
   NAND2_X1 U385 (.ZN(n1306), 
	.A2(n1302), 
	.A1(FE_OFN184_UUT_Mpath_out_regB_0_));
   MUX2_X1 U386 (.Z(n1304), 
	.S(n1143), 
	.B(n1309), 
	.A(n1308));
   NAND2_X1 U387 (.ZN(n1309), 
	.A2(n1154), 
	.A1(n1267));
   NAND2_X1 U388 (.ZN(n1308), 
	.A2(n1154), 
	.A1(n1310));
   NAND2_X1 U389 (.ZN(B[25]), 
	.A2(n1312), 
	.A1(n1311));
   MUX2_X1 U390 (.Z(n1312), 
	.S(n1143), 
	.B(n1314), 
	.A(n1313));
   NAND2_X1 U391 (.ZN(n1314), 
	.A2(n1267), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   OAI21_X1 U392 (.ZN(n1267), 
	.B2(n1150), 
	.B1(n1266), 
	.A(n1315));
   MUX2_X1 U393 (.Z(n1315), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1316));
   NAND2_X1 U394 (.ZN(n1316), 
	.A2(n1150), 
	.A1(n1317));
   NAND2_X1 U395 (.ZN(n1313), 
	.A2(n1310), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U396 (.Z(n1311), 
	.S(n1143), 
	.B(n1319), 
	.A(n1318));
   NAND2_X1 U397 (.ZN(n1319), 
	.A2(n1154), 
	.A1(n1294));
   NAND2_X1 U398 (.ZN(n1318), 
	.A2(n1154), 
	.A1(n1320));
   NAND2_X1 U399 (.ZN(B[24]), 
	.A2(n1322), 
	.A1(n1321));
   MUX2_X1 U400 (.Z(n1322), 
	.S(n1143), 
	.B(n1324), 
	.A(n1323));
   NAND2_X1 U401 (.ZN(n1324), 
	.A2(n1294), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   OAI21_X1 U402 (.ZN(n1294), 
	.B2(n1151), 
	.B1(n1266), 
	.A(n1325));
   MUX2_X1 U403 (.Z(n1325), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1326));
   NAND2_X1 U404 (.ZN(n1326), 
	.A2(n1150), 
	.A1(n1327));
   NAND2_X1 U405 (.ZN(n1323), 
	.A2(n1320), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U406 (.Z(n1321), 
	.S(n1143), 
	.B(n1329), 
	.A(n1328));
   NAND2_X1 U407 (.ZN(n1329), 
	.A2(n1154), 
	.A1(n1298));
   NAND2_X1 U408 (.ZN(n1328), 
	.A2(n1154), 
	.A1(n1330));
   NAND2_X1 U409 (.ZN(B[23]), 
	.A2(n1332), 
	.A1(n1331));
   MUX2_X1 U410 (.Z(n1332), 
	.S(n1143), 
	.B(n1334), 
	.A(n1333));
   NAND2_X1 U411 (.ZN(n1334), 
	.A2(n1298), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U412 (.ZN(n1298), 
	.A2(n1336), 
	.A1(n1335));
   NAND3_X1 U413 (.ZN(n1336), 
	.A3(n1337), 
	.A2(n1113), 
	.A1(n1152));
   MUX2_X1 U414 (.Z(n1335), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1338));
   NAND2_X1 U415 (.ZN(n1338), 
	.A2(n1317), 
	.A1(n1146));
   NAND2_X1 U416 (.ZN(n1333), 
	.A2(n1330), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U417 (.Z(n1331), 
	.S(n1142), 
	.B(n1340), 
	.A(n1339));
   NAND2_X1 U418 (.ZN(n1340), 
	.A2(n1154), 
	.A1(n1302));
   NAND2_X1 U419 (.ZN(n1339), 
	.A2(n1154), 
	.A1(n1341));
   NAND2_X1 U420 (.ZN(B[22]), 
	.A2(n1343), 
	.A1(n1342));
   MUX2_X1 U421 (.Z(n1343), 
	.S(n1142), 
	.B(n1345), 
	.A(n1344));
   NAND2_X1 U422 (.ZN(n1345), 
	.A2(n1302), 
	.A1(SH[0]));
   NAND2_X1 U423 (.ZN(n1302), 
	.A2(n1347), 
	.A1(n1346));
   NAND3_X1 U424 (.ZN(n1347), 
	.A3(n1348), 
	.A2(n1112), 
	.A1(n1152));
   MUX2_X1 U425 (.Z(n1346), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1349));
   NAND2_X1 U426 (.ZN(n1349), 
	.A2(n1327), 
	.A1(n1146));
   NAND2_X1 U427 (.ZN(n1344), 
	.A2(n1341), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U428 (.Z(n1342), 
	.S(n1142), 
	.B(n1308), 
	.A(n1350));
   NAND2_X1 U430 (.ZN(n1350), 
	.A2(n1155), 
	.A1(n1352));
   NAND2_X1 U431 (.ZN(B[21]), 
	.A2(n1354), 
	.A1(n1353));
   MUX2_X1 U432 (.Z(n1354), 
	.S(n1142), 
	.B(n1356), 
	.A(n1355));
   NAND2_X1 U433 (.ZN(n1356), 
	.A2(n1310), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U434 (.ZN(n1310), 
	.A2(n1358), 
	.A1(n1357));
   NAND3_X1 U435 (.ZN(n1358), 
	.A3(n1359), 
	.A2(n1113), 
	.A1(n1152));
   MUX2_X1 U436 (.Z(n1357), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1360));
   NAND2_X1 U437 (.ZN(n1360), 
	.A2(n1337), 
	.A1(n1146));
   NAND2_X1 U438 (.ZN(n1355), 
	.A2(n1352), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U439 (.Z(n1353), 
	.S(n1142), 
	.B(n1362), 
	.A(n1361));
   NAND2_X1 U440 (.ZN(n1362), 
	.A2(n1155), 
	.A1(n1320));
   NAND2_X1 U441 (.ZN(n1361), 
	.A2(n1155), 
	.A1(n1363));
   NAND2_X1 U442 (.ZN(B[20]), 
	.A2(n1365), 
	.A1(n1364));
   MUX2_X1 U443 (.Z(n1365), 
	.S(n1142), 
	.B(n1367), 
	.A(n1366));
   NAND2_X1 U444 (.ZN(n1367), 
	.A2(n1320), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   NAND2_X1 U445 (.ZN(n1320), 
	.A2(n1369), 
	.A1(n1368));
   NAND3_X1 U446 (.ZN(n1369), 
	.A3(n1370), 
	.A2(n1112), 
	.A1(n1152));
   MUX2_X1 U447 (.Z(n1368), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1371));
   NAND2_X1 U448 (.ZN(n1371), 
	.A2(n1348), 
	.A1(n1146));
   NAND2_X1 U449 (.ZN(n1366), 
	.A2(n1363), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U450 (.Z(n1364), 
	.S(n1142), 
	.B(n1373), 
	.A(n1372));
   NAND2_X1 U451 (.ZN(n1373), 
	.A2(n1155), 
	.A1(n1330));
   NAND2_X1 U452 (.ZN(n1372), 
	.A2(n1155), 
	.A1(n1374));
   NAND2_X1 U453 (.ZN(B[1]), 
	.A2(n1376), 
	.A1(n1375));
   MUX2_X1 U454 (.Z(n1376), 
	.S(n1142), 
	.B(n1378), 
	.A(n1377));
   NAND2_X1 U455 (.ZN(n1378), 
	.A2(n1221), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U456 (.ZN(n1221), 
	.A2(n1380), 
	.A1(n1379));
   MUX2_X1 U457 (.Z(n1380), 
	.S(n1148), 
	.B(n1382), 
	.A(n1381));
   NAND2_X1 U458 (.ZN(n1382), 
	.A2(n1255), 
	.A1(SH[3]));
   NAND2_X1 U459 (.ZN(n1381), 
	.A2(n1383), 
	.A1(SH[3]));
   MUX2_X1 U460 (.Z(n1379), 
	.S(n1148), 
	.B(n1256), 
	.A(n1384));
   NAND2_X1 U462 (.ZN(n1384), 
	.A2(n1109), 
	.A1(n1386));
   NAND2_X1 U463 (.ZN(n1377), 
	.A2(n1291), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U464 (.ZN(n1291), 
	.A2(n1388), 
	.A1(n1387));
   MUX2_X1 U465 (.Z(n1388), 
	.S(n1148), 
	.B(n1390), 
	.A(n1389));
   NAND2_X1 U466 (.ZN(n1390), 
	.A2(n1391), 
	.A1(SH[3]));
   NAND2_X1 U467 (.ZN(n1389), 
	.A2(n1258), 
	.A1(SH[3]));
   MUX2_X1 U468 (.Z(n1387), 
	.S(n1148), 
	.B(n1393), 
	.A(n1392));
   NAND2_X1 U469 (.ZN(n1393), 
	.A2(n1109), 
	.A1(n1394));
   NAND2_X1 U470 (.ZN(n1392), 
	.A2(n1109), 
	.A1(n1395));
   MUX2_X1 U471 (.Z(n1375), 
	.S(n1142), 
	.B(n1397), 
	.A(n1396));
   NAND2_X1 U472 (.ZN(n1397), 
	.A2(n1155), 
	.A1(n1228));
   NAND2_X1 U473 (.ZN(n1396), 
	.A2(n1155), 
	.A1(n1398));
   NAND2_X1 U474 (.ZN(B[19]), 
	.A2(n1400), 
	.A1(n1399));
   MUX2_X1 U475 (.Z(n1400), 
	.S(n1142), 
	.B(n1402), 
	.A(n1401));
   NAND2_X1 U476 (.ZN(n1402), 
	.A2(n1330), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U477 (.ZN(n1330), 
	.A2(n1404), 
	.A1(n1403));
   NAND3_X1 U478 (.ZN(n1404), 
	.A3(n1405), 
	.A2(n1112), 
	.A1(n1152));
   MUX2_X1 U479 (.Z(n1403), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1406));
   NAND2_X1 U480 (.ZN(n1406), 
	.A2(n1359), 
	.A1(n1146));
   NAND2_X1 U481 (.ZN(n1401), 
	.A2(n1374), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   MUX2_X1 U482 (.Z(n1399), 
	.S(n1142), 
	.B(n1408), 
	.A(n1407));
   NAND2_X1 U483 (.ZN(n1408), 
	.A2(n1155), 
	.A1(n1341));
   NAND2_X1 U484 (.ZN(n1407), 
	.A2(n1155), 
	.A1(n1409));
   NAND2_X1 U485 (.ZN(B[18]), 
	.A2(n1411), 
	.A1(n1410));
   MUX2_X1 U486 (.Z(n1411), 
	.S(n1142), 
	.B(n1413), 
	.A(n1412));
   NAND2_X1 U487 (.ZN(n1413), 
	.A2(n1341), 
	.A1(SH[0]));
   NAND2_X1 U488 (.ZN(n1341), 
	.A2(n1415), 
	.A1(n1414));
   NAND3_X1 U489 (.ZN(n1415), 
	.A3(n1416), 
	.A2(n1112), 
	.A1(n1152));
   MUX2_X1 U490 (.Z(n1414), 
	.S(SH[3]), 
	.B(n1266), 
	.A(n1417));
   NAND2_X1 U491 (.ZN(n1417), 
	.A2(n1370), 
	.A1(n1146));
   NAND2_X1 U492 (.ZN(n1412), 
	.A2(n1409), 
	.A1(SH[0]));
   MUX2_X1 U493 (.Z(n1410), 
	.S(n1142), 
	.B(n1350), 
	.A(n1418));
   NAND2_X1 U495 (.ZN(n1418), 
	.A2(n1155), 
	.A1(n1420));
   NAND2_X1 U496 (.ZN(B[17]), 
	.A2(n1422), 
	.A1(n1421));
   MUX2_X1 U497 (.Z(n1422), 
	.S(n1142), 
	.B(n1424), 
	.A(n1423));
   NAND2_X1 U498 (.ZN(n1424), 
	.A2(n1352), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   NAND2_X1 U499 (.ZN(n1352), 
	.A2(n1426), 
	.A1(n1425));
   MUX2_X1 U500 (.Z(n1426), 
	.S(n1148), 
	.B(n1428), 
	.A(n1427));
   NAND2_X1 U501 (.ZN(n1428), 
	.A2(\A[31] ), 
	.A1(SH[3]));
   NAND2_X1 U502 (.ZN(n1427), 
	.A2(n1317), 
	.A1(SH[3]));
   MUX2_X1 U503 (.Z(n1425), 
	.S(n1148), 
	.B(n1430), 
	.A(n1429));
   NAND2_X1 U504 (.ZN(n1430), 
	.A2(n1109), 
	.A1(n1405));
   NAND2_X1 U505 (.ZN(n1429), 
	.A2(n1110), 
	.A1(n1431));
   NAND2_X1 U506 (.ZN(n1423), 
	.A2(n1420), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U507 (.Z(n1421), 
	.S(n1142), 
	.B(n1433), 
	.A(n1432));
   NAND2_X1 U508 (.ZN(n1433), 
	.A2(n1156), 
	.A1(n1363));
   NAND2_X1 U509 (.ZN(n1432), 
	.A2(n1156), 
	.A1(n1434));
   NAND2_X1 U510 (.ZN(B[16]), 
	.A2(n1436), 
	.A1(n1435));
   MUX2_X1 U511 (.Z(n1436), 
	.S(n1142), 
	.B(n1366), 
	.A(n1437));
   NAND2_X1 U513 (.ZN(n1363), 
	.A2(n1440), 
	.A1(n1439));
   MUX2_X1 U514 (.Z(n1440), 
	.S(n1148), 
	.B(n1442), 
	.A(n1441));
   NAND2_X1 U515 (.ZN(n1442), 
	.A2(\A[31] ), 
	.A1(SH[3]));
   NAND2_X1 U516 (.ZN(n1441), 
	.A2(n1327), 
	.A1(SH[3]));
   MUX2_X1 U517 (.Z(n1439), 
	.S(n1148), 
	.B(n1444), 
	.A(n1443));
   NAND2_X1 U518 (.ZN(n1444), 
	.A2(n1110), 
	.A1(n1416));
   NAND2_X1 U519 (.ZN(n1443), 
	.A2(n1110), 
	.A1(n1445));
   NAND2_X1 U520 (.ZN(n1437), 
	.A2(n1434), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U521 (.Z(n1435), 
	.S(n1141), 
	.B(n1447), 
	.A(n1446));
   NAND2_X1 U522 (.ZN(n1447), 
	.A2(n1156), 
	.A1(n1374));
   NAND2_X1 U523 (.ZN(n1446), 
	.A2(n1156), 
	.A1(n1448));
   NAND2_X1 U524 (.ZN(B[15]), 
	.A2(n1450), 
	.A1(n1449));
   MUX2_X1 U525 (.Z(n1450), 
	.S(n1141), 
	.B(n1452), 
	.A(n1451));
   NAND2_X1 U526 (.ZN(n1452), 
	.A2(n1374), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   NAND2_X1 U527 (.ZN(n1374), 
	.A2(n1454), 
	.A1(n1453));
   MUX2_X1 U528 (.Z(n1454), 
	.S(n1148), 
	.B(n1456), 
	.A(n1455));
   NAND2_X1 U529 (.ZN(n1456), 
	.A2(n1317), 
	.A1(SH[3]));
   INV_X1 U530 (.ZN(n1317), 
	.A(n1457));
   MUX2_X1 U531 (.Z(n1457), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1458));
   NAND2_X1 U532 (.ZN(n1455), 
	.A2(n1337), 
	.A1(SH[3]));
   MUX2_X1 U533 (.Z(n1453), 
	.S(n1148), 
	.B(n1429), 
	.A(n1459));
   NAND2_X1 U535 (.ZN(n1459), 
	.A2(n1110), 
	.A1(n1461));
   NAND2_X1 U536 (.ZN(n1451), 
	.A2(n1448), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U537 (.Z(n1449), 
	.S(n1141), 
	.B(n1463), 
	.A(n1462));
   NAND2_X1 U538 (.ZN(n1463), 
	.A2(n1156), 
	.A1(n1409));
   NAND2_X1 U539 (.ZN(n1462), 
	.A2(n1156), 
	.A1(n1464));
   NAND2_X1 U540 (.ZN(B[14]), 
	.A2(n1466), 
	.A1(n1465));
   MUX2_X1 U541 (.Z(n1466), 
	.S(n1141), 
	.B(n1468), 
	.A(n1467));
   NAND2_X1 U542 (.ZN(n1468), 
	.A2(n1409), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   NAND2_X1 U543 (.ZN(n1409), 
	.A2(n1470), 
	.A1(n1469));
   MUX2_X1 U544 (.Z(n1470), 
	.S(n1148), 
	.B(n1472), 
	.A(n1471));
   NAND2_X1 U545 (.ZN(n1472), 
	.A2(n1327), 
	.A1(SH[3]));
   INV_X1 U546 (.ZN(n1327), 
	.A(n1473));
   MUX2_X1 U547 (.Z(n1473), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1474));
   NAND2_X1 U548 (.ZN(n1471), 
	.A2(n1348), 
	.A1(SH[3]));
   MUX2_X1 U549 (.Z(n1469), 
	.S(n1148), 
	.B(n1443), 
	.A(n1475));
   NAND2_X1 U551 (.ZN(n1475), 
	.A2(n1110), 
	.A1(n1237));
   NAND2_X1 U552 (.ZN(n1467), 
	.A2(n1464), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U553 (.Z(n1465), 
	.S(n1141), 
	.B(n1478), 
	.A(n1477));
   NAND2_X1 U554 (.ZN(n1478), 
	.A2(n1156), 
	.A1(n1420));
   NAND2_X1 U555 (.ZN(n1477), 
	.A2(n1156), 
	.A1(n1193));
   NAND2_X1 U556 (.ZN(B[13]), 
	.A2(n1480), 
	.A1(n1479));
   MUX2_X1 U557 (.Z(n1480), 
	.S(n1141), 
	.B(n1423), 
	.A(n1481));
   NAND2_X1 U559 (.ZN(n1420), 
	.A2(n1484), 
	.A1(n1483));
   MUX2_X1 U560 (.Z(n1484), 
	.S(n1148), 
	.B(n1486), 
	.A(n1485));
   NAND2_X1 U561 (.ZN(n1486), 
	.A2(n1337), 
	.A1(SH[3]));
   INV_X1 U562 (.ZN(n1337), 
	.A(n1487));
   MUX2_X1 U563 (.Z(n1487), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1488));
   NAND2_X1 U564 (.ZN(n1485), 
	.A2(n1359), 
	.A1(SH[3]));
   MUX2_X1 U565 (.Z(n1483), 
	.S(n1148), 
	.B(n1459), 
	.A(n1489));
   NAND2_X1 U567 (.ZN(n1489), 
	.A2(n1110), 
	.A1(n1254));
   NAND2_X1 U568 (.ZN(n1481), 
	.A2(n1193), 
	.A1(FE_OFN183_UUT_Mpath_out_regB_0_));
   MUX2_X1 U569 (.Z(n1479), 
	.S(n1141), 
	.B(n1432), 
	.A(n1491));
   NAND2_X1 U571 (.ZN(n1491), 
	.A2(n1156), 
	.A1(n1197));
   NAND2_X1 U572 (.ZN(B[12]), 
	.A2(n1494), 
	.A1(n1493));
   MUX2_X1 U573 (.Z(n1494), 
	.S(n1141), 
	.B(n1496), 
	.A(n1495));
   NAND2_X1 U574 (.ZN(n1496), 
	.A2(n1434), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U575 (.ZN(n1434), 
	.A2(n1498), 
	.A1(n1497));
   MUX2_X1 U576 (.Z(n1498), 
	.S(n1147), 
	.B(n1500), 
	.A(n1499));
   NAND2_X1 U577 (.ZN(n1500), 
	.A2(n1348), 
	.A1(SH[3]));
   INV_X1 U578 (.ZN(n1348), 
	.A(n1501));
   MUX2_X1 U579 (.Z(n1501), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1502));
   NAND2_X1 U580 (.ZN(n1499), 
	.A2(n1370), 
	.A1(SH[3]));
   MUX2_X1 U581 (.Z(n1497), 
	.S(n1147), 
	.B(n1475), 
	.A(n1503));
   NAND2_X1 U583 (.ZN(n1503), 
	.A2(n1110), 
	.A1(n1238));
   NAND2_X1 U584 (.ZN(n1495), 
	.A2(n1197), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U585 (.ZN(n1197), 
	.A2(n1506), 
	.A1(n1505));
   MUX2_X1 U586 (.Z(n1506), 
	.S(n1147), 
	.B(n1508), 
	.A(n1507));
   NAND2_X1 U587 (.ZN(n1508), 
	.A2(n1416), 
	.A1(SH[3]));
   NAND2_X1 U588 (.ZN(n1507), 
	.A2(n1445), 
	.A1(SH[3]));
   MUX2_X1 U589 (.Z(n1505), 
	.S(n1147), 
	.B(n1510), 
	.A(n1509));
   NAND2_X1 U590 (.ZN(n1510), 
	.A2(n1111), 
	.A1(n1276));
   NAND2_X1 U591 (.ZN(n1509), 
	.A2(n1111), 
	.A1(n1284));
   MUX2_X1 U592 (.Z(n1493), 
	.S(n1141), 
	.B(n1512), 
	.A(n1511));
   NAND2_X1 U593 (.ZN(n1512), 
	.A2(n1157), 
	.A1(n1448));
   NAND2_X1 U594 (.ZN(n1511), 
	.A2(n1156), 
	.A1(n1205));
   NAND2_X1 U595 (.ZN(B[11]), 
	.A2(n1514), 
	.A1(n1513));
   MUX2_X1 U596 (.Z(n1514), 
	.S(n1141), 
	.B(n1516), 
	.A(n1515));
   NAND2_X1 U597 (.ZN(n1516), 
	.A2(n1448), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U598 (.ZN(n1448), 
	.A2(n1518), 
	.A1(n1517));
   MUX2_X1 U599 (.Z(n1518), 
	.S(n1147), 
	.B(n1520), 
	.A(n1519));
   NAND2_X1 U600 (.ZN(n1520), 
	.A2(n1359), 
	.A1(SH[3]));
   INV_X1 U601 (.ZN(n1359), 
	.A(n1521));
   MUX2_X1 U602 (.Z(n1521), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1522));
   NAND2_X1 U603 (.ZN(n1519), 
	.A2(n1405), 
	.A1(SH[3]));
   MUX2_X1 U604 (.Z(n1517), 
	.S(n1147), 
	.B(n1524), 
	.A(n1523));
   NAND2_X1 U605 (.ZN(n1524), 
	.A2(n1111), 
	.A1(n1254));
   NAND2_X1 U606 (.ZN(n1523), 
	.A2(n1111), 
	.A1(n1255));
   NAND2_X1 U607 (.ZN(n1515), 
	.A2(n1205), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U608 (.ZN(n1205), 
	.A2(n1526), 
	.A1(n1525));
   MUX2_X1 U609 (.Z(n1526), 
	.S(n1147), 
	.B(n1528), 
	.A(n1527));
   NAND2_X1 U610 (.ZN(n1528), 
	.A2(n1431), 
	.A1(SH[3]));
   NAND2_X1 U611 (.ZN(n1527), 
	.A2(n1461), 
	.A1(SH[3]));
   MUX2_X1 U612 (.Z(n1525), 
	.S(n1147), 
	.B(n1530), 
	.A(n1529));
   NAND2_X1 U613 (.ZN(n1530), 
	.A2(n1111), 
	.A1(n1383));
   NAND2_X1 U614 (.ZN(n1529), 
	.A2(n1111), 
	.A1(n1391));
   MUX2_X1 U615 (.Z(n1513), 
	.S(n1141), 
	.B(n1532), 
	.A(n1531));
   NAND2_X1 U616 (.ZN(n1532), 
	.A2(n1157), 
	.A1(n1464));
   NAND2_X1 U617 (.ZN(n1531), 
	.A2(n1156), 
	.A1(n1213));
   NAND2_X1 U618 (.ZN(B[10]), 
	.A2(n1534), 
	.A1(n1533));
   MUX2_X1 U619 (.Z(n1534), 
	.S(n1141), 
	.B(n1536), 
	.A(n1535));
   NAND2_X1 U620 (.ZN(n1536), 
	.A2(n1464), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U621 (.ZN(n1464), 
	.A2(n1538), 
	.A1(n1537));
   MUX2_X1 U622 (.Z(n1538), 
	.S(n1147), 
	.B(n1540), 
	.A(n1539));
   NAND2_X1 U623 (.ZN(n1540), 
	.A2(n1370), 
	.A1(SH[3]));
   INV_X1 U624 (.ZN(n1370), 
	.A(n1541));
   MUX2_X1 U625 (.Z(n1541), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1542));
   NAND2_X1 U626 (.ZN(n1539), 
	.A2(n1416), 
	.A1(SH[3]));
   INV_X1 U627 (.ZN(n1416), 
	.A(n1543));
   MUX2_X1 U628 (.Z(n1543), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1544));
   MUX2_X1 U629 (.Z(n1537), 
	.S(n1147), 
	.B(n1546), 
	.A(n1510));
   NAND2_X1 U630 (.ZN(n1546), 
	.A2(n1111), 
	.A1(n1238));
   INV_X1 U631 (.ZN(n1238), 
	.A(n1547));
   MUX2_X1 U632 (.Z(n1547), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1548));
   NAND2_X1 U634 (.ZN(n1535), 
	.A2(n1213), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U635 (.ZN(n1213), 
	.A2(n1550), 
	.A1(n1549));
   MUX2_X1 U636 (.Z(n1550), 
	.S(n1147), 
	.B(n1552), 
	.A(n1551));
   NAND2_X1 U637 (.ZN(n1552), 
	.A2(n1445), 
	.A1(SH[3]));
   INV_X1 U638 (.ZN(n1445), 
	.A(n1553));
   MUX2_X1 U639 (.Z(n1553), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1554));
   NAND2_X1 U640 (.ZN(n1551), 
	.A2(n1237), 
	.A1(SH[3]));
   INV_X1 U641 (.ZN(n1237), 
	.A(n1555));
   MUX2_X1 U642 (.Z(n1555), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1556));
   MUX2_X1 U643 (.Z(n1549), 
	.S(n1147), 
	.B(n1509), 
	.A(n1557));
   NAND2_X1 U645 (.ZN(n1557), 
	.A2(n1111), 
	.A1(n1241));
   MUX2_X1 U646 (.Z(n1533), 
	.S(n1141), 
	.B(n1560), 
	.A(n1559));
   NAND2_X1 U647 (.ZN(n1560), 
	.A2(n1157), 
	.A1(n1193));
   NAND2_X1 U648 (.ZN(n1193), 
	.A2(n1562), 
	.A1(n1561));
   MUX2_X1 U649 (.Z(n1562), 
	.S(n1147), 
	.B(n1564), 
	.A(n1563));
   NAND2_X1 U650 (.ZN(n1564), 
	.A2(n1405), 
	.A1(SH[3]));
   INV_X1 U651 (.ZN(n1405), 
	.A(n1565));
   MUX2_X1 U652 (.Z(n1565), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1566));
   NAND2_X1 U653 (.ZN(n1563), 
	.A2(n1431), 
	.A1(SH[3]));
   INV_X1 U654 (.ZN(n1431), 
	.A(n1567));
   MUX2_X1 U655 (.Z(n1567), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1568));
   MUX2_X1 U656 (.Z(n1561), 
	.S(n1147), 
	.B(n1523), 
	.A(n1530));
   INV_X1 U658 (.ZN(n1255), 
	.A(n1571));
   MUX2_X1 U659 (.Z(n1571), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1572));
   NAND2_X1 U661 (.ZN(n1559), 
	.A2(n1157), 
	.A1(n1194));
   NAND2_X1 U662 (.ZN(n1194), 
	.A2(n1574), 
	.A1(n1573));
   MUX2_X1 U663 (.Z(n1574), 
	.S(n1147), 
	.B(n1576), 
	.A(n1575));
   NAND2_X1 U664 (.ZN(n1576), 
	.A2(n1461), 
	.A1(SH[3]));
   INV_X1 U665 (.ZN(n1461), 
	.A(n1577));
   MUX2_X1 U666 (.Z(n1577), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1578));
   NAND2_X1 U667 (.ZN(n1575), 
	.A2(n1254), 
	.A1(SH[3]));
   INV_X1 U668 (.ZN(n1254), 
	.A(n1579));
   MUX2_X1 U669 (.Z(n1579), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1580));
   MUX2_X1 U670 (.Z(n1573), 
	.S(n1146), 
	.B(n1582), 
	.A(n1581));
   NAND2_X1 U671 (.ZN(n1582), 
	.A2(n1112), 
	.A1(n1391));
   NAND2_X1 U672 (.ZN(n1581), 
	.A2(n1112), 
	.A1(n1258));
   NAND2_X1 U673 (.ZN(B[0]), 
	.A2(n1584), 
	.A1(n1583));
   MUX2_X1 U674 (.Z(n1584), 
	.S(n1141), 
	.B(n1586), 
	.A(n1585));
   NAND2_X1 U675 (.ZN(n1586), 
	.A2(n1228), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U676 (.ZN(n1228), 
	.A2(n1588), 
	.A1(n1587));
   MUX2_X1 U677 (.Z(n1588), 
	.S(n1146), 
	.B(n1590), 
	.A(n1589));
   NAND2_X1 U678 (.ZN(n1590), 
	.A2(n1276), 
	.A1(SH[3]));
   INV_X1 U679 (.ZN(n1276), 
	.A(n1591));
   MUX2_X1 U680 (.Z(n1591), 
	.S(SH[4]), 
	.B(n1266), 
	.A(n1592));
   INV_X1 U681 (.ZN(n1266), 
	.A(\A[31] ));
   NAND2_X1 U682 (.ZN(n1589), 
	.A2(n1284), 
	.A1(SH[3]));
   INV_X1 U683 (.ZN(n1284), 
	.A(n1593));
   MUX2_X1 U684 (.Z(n1593), 
	.S(SH[4]), 
	.B(n1474), 
	.A(n1594));
   MUX2_X1 U685 (.Z(n1587), 
	.S(n1146), 
	.B(n1596), 
	.A(n1595));
   NAND2_X1 U686 (.ZN(n1596), 
	.A2(n1112), 
	.A1(n1279));
   INV_X1 U687 (.ZN(n1279), 
	.A(n1597));
   MUX2_X1 U688 (.Z(n1597), 
	.S(SH[4]), 
	.B(n1544), 
	.A(n1598));
   NAND2_X1 U689 (.ZN(n1595), 
	.A2(n1112), 
	.A1(n1287));
   INV_X1 U690 (.ZN(n1287), 
	.A(n1599));
   MUX2_X1 U691 (.Z(n1599), 
	.S(SH[4]), 
	.B(n1554), 
	.A(n1600));
   NAND2_X1 U692 (.ZN(n1585), 
	.A2(n1398), 
	.A1(FE_OFN180_UUT_Mpath_out_regB_0_));
   NAND2_X1 U693 (.ZN(n1398), 
	.A2(n1602), 
	.A1(n1601));
   MUX2_X1 U694 (.Z(n1602), 
	.S(n1146), 
	.B(n1604), 
	.A(n1603));
   NAND2_X1 U695 (.ZN(n1604), 
	.A2(n1241), 
	.A1(FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_));
   INV_X1 U696 (.ZN(n1241), 
	.A(n1605));
   MUX2_X1 U697 (.Z(n1605), 
	.S(SH[4]), 
	.B(n1502), 
	.A(n1606));
   NAND2_X1 U698 (.ZN(n1603), 
	.A2(n1242), 
	.A1(SH[3]));
   INV_X1 U699 (.ZN(n1242), 
	.A(n1607));
   MUX2_X1 U700 (.Z(n1607), 
	.S(SH[4]), 
	.B(n1542), 
	.A(n1608));
   MUX2_X1 U701 (.Z(n1601), 
	.S(n1147), 
	.B(n1610), 
	.A(n1609));
   NAND2_X1 U702 (.ZN(n1610), 
	.A2(n1112), 
	.A1(n1288));
   INV_X1 U703 (.ZN(n1288), 
	.A(n1611));
   MUX2_X1 U704 (.Z(n1611), 
	.S(FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(n1556), 
	.A(n1612));
   NAND2_X1 U705 (.ZN(n1609), 
	.A2(n1112), 
	.A1(n1613));
   MUX2_X1 U706 (.Z(n1613), 
	.S(FE_OFN160_UUT_Mpath_out_regB_4_), 
	.B(A[17]), 
	.A(A[1]));
   MUX2_X1 U707 (.Z(n1583), 
	.S(n1142), 
	.B(n1615), 
	.A(n1614));
   NAND2_X1 U708 (.ZN(n1615), 
	.A2(n1157), 
	.A1(n1245));
   NAND2_X1 U709 (.ZN(n1245), 
	.A2(n1617), 
	.A1(n1616));
   MUX2_X1 U710 (.Z(n1617), 
	.S(n1146), 
	.B(n1619), 
	.A(n1618));
   NAND2_X1 U711 (.ZN(n1619), 
	.A2(n1383), 
	.A1(SH[3]));
   INV_X1 U712 (.ZN(n1383), 
	.A(n1620));
   MUX2_X1 U713 (.Z(n1620), 
	.S(SH[4]), 
	.B(n1458), 
	.A(n1621));
   NAND2_X1 U714 (.ZN(n1618), 
	.A2(n1391), 
	.A1(SH[3]));
   INV_X1 U715 (.ZN(n1391), 
	.A(n1622));
   MUX2_X1 U716 (.Z(n1622), 
	.S(SH[4]), 
	.B(n1488), 
	.A(n1623));
   MUX2_X1 U717 (.Z(n1616), 
	.S(n1146), 
	.B(n1625), 
	.A(n1624));
   NAND2_X1 U718 (.ZN(n1625), 
	.A2(n1112), 
	.A1(n1386));
   INV_X1 U719 (.ZN(n1386), 
	.A(n1626));
   MUX2_X1 U720 (.Z(n1626), 
	.S(SH[4]), 
	.B(n1568), 
	.A(n1627));
   NAND2_X1 U721 (.ZN(n1624), 
	.A2(n1112), 
	.A1(n1394));
   INV_X1 U722 (.ZN(n1394), 
	.A(n1628));
   MUX2_X1 U723 (.Z(n1628), 
	.S(SH[4]), 
	.B(n1578), 
	.A(n1629));
   OAI21_X1 U724 (.ZN(n1614), 
	.B2(n1631), 
	.B1(n1630), 
	.A(n1157));
   MUX2_X1 U725 (.Z(n1631), 
	.S(n1146), 
	.B(n1633), 
	.A(n1632));
   AND2_X1 U726 (.ZN(n1633), 
	.A2(n1112), 
	.A1(n1395));
   INV_X1 U727 (.ZN(n1395), 
	.A(n1634));
   MUX2_X1 U728 (.Z(n1634), 
	.S(SH[4]), 
	.B(n1580), 
	.A(n1635));
   AND2_X1 U729 (.ZN(n1632), 
	.A2(n1112), 
	.A1(n1636));
   MUX2_X1 U730 (.Z(n1636), 
	.S(SH[4]), 
	.B(A[16]), 
	.A(A[0]));
   MUX2_X1 U731 (.Z(n1630), 
	.S(n1147), 
	.B(n1638), 
	.A(n1637));
   AND2_X1 U732 (.ZN(n1638), 
	.A2(n1258), 
	.A1(SH[3]));
   INV_X1 U733 (.ZN(n1258), 
	.A(n1639));
   MUX2_X1 U734 (.Z(n1639), 
	.S(SH[4]), 
	.B(n1522), 
	.A(n1640));
   AND2_X1 U735 (.ZN(n1637), 
	.A2(n1259), 
	.A1(SH[3]));
   INV_X1 U736 (.ZN(n1259), 
	.A(n1641));
   MUX2_X1 U737 (.Z(n1641), 
	.S(SH[4]), 
	.B(n1566), 
	.A(n1642));
endmodule

module up_island_DW_rightsh_1 (
	A, 
	SH, 
	B, 
	DATA_TC, 
	FE_OFN169_UUT_Mpath_out_regB_2_, 
	FE_OFN175_UUT_Mpath_out_regB_1_, 
	FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_);
   input [31:0] A;
   input [4:0] SH;
   output [31:0] B;
   input DATA_TC;
   input FE_OFN169_UUT_Mpath_out_regB_2_;
   input FE_OFN175_UUT_Mpath_out_regB_1_;
   input FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_;

   // Internal wires
   wire n378;
   wire n379;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n392;
   wire n394;
   wire n395;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;

   INV_X1 U174 (.ZN(n585), 
	.A(A[18]));
   INV_X1 U175 (.ZN(n572), 
	.A(A[15]));
   INV_X1 U176 (.ZN(n583), 
	.A(A[19]));
   INV_X1 U177 (.ZN(n581), 
	.A(A[20]));
   INV_X1 U178 (.ZN(n579), 
	.A(A[21]));
   INV_X1 U179 (.ZN(n438), 
	.A(A[9]));
   INV_X1 U180 (.ZN(n584), 
	.A(A[10]));
   INV_X1 U181 (.ZN(n575), 
	.A(A[22]));
   INV_X1 U182 (.ZN(n573), 
	.A(A[23]));
   INV_X1 U183 (.ZN(n486), 
	.A(A[8]));
   INV_X1 U184 (.ZN(n487), 
	.A(A[16]));
   INV_X1 U185 (.ZN(n439), 
	.A(A[17]));
   NAND2_X1 U186 (.ZN(n563), 
	.A2(n384), 
	.A1(A[28]));
   INV_X1 U187 (.ZN(n592), 
	.A(A[28]));
   NAND2_X1 U188 (.ZN(n562), 
	.A2(n385), 
	.A1(A[27]));
   INV_X1 U189 (.ZN(n599), 
	.A(A[27]));
   NAND2_X1 U190 (.ZN(n503), 
	.A2(n382), 
	.A1(A[25]));
   INV_X1 U191 (.ZN(n601), 
	.A(A[25]));
   NAND2_X1 U192 (.ZN(n561), 
	.A2(n383), 
	.A1(A[30]));
   INV_X1 U193 (.ZN(n590), 
	.A(A[30]));
   INV_X1 U194 (.ZN(n593), 
	.A(A[7]));
   INV_X1 U195 (.ZN(n574), 
	.A(A[14]));
   INV_X1 U196 (.ZN(n578), 
	.A(A[13]));
   INV_X1 U197 (.ZN(n582), 
	.A(A[11]));
   INV_X1 U198 (.ZN(n580), 
	.A(A[12]));
   NAND2_X1 U199 (.ZN(n560), 
	.A2(n384), 
	.A1(A[29]));
   INV_X1 U200 (.ZN(n591), 
	.A(A[29]));
   INV_X1 U201 (.ZN(n595), 
	.A(A[5]));
   NAND2_X1 U202 (.ZN(n504), 
	.A2(n385), 
	.A1(A[26]));
   INV_X1 U203 (.ZN(n600), 
	.A(A[26]));
   NAND2_X1 U204 (.ZN(n509), 
	.A2(n382), 
	.A1(A[24]));
   INV_X1 U205 (.ZN(n602), 
	.A(A[24]));
   INV_X1 U206 (.ZN(n594), 
	.A(A[6]));
   INV_X1 U207 (.ZN(n596), 
	.A(A[4]));
   INV_X1 U208 (.ZN(n605), 
	.A(A[3]));
   INV_X1 U209 (.ZN(n606), 
	.A(A[2]));
   INV_X1 U210 (.ZN(n397), 
	.A(SH[0]));
   INV_X1 U211 (.ZN(n609), 
	.A(A[1]));
   INV_X1 U212 (.ZN(n378), 
	.A(SH[4]));
   INV_X1 U213 (.ZN(n379), 
	.A(SH[4]));
   INV_X1 U216 (.ZN(n382), 
	.A(SH[3]));
   INV_X1 U217 (.ZN(n383), 
	.A(SH[3]));
   INV_X1 U218 (.ZN(n384), 
	.A(SH[3]));
   INV_X1 U219 (.ZN(n385), 
	.A(SH[3]));
   INV_X1 U226 (.ZN(n392), 
	.A(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_));
   INV_X1 U228 (.ZN(n394), 
	.A(n397));
   INV_X1 U229 (.ZN(n395), 
	.A(n397));
   MUX2_X1 U231 (.Z(B[9]), 
	.S(SH[2]), 
	.B(n399), 
	.A(n398));
   MUX2_X1 U232 (.Z(B[8]), 
	.S(SH[2]), 
	.B(n401), 
	.A(n400));
   MUX2_X1 U233 (.Z(B[7]), 
	.S(SH[2]), 
	.B(n403), 
	.A(n402));
   MUX2_X1 U234 (.Z(B[6]), 
	.S(SH[2]), 
	.B(n405), 
	.A(n404));
   MUX2_X1 U235 (.Z(B[5]), 
	.S(SH[2]), 
	.B(n398), 
	.A(n406));
   INV_X1 U236 (.ZN(n398), 
	.A(n407));
   MUX2_X1 U237 (.Z(n407), 
	.S(SH[4]), 
	.B(n409), 
	.A(n408));
   MUX2_X1 U238 (.Z(n408), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n411), 
	.A(n410));
   MUX2_X1 U239 (.Z(B[4]), 
	.S(SH[2]), 
	.B(n400), 
	.A(n412));
   INV_X1 U240 (.ZN(n400), 
	.A(n413));
   MUX2_X1 U241 (.Z(n413), 
	.S(SH[4]), 
	.B(n415), 
	.A(n414));
   MUX2_X1 U242 (.Z(n414), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n417), 
	.A(n416));
   MUX2_X1 U243 (.Z(B[3]), 
	.S(SH[2]), 
	.B(n402), 
	.A(n418));
   INV_X1 U244 (.ZN(n402), 
	.A(n419));
   MUX2_X1 U245 (.Z(n419), 
	.S(SH[4]), 
	.B(n421), 
	.A(n420));
   MUX2_X1 U246 (.Z(n420), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n410), 
	.A(n422));
   MUX2_X1 U247 (.Z(n410), 
	.S(n394), 
	.B(n424), 
	.A(n423));
   MUX2_X1 U248 (.Z(n418), 
	.S(SH[4]), 
	.B(n426), 
	.A(n425));
   MUX2_X1 U249 (.Z(n425), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n428), 
	.A(n427));
   INV_X1 U250 (.ZN(n428), 
	.A(n429));
   NOR2_X1 U251 (.ZN(B[31]), 
	.A2(n430), 
	.A1(SH[2]));
   NOR2_X1 U252 (.ZN(B[30]), 
	.A2(n431), 
	.A1(SH[2]));
   MUX2_X1 U253 (.Z(B[2]), 
	.S(SH[2]), 
	.B(n404), 
	.A(n432));
   INV_X1 U254 (.ZN(n404), 
	.A(n433));
   MUX2_X1 U255 (.Z(n433), 
	.S(SH[4]), 
	.B(n435), 
	.A(n434));
   MUX2_X1 U256 (.Z(n434), 
	.S(SH[1]), 
	.B(n416), 
	.A(n436));
   MUX2_X1 U257 (.Z(n416), 
	.S(n394), 
	.B(n423), 
	.A(n437));
   MUX2_X1 U258 (.Z(n423), 
	.S(SH[3]), 
	.B(n439), 
	.A(n438));
   MUX2_X1 U259 (.Z(n432), 
	.S(SH[4]), 
	.B(n441), 
	.A(n440));
   MUX2_X1 U260 (.Z(n440), 
	.S(SH[1]), 
	.B(n443), 
	.A(n442));
   INV_X1 U261 (.ZN(n443), 
	.A(n444));
   NOR2_X1 U262 (.ZN(B[29]), 
	.A2(n445), 
	.A1(SH[2]));
   NOR2_X1 U263 (.ZN(B[28]), 
	.A2(n446), 
	.A1(FE_OFN169_UUT_Mpath_out_regB_2_));
   MUX2_X1 U264 (.Z(B[27]), 
	.S(SH[2]), 
	.B(n448), 
	.A(n447));
   INV_X1 U265 (.ZN(n448), 
	.A(n430));
   NAND2_X1 U266 (.ZN(n430), 
	.A2(n379), 
	.A1(n449));
   INV_X1 U267 (.ZN(n449), 
	.A(n450));
   MUX2_X1 U268 (.Z(B[26]), 
	.S(SH[2]), 
	.B(n452), 
	.A(n451));
   INV_X1 U269 (.ZN(n452), 
	.A(n431));
   NAND2_X1 U270 (.ZN(n431), 
	.A2(n379), 
	.A1(n453));
   INV_X1 U271 (.ZN(n453), 
	.A(n454));
   MUX2_X1 U272 (.Z(B[25]), 
	.S(FE_OFN169_UUT_Mpath_out_regB_2_), 
	.B(n456), 
	.A(n455));
   INV_X1 U273 (.ZN(n456), 
	.A(n445));
   NAND2_X1 U274 (.ZN(n445), 
	.A2(n379), 
	.A1(n457));
   INV_X1 U275 (.ZN(n457), 
	.A(n458));
   MUX2_X1 U276 (.Z(B[24]), 
	.S(SH[2]), 
	.B(n460), 
	.A(n459));
   INV_X1 U277 (.ZN(n460), 
	.A(n446));
   NAND2_X1 U278 (.ZN(n446), 
	.A2(n379), 
	.A1(n461));
   INV_X1 U279 (.ZN(n461), 
	.A(n462));
   MUX2_X1 U280 (.Z(B[23]), 
	.S(SH[2]), 
	.B(n447), 
	.A(n463));
   INV_X1 U281 (.ZN(n447), 
	.A(n464));
   NAND2_X1 U282 (.ZN(n464), 
	.A2(n378), 
	.A1(n465));
   INV_X1 U283 (.ZN(n465), 
	.A(n466));
   MUX2_X1 U284 (.Z(B[22]), 
	.S(SH[2]), 
	.B(n451), 
	.A(n467));
   INV_X1 U285 (.ZN(n451), 
	.A(n468));
   NAND2_X1 U286 (.ZN(n468), 
	.A2(n378), 
	.A1(n469));
   INV_X1 U287 (.ZN(n469), 
	.A(n470));
   MUX2_X1 U288 (.Z(B[21]), 
	.S(SH[2]), 
	.B(n455), 
	.A(n471));
   INV_X1 U289 (.ZN(n455), 
	.A(n472));
   NAND2_X1 U290 (.ZN(n472), 
	.A2(n378), 
	.A1(n473));
   INV_X1 U291 (.ZN(n473), 
	.A(n409));
   MUX2_X1 U292 (.Z(n409), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n475), 
	.A(n474));
   MUX2_X1 U293 (.Z(B[20]), 
	.S(SH[2]), 
	.B(n459), 
	.A(n476));
   INV_X1 U294 (.ZN(n459), 
	.A(n477));
   NAND2_X1 U295 (.ZN(n477), 
	.A2(n378), 
	.A1(n478));
   INV_X1 U296 (.ZN(n478), 
	.A(n415));
   MUX2_X1 U297 (.Z(n415), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n480), 
	.A(n479));
   MUX2_X1 U298 (.Z(B[1]), 
	.S(SH[2]), 
	.B(n406), 
	.A(n481));
   INV_X1 U299 (.ZN(n406), 
	.A(n482));
   MUX2_X1 U300 (.Z(n482), 
	.S(SH[4]), 
	.B(n484), 
	.A(n483));
   MUX2_X1 U301 (.Z(n483), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n422), 
	.A(n429));
   MUX2_X1 U302 (.Z(n422), 
	.S(n394), 
	.B(n437), 
	.A(n485));
   MUX2_X1 U303 (.Z(n437), 
	.S(SH[3]), 
	.B(n487), 
	.A(n486));
   MUX2_X1 U304 (.Z(n429), 
	.S(n394), 
	.B(n489), 
	.A(n488));
   MUX2_X1 U305 (.Z(n481), 
	.S(SH[4]), 
	.B(n491), 
	.A(n490));
   MUX2_X1 U306 (.Z(n490), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n427), 
	.A(n492));
   INV_X1 U307 (.ZN(n427), 
	.A(n493));
   MUX2_X1 U308 (.Z(n493), 
	.S(n394), 
	.B(n495), 
	.A(n494));
   MUX2_X1 U309 (.Z(n492), 
	.S(n394), 
	.B(n497), 
	.A(n496));
   INV_X1 U310 (.ZN(n497), 
	.A(n498));
   MUX2_X1 U311 (.Z(B[19]), 
	.S(SH[2]), 
	.B(n463), 
	.A(n499));
   INV_X1 U312 (.ZN(n463), 
	.A(n500));
   NAND2_X1 U313 (.ZN(n500), 
	.A2(n378), 
	.A1(n501));
   INV_X1 U314 (.ZN(n501), 
	.A(n421));
   MUX2_X1 U315 (.Z(n421), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n474), 
	.A(n502));
   MUX2_X1 U316 (.Z(n474), 
	.S(n394), 
	.B(n504), 
	.A(n503));
   MUX2_X1 U317 (.Z(B[18]), 
	.S(SH[2]), 
	.B(n467), 
	.A(n505));
   INV_X1 U318 (.ZN(n467), 
	.A(n506));
   NAND2_X1 U319 (.ZN(n506), 
	.A2(n378), 
	.A1(n507));
   INV_X1 U320 (.ZN(n507), 
	.A(n435));
   MUX2_X1 U321 (.Z(n435), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n479), 
	.A(n508));
   MUX2_X1 U322 (.Z(n479), 
	.S(n394), 
	.B(n503), 
	.A(n509));
   MUX2_X1 U323 (.Z(B[17]), 
	.S(SH[2]), 
	.B(n471), 
	.A(n510));
   INV_X1 U324 (.ZN(n471), 
	.A(n511));
   NAND2_X1 U325 (.ZN(n511), 
	.A2(n378), 
	.A1(n512));
   INV_X1 U326 (.ZN(n512), 
	.A(n484));
   MUX2_X1 U327 (.Z(n484), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n502), 
	.A(n513));
   MUX2_X1 U328 (.Z(n502), 
	.S(n394), 
	.B(n509), 
	.A(n514));
   MUX2_X1 U329 (.Z(B[16]), 
	.S(SH[2]), 
	.B(n476), 
	.A(n515));
   INV_X1 U330 (.ZN(n476), 
	.A(n516));
   NAND2_X1 U331 (.ZN(n516), 
	.A2(n378), 
	.A1(n517));
   INV_X1 U332 (.ZN(n517), 
	.A(n518));
   MUX2_X1 U333 (.Z(B[15]), 
	.S(SH[2]), 
	.B(n499), 
	.A(n519));
   INV_X1 U334 (.ZN(n499), 
	.A(n520));
   NAND2_X1 U335 (.ZN(n520), 
	.A2(n378), 
	.A1(n426));
   INV_X1 U336 (.ZN(n426), 
	.A(n521));
   MUX2_X1 U337 (.Z(n521), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n513), 
	.A(n522));
   MUX2_X1 U338 (.Z(n513), 
	.S(n394), 
	.B(n524), 
	.A(n523));
   MUX2_X1 U339 (.Z(B[14]), 
	.S(SH[2]), 
	.B(n505), 
	.A(n525));
   INV_X1 U340 (.ZN(n505), 
	.A(n526));
   NAND2_X1 U341 (.ZN(n526), 
	.A2(n378), 
	.A1(n441));
   INV_X1 U342 (.ZN(n441), 
	.A(n527));
   MUX2_X1 U343 (.Z(n527), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n529), 
	.A(n528));
   MUX2_X1 U344 (.Z(B[13]), 
	.S(SH[2]), 
	.B(n510), 
	.A(n399));
   INV_X1 U345 (.ZN(n510), 
	.A(n530));
   NAND2_X1 U346 (.ZN(n530), 
	.A2(n378), 
	.A1(n491));
   INV_X1 U347 (.ZN(n491), 
	.A(n531));
   MUX2_X1 U348 (.Z(n531), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n522), 
	.A(n532));
   MUX2_X1 U349 (.Z(n522), 
	.S(n394), 
	.B(n534), 
	.A(n533));
   INV_X1 U350 (.ZN(n399), 
	.A(n535));
   MUX2_X1 U351 (.Z(n535), 
	.S(SH[4]), 
	.B(n458), 
	.A(n536));
   MUX2_X1 U352 (.Z(n458), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n538), 
	.A(n537));
   MUX2_X1 U353 (.Z(n536), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n540), 
	.A(n539));
   MUX2_X1 U354 (.Z(B[12]), 
	.S(SH[2]), 
	.B(n515), 
	.A(n401));
   INV_X1 U355 (.ZN(n515), 
	.A(n541));
   NAND2_X1 U356 (.ZN(n541), 
	.A2(n378), 
	.A1(n542));
   INV_X1 U357 (.ZN(n401), 
	.A(n543));
   MUX2_X1 U358 (.Z(n543), 
	.S(SH[4]), 
	.B(n462), 
	.A(n544));
   MUX2_X1 U359 (.Z(n462), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n546), 
	.A(n545));
   MUX2_X1 U360 (.Z(n544), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n548), 
	.A(n547));
   MUX2_X1 U361 (.Z(B[11]), 
	.S(SH[2]), 
	.B(n519), 
	.A(n403));
   INV_X1 U362 (.ZN(n519), 
	.A(n549));
   MUX2_X1 U363 (.Z(n549), 
	.S(SH[4]), 
	.B(n450), 
	.A(n550));
   NAND2_X1 U364 (.ZN(n450), 
	.A2(n392), 
	.A1(n551));
   INV_X1 U365 (.ZN(n551), 
	.A(n538));
   NAND2_X1 U366 (.ZN(n538), 
	.A2(n397), 
	.A1(n552));
   INV_X1 U367 (.ZN(n552), 
	.A(n553));
   MUX2_X1 U368 (.Z(n550), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n532), 
	.A(n540));
   MUX2_X1 U369 (.Z(n532), 
	.S(n394), 
	.B(n555), 
	.A(n554));
   MUX2_X1 U370 (.Z(n540), 
	.S(n395), 
	.B(n557), 
	.A(n556));
   INV_X1 U371 (.ZN(n403), 
	.A(n558));
   MUX2_X1 U372 (.Z(n558), 
	.S(SH[4]), 
	.B(n466), 
	.A(n559));
   MUX2_X1 U373 (.Z(n466), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n537), 
	.A(n475));
   MUX2_X1 U374 (.Z(n537), 
	.S(n395), 
	.B(n561), 
	.A(n560));
   MUX2_X1 U375 (.Z(n475), 
	.S(n395), 
	.B(n563), 
	.A(n562));
   MUX2_X1 U376 (.Z(n559), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n539), 
	.A(n411));
   MUX2_X1 U377 (.Z(n539), 
	.S(n395), 
	.B(n565), 
	.A(n564));
   MUX2_X1 U378 (.Z(n411), 
	.S(n395), 
	.B(n567), 
	.A(n566));
   MUX2_X1 U379 (.Z(B[10]), 
	.S(SH[2]), 
	.B(n525), 
	.A(n405));
   INV_X1 U380 (.ZN(n525), 
	.A(n568));
   MUX2_X1 U381 (.Z(n568), 
	.S(SH[4]), 
	.B(n454), 
	.A(n569));
   NAND2_X1 U382 (.ZN(n454), 
	.A2(n392), 
	.A1(n570));
   INV_X1 U383 (.ZN(n570), 
	.A(n546));
   MUX2_X1 U384 (.Z(n546), 
	.S(n395), 
	.B(n553), 
	.A(n561));
   NAND2_X1 U385 (.ZN(n553), 
	.A2(n383), 
	.A1(A[31]));
   MUX2_X1 U386 (.Z(n569), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n571), 
	.A(n548));
   MUX2_X1 U387 (.Z(n548), 
	.S(n395), 
	.B(n556), 
	.A(n565));
   MUX2_X1 U388 (.Z(n556), 
	.S(SH[3]), 
	.B(n573), 
	.A(n572));
   MUX2_X1 U389 (.Z(n565), 
	.S(SH[3]), 
	.B(n575), 
	.A(n574));
   INV_X1 U390 (.ZN(n405), 
	.A(n576));
   MUX2_X1 U391 (.Z(n576), 
	.S(SH[4]), 
	.B(n470), 
	.A(n577));
   MUX2_X1 U392 (.Z(n470), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n545), 
	.A(n480));
   MUX2_X1 U393 (.Z(n545), 
	.S(n395), 
	.B(n560), 
	.A(n563));
   MUX2_X1 U394 (.Z(n480), 
	.S(n395), 
	.B(n562), 
	.A(n504));
   MUX2_X1 U395 (.Z(n577), 
	.S(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n547), 
	.A(n417));
   MUX2_X1 U396 (.Z(n547), 
	.S(n395), 
	.B(n564), 
	.A(n567));
   MUX2_X1 U397 (.Z(n564), 
	.S(SH[3]), 
	.B(n579), 
	.A(n578));
   MUX2_X1 U398 (.Z(n567), 
	.S(SH[3]), 
	.B(n581), 
	.A(n580));
   MUX2_X1 U399 (.Z(n417), 
	.S(n395), 
	.B(n566), 
	.A(n424));
   MUX2_X1 U400 (.Z(n566), 
	.S(SH[3]), 
	.B(n583), 
	.A(n582));
   MUX2_X1 U401 (.Z(n424), 
	.S(SH[3]), 
	.B(n585), 
	.A(n584));
   MUX2_X1 U402 (.Z(B[0]), 
	.S(SH[2]), 
	.B(n412), 
	.A(n586));
   INV_X1 U403 (.ZN(n412), 
	.A(n587));
   MUX2_X1 U404 (.Z(n587), 
	.S(SH[4]), 
	.B(n518), 
	.A(n588));
   MUX2_X1 U405 (.Z(n518), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n508), 
	.A(n529));
   MUX2_X1 U406 (.Z(n508), 
	.S(n395), 
	.B(n514), 
	.A(n524));
   MUX2_X1 U407 (.Z(n514), 
	.S(SH[3]), 
	.B(n589), 
	.A(n573));
   INV_X1 U408 (.ZN(n589), 
	.A(A[31]));
   MUX2_X1 U409 (.Z(n524), 
	.S(SH[3]), 
	.B(n590), 
	.A(n575));
   MUX2_X1 U410 (.Z(n529), 
	.S(n394), 
	.B(n523), 
	.A(n534));
   MUX2_X1 U411 (.Z(n523), 
	.S(SH[3]), 
	.B(n591), 
	.A(n579));
   MUX2_X1 U412 (.Z(n534), 
	.S(SH[3]), 
	.B(n592), 
	.A(n581));
   MUX2_X1 U413 (.Z(n588), 
	.S(SH[1]), 
	.B(n436), 
	.A(n444));
   MUX2_X1 U414 (.Z(n436), 
	.S(n394), 
	.B(n485), 
	.A(n489));
   MUX2_X1 U415 (.Z(n485), 
	.S(SH[3]), 
	.B(n572), 
	.A(n593));
   MUX2_X1 U416 (.Z(n489), 
	.S(SH[3]), 
	.B(n574), 
	.A(n594));
   MUX2_X1 U417 (.Z(n444), 
	.S(n394), 
	.B(n488), 
	.A(n495));
   MUX2_X1 U418 (.Z(n488), 
	.S(SH[3]), 
	.B(n578), 
	.A(n595));
   MUX2_X1 U419 (.Z(n495), 
	.S(SH[3]), 
	.B(n580), 
	.A(n596));
   MUX2_X1 U420 (.Z(n586), 
	.S(SH[4]), 
	.B(n542), 
	.A(n597));
   INV_X1 U421 (.ZN(n542), 
	.A(n598));
   MUX2_X1 U422 (.Z(n598), 
	.S(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.B(n528), 
	.A(n571));
   MUX2_X1 U423 (.Z(n528), 
	.S(n394), 
	.B(n533), 
	.A(n555));
   MUX2_X1 U424 (.Z(n533), 
	.S(SH[3]), 
	.B(n599), 
	.A(n583));
   MUX2_X1 U425 (.Z(n555), 
	.S(SH[3]), 
	.B(n600), 
	.A(n585));
   MUX2_X1 U426 (.Z(n571), 
	.S(n394), 
	.B(n554), 
	.A(n557));
   MUX2_X1 U427 (.Z(n554), 
	.S(SH[3]), 
	.B(n601), 
	.A(n439));
   MUX2_X1 U428 (.Z(n557), 
	.S(SH[3]), 
	.B(n602), 
	.A(n487));
   MUX2_X1 U429 (.Z(n597), 
	.S(SH[1]), 
	.B(n442), 
	.A(n603));
   INV_X1 U430 (.ZN(n442), 
	.A(n604));
   MUX2_X1 U431 (.Z(n604), 
	.S(n394), 
	.B(n494), 
	.A(n498));
   MUX2_X1 U432 (.Z(n494), 
	.S(SH[3]), 
	.B(n582), 
	.A(n605));
   MUX2_X1 U433 (.Z(n498), 
	.S(SH[3]), 
	.B(n584), 
	.A(n606));
   MUX2_X1 U434 (.Z(n603), 
	.S(n394), 
	.B(n496), 
	.A(n607));
   INV_X1 U435 (.ZN(n496), 
	.A(n608));
   MUX2_X1 U436 (.Z(n608), 
	.S(SH[3]), 
	.B(n438), 
	.A(n609));
   MUX2_X1 U437 (.Z(n607), 
	.S(SH[3]), 
	.B(A[8]), 
	.A(A[0]));
endmodule

module up_island_DW_mult_tc_1 (
	a, 
	b, 
	product, 
	FE_PT1_n796, 
	FE_PT1_n705, 
	FE_PT1_n654, 
	FE_PT1_n617, 
	FE_PT1_n582, 
	n531, 
	FE_PT1_n477, 
	n338, 
	FE_PT1_n808, 
	FE_PT1_n949);
   input [31:0] a;
   input [31:0] b;
   output [63:0] product;
   input FE_PT1_n796;
   input FE_PT1_n705;
   input FE_PT1_n654;
   input FE_PT1_n617;
   input FE_PT1_n582;
   input n531;
   input FE_PT1_n477;
   input n338;
   input FE_PT1_n808;
   input FE_PT1_n949;

   // Internal wires
   wire FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_;
   wire FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_;
   wire FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_;
   wire FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_;
   wire FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_;
   wire FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_;
   wire FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_;
   wire FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_;
   wire FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_;
   wire FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_;
   wire FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_;
   wire FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_;
   wire FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_;
   wire FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_;
   wire FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_;
   wire FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_;
   wire FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_;
   wire FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_;
   wire FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_;
   wire FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_;
   wire FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_;
   wire FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_;
   wire FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_;
   wire FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_;
   wire FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_;
   wire FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_;
   wire FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_;
   wire FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_;
   wire FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_;
   wire FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_;
   wire FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_;
   wire FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_;
   wire FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_;
   wire FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_;
   wire FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_;
   wire FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_;
   wire FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_;
   wire FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_;
   wire FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_;
   wire FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_;
   wire FE_OFN81_n3137;
   wire FE_OFN78_n3121;
   wire FE_OFN75_n3136;
   wire FE_OFN72_n3120;
   wire FE_OFN70_n3135;
   wire FE_OFN67_n3119;
   wire FE_OFN66_n3134;
   wire FE_OFN65_n3118;
   wire FE_OFN64_n3133;
   wire FE_OFN61_n3117;
   wire FE_OFN58_n3132;
   wire FE_OFN55_n3116;
   wire FE_OFN52_n3131;
   wire FE_OFN51_n3115;
   wire FE_OFN48_n3130;
   wire FE_OFN47_n3114;
   wire FE_OFN46_n3129;
   wire FE_OFN45_n3113;
   wire FE_OFN44_n3128;
   wire FE_OFN43_n3112;
   wire FE_OFN42_n3127;
   wire FE_OFN41_n3111;
   wire FE_OFN40_n3126;
   wire FE_OFN39_n3110;
   wire FE_OFN38_n3125;
   wire FE_OFN37_n3109;
   wire FE_OFN36_n3124;
   wire FE_OFN35_n3123;
   wire FE_OFN34_n3107;
   wire FE_OFN33_n3108;
   wire FE_OFN32_n765;
   wire n8;
   wire n10;
   wire n14;
   wire n15;
   wire n24;
   wire n26;
   wire n30;
   wire n31;
   wire n40;
   wire n60;
   wire n82;
   wire n83;
   wire n92;
   wire n94;
   wire n98;
   wire n99;
   wire n108;
   wire n110;
   wire n114;
   wire n115;
   wire n124;
   wire n126;
   wire n130;
   wire n131;
   wire n140;
   wire n142;
   wire n146;
   wire n147;
   wire n156;
   wire n158;
   wire n162;
   wire n163;
   wire n167;
   wire n172;
   wire n173;
   wire n174;
   wire n178;
   wire n179;
   wire n188;
   wire n189;
   wire n190;
   wire n194;
   wire n195;
   wire n204;
   wire n205;
   wire n206;
   wire n210;
   wire n211;
   wire n220;
   wire n221;
   wire n222;
   wire n226;
   wire n227;
   wire n236;
   wire n238;
   wire n242;
   wire n243;
   wire n252;
   wire n254;
   wire n258;
   wire n259;
   wire n263;
   wire n268;
   wire n270;
   wire n274;
   wire n275;
   wire n284;
   wire n286;
   wire n290;
   wire n291;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1013;
   wire n1016;
   wire n1020;
   wire n1025;
   wire n1026;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1038;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1060;
   wire n1061;
   wire n1069;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3145;
   wire n3146;
   wire n3153;

   BUF_X2 FE_OFC178_UUT_Mpath_the_mult_x_operand1_31_ (.Z(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(a[31]));
   BUF_X2 FE_OFC174_UUT_Mpath_the_mult_x_operand1_23_ (.Z(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(a[23]));
   BUF_X2 FE_OFC172_UUT_Mpath_the_mult_x_operand1_1_ (.Z(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(a[1]));
   BUF_X1 FE_OFC166_UUT_Mpath_the_mult_x_operand1_3_ (.Z(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(a[3]));
   CLKBUF_X1 FE_OFC161_UUT_Mpath_the_mult_x_operand2_3_ (.Z(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_), 
	.A(b[3]));
   CLKBUF_X1 FE_OFC158_UUT_Mpath_the_mult_x_operand2_4_ (.Z(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_), 
	.A(b[4]));
   BUF_X2 FE_OFC157_UUT_Mpath_the_mult_x_operand1_5_ (.Z(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(a[5]));
   CLKBUF_X1 FE_OFC155_UUT_Mpath_the_mult_x_operand2_5_ (.Z(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_), 
	.A(b[5]));
   CLKBUF_X1 FE_OFC154_UUT_Mpath_the_mult_x_operand2_6_ (.Z(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_), 
	.A(b[6]));
   BUF_X2 FE_OFC153_UUT_Mpath_the_mult_x_operand1_7_ (.Z(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(a[7]));
   CLKBUF_X1 FE_OFC151_UUT_Mpath_the_mult_x_operand2_7_ (.Z(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_), 
	.A(b[7]));
   BUF_X2 FE_OFC150_UUT_Mpath_the_mult_x_operand1_9_ (.Z(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(a[9]));
   CLKBUF_X1 FE_OFC148_UUT_Mpath_the_mult_x_operand2_9_ (.Z(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_), 
	.A(b[9]));
   BUF_X2 FE_OFC147_UUT_Mpath_the_mult_x_operand1_11_ (.Z(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(a[11]));
   CLKBUF_X1 FE_OFC145_UUT_Mpath_the_mult_x_operand2_11_ (.Z(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_), 
	.A(b[11]));
   CLKBUF_X1 FE_OFC144_UUT_Mpath_the_mult_x_operand2_12_ (.Z(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_), 
	.A(b[12]));
   BUF_X2 FE_OFC143_UUT_Mpath_the_mult_x_operand1_13_ (.Z(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(a[13]));
   CLKBUF_X1 FE_OFC141_UUT_Mpath_the_mult_x_operand2_13_ (.Z(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_), 
	.A(b[13]));
   BUF_X2 FE_OFC139_UUT_Mpath_the_mult_x_operand1_15_ (.Z(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(a[15]));
   BUF_X2 FE_OFC135_UUT_Mpath_the_mult_x_operand1_17_ (.Z(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(a[17]));
   CLKBUF_X1 FE_OFC132_UUT_Mpath_the_mult_x_operand2_18_ (.Z(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_), 
	.A(b[18]));
   BUF_X1 FE_OFC131_UUT_Mpath_the_mult_x_operand1_19_ (.Z(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(a[19]));
   CLKBUF_X1 FE_OFC128_UUT_Mpath_the_mult_x_operand2_20_ (.Z(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_), 
	.A(b[20]));
   BUF_X2 FE_OFC127_UUT_Mpath_the_mult_x_operand1_21_ (.Z(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(a[21]));
   CLKBUF_X1 FE_OFC125_UUT_Mpath_the_mult_x_operand2_21_ (.Z(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_), 
	.A(b[21]));
   CLKBUF_X1 FE_OFC124_UUT_Mpath_the_mult_x_operand2_22_ (.Z(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_), 
	.A(b[22]));
   CLKBUF_X1 FE_OFC123_UUT_Mpath_the_mult_x_operand2_24_ (.Z(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_), 
	.A(b[24]));
   BUF_X2 FE_OFC122_UUT_Mpath_the_mult_x_operand1_25_ (.Z(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(a[25]));
   CLKBUF_X1 FE_OFC119_UUT_Mpath_the_mult_x_operand2_26_ (.Z(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_), 
	.A(b[26]));
   BUF_X2 FE_OFC118_UUT_Mpath_the_mult_x_operand1_27_ (.Z(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(a[27]));
   CLKBUF_X1 FE_OFC116_UUT_Mpath_the_mult_x_operand2_27_ (.Z(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_), 
	.A(b[27]));
   CLKBUF_X1 FE_OFC115_UUT_Mpath_the_mult_x_operand2_28_ (.Z(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_), 
	.A(b[28]));
   BUF_X2 FE_OFC114_UUT_Mpath_the_mult_x_operand1_29_ (.Z(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(a[29]));
   CLKBUF_X1 FE_OFC112_UUT_Mpath_the_mult_x_operand2_29_ (.Z(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_), 
	.A(b[29]));
   CLKBUF_X1 FE_OFC111_UUT_Mpath_the_mult_x_operand2_30_ (.Z(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_), 
	.A(b[30]));
   CLKBUF_X1 FE_OFC110_UUT_Mpath_the_mult_x_operand2_23_ (.Z(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_), 
	.A(b[23]));
   CLKBUF_X1 FE_OFC109_UUT_Mpath_the_mult_x_operand2_8_ (.Z(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_), 
	.A(b[8]));
   CLKBUF_X1 FE_OFC108_UUT_Mpath_the_mult_x_operand2_10_ (.Z(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_), 
	.A(b[10]));
   CLKBUF_X1 FE_OFC107_UUT_Mpath_the_mult_x_operand2_31_ (.Z(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_), 
	.A(b[31]));
   BUF_X1 FE_OFC106_UUT_Mpath_the_mult_x_operand2_0_ (.Z(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_), 
	.A(b[0]));
   BUF_X2 FE_OFC81_n3137 (.Z(FE_OFN81_n3137), 
	.A(n3137));
   BUF_X2 FE_OFC78_n3121 (.Z(FE_OFN78_n3121), 
	.A(n3121));
   BUF_X2 FE_OFC75_n3136 (.Z(FE_OFN75_n3136), 
	.A(n3136));
   BUF_X2 FE_OFC72_n3120 (.Z(FE_OFN72_n3120), 
	.A(n3120));
   BUF_X2 FE_OFC70_n3135 (.Z(FE_OFN70_n3135), 
	.A(n3135));
   BUF_X2 FE_OFC67_n3119 (.Z(FE_OFN67_n3119), 
	.A(n3119));
   BUF_X2 FE_OFC66_n3134 (.Z(FE_OFN66_n3134), 
	.A(n3134));
   BUF_X2 FE_OFC65_n3118 (.Z(FE_OFN65_n3118), 
	.A(n3118));
   BUF_X2 FE_OFC64_n3133 (.Z(FE_OFN64_n3133), 
	.A(n3133));
   BUF_X2 FE_OFC61_n3117 (.Z(FE_OFN61_n3117), 
	.A(n3117));
   BUF_X2 FE_OFC58_n3132 (.Z(FE_OFN58_n3132), 
	.A(n3132));
   BUF_X2 FE_OFC55_n3116 (.Z(FE_OFN55_n3116), 
	.A(n3116));
   BUF_X2 FE_OFC52_n3131 (.Z(FE_OFN52_n3131), 
	.A(n3131));
   BUF_X2 FE_OFC51_n3115 (.Z(FE_OFN51_n3115), 
	.A(n3115));
   BUF_X2 FE_OFC48_n3130 (.Z(FE_OFN48_n3130), 
	.A(n3130));
   BUF_X2 FE_OFC47_n3114 (.Z(FE_OFN47_n3114), 
	.A(n3114));
   BUF_X2 FE_OFC46_n3129 (.Z(FE_OFN46_n3129), 
	.A(n3129));
   BUF_X2 FE_OFC45_n3113 (.Z(FE_OFN45_n3113), 
	.A(n3113));
   BUF_X2 FE_OFC44_n3128 (.Z(FE_OFN44_n3128), 
	.A(n3128));
   BUF_X2 FE_OFC43_n3112 (.Z(FE_OFN43_n3112), 
	.A(n3112));
   BUF_X2 FE_OFC42_n3127 (.Z(FE_OFN42_n3127), 
	.A(n3127));
   BUF_X2 FE_OFC41_n3111 (.Z(FE_OFN41_n3111), 
	.A(n3111));
   BUF_X2 FE_OFC40_n3126 (.Z(FE_OFN40_n3126), 
	.A(n3126));
   BUF_X2 FE_OFC39_n3110 (.Z(FE_OFN39_n3110), 
	.A(n3110));
   BUF_X2 FE_OFC38_n3125 (.Z(FE_OFN38_n3125), 
	.A(n3125));
   BUF_X2 FE_OFC37_n3109 (.Z(FE_OFN37_n3109), 
	.A(n3109));
   BUF_X2 FE_OFC36_n3124 (.Z(FE_OFN36_n3124), 
	.A(n3124));
   BUF_X2 FE_OFC35_n3123 (.Z(FE_OFN35_n3123), 
	.A(n3123));
   BUF_X2 FE_OFC34_n3107 (.Z(FE_OFN34_n3107), 
	.A(n3107));
   BUF_X2 FE_OFC33_n3108 (.Z(FE_OFN33_n3108), 
	.A(n3108));
   CLKBUF_X2 FE_OFC32_n765 (.Z(FE_OFN32_n765), 
	.A(n765));
   NAND2_X1 OR_NOTi (.ZN(n3058), 
	.A2(a[1]), 
	.A1(n263));
   NAND2_X1 AND_NOTi (.ZN(n291), 
	.A2(n290), 
	.A1(b[0]));
   INV_X1 U2 (.ZN(product[0]), 
	.A(n291));
   INV_X1 U11 (.ZN(n290), 
	.A(n3138));
   OAI21_X1 AO21i (.ZN(n2499), 
	.B2(n290), 
	.B1(n284), 
	.A(n286));
   INV_X1 U3 (.ZN(n286), 
	.A(n3026));
   INV_X1 U12 (.ZN(n284), 
	.A(n3122));
   NAND2_X1 OR_NOTi1 (.ZN(n3025), 
	.A2(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A1(n263));
   NAND2_X1 AND_NOTi1 (.ZN(n275), 
	.A2(n274), 
	.A1(b[0]));
   INV_X1 U22 (.ZN(n2498), 
	.A(n275));
   INV_X1 U14 (.ZN(n274), 
	.A(FE_OFN81_n3137));
   OAI21_X1 AO21i1 (.ZN(n2467), 
	.B2(n274), 
	.B1(n268), 
	.A(n270));
   INV_X1 U31 (.ZN(n270), 
	.A(n2993));
   INV_X1 U15 (.ZN(n268), 
	.A(FE_OFN78_n3121));
   NAND2_X1 OR_NOTi2 (.ZN(n2992), 
	.A2(a[5]), 
	.A1(n263));
   INV_X1 U16 (.ZN(n263), 
	.A(b[0]));
   NAND2_X1 AND_NOTi2 (.ZN(n259), 
	.A2(n258), 
	.A1(b[0]));
   INV_X1 U24 (.ZN(n2466), 
	.A(n259));
   INV_X1 U17 (.ZN(n258), 
	.A(FE_OFN75_n3136));
   OAI21_X1 AO21i2 (.ZN(n2435), 
	.B2(n258), 
	.B1(n252), 
	.A(n254));
   INV_X1 U32 (.ZN(n254), 
	.A(n2960));
   INV_X1 U18 (.ZN(n252), 
	.A(FE_OFN72_n3120));
   NAND2_X1 OR_NOTi3 (.ZN(n2959), 
	.A2(a[7]), 
	.A1(n263));
   NAND2_X1 AND_NOTi3 (.ZN(n243), 
	.A2(n242), 
	.A1(b[0]));
   INV_X1 U26 (.ZN(n2434), 
	.A(n243));
   INV_X1 U110 (.ZN(n242), 
	.A(FE_OFN70_n3135));
   OAI21_X1 AO21i3 (.ZN(n2403), 
	.B2(n242), 
	.B1(n236), 
	.A(n238));
   INV_X1 U33 (.ZN(n238), 
	.A(n2927));
   INV_X1 U111 (.ZN(n236), 
	.A(FE_OFN67_n3119));
   NAND2_X1 OR_NOTi4 (.ZN(n2926), 
	.A2(a[9]), 
	.A1(n263));
   NAND2_X1 AND_NOTi4 (.ZN(n227), 
	.A2(n226), 
	.A1(b[0]));
   INV_X1 U28 (.ZN(n2402), 
	.A(n227));
   INV_X1 U113 (.ZN(n226), 
	.A(n3134));
   OAI21_X1 AO21i4 (.ZN(n2371), 
	.B2(n221), 
	.B1(n220), 
	.A(n222));
   INV_X1 U34 (.ZN(n222), 
	.A(n2894));
   INV_X1 U29 (.ZN(n221), 
	.A(FE_OFN66_n3134));
   INV_X1 U114 (.ZN(n220), 
	.A(FE_OFN65_n3118));
   NAND2_X1 OR_NOTi5 (.ZN(n2893), 
	.A2(a[11]), 
	.A1(n263));
   NAND2_X1 AND_NOTi5 (.ZN(n211), 
	.A2(n210), 
	.A1(b[0]));
   INV_X1 U210 (.ZN(n2370), 
	.A(n211));
   INV_X1 U116 (.ZN(n210), 
	.A(n3133));
   OAI21_X1 AO21i5 (.ZN(n2339), 
	.B2(n205), 
	.B1(n204), 
	.A(n206));
   INV_X1 U35 (.ZN(n206), 
	.A(n2861));
   INV_X1 U211 (.ZN(n205), 
	.A(FE_OFN64_n3133));
   INV_X1 U117 (.ZN(n204), 
	.A(FE_OFN61_n3117));
   NAND2_X1 OR_NOTi6 (.ZN(n2860), 
	.A2(a[13]), 
	.A1(n263));
   NAND2_X1 AND_NOTi6 (.ZN(n195), 
	.A2(n194), 
	.A1(b[0]));
   INV_X1 U212 (.ZN(n2338), 
	.A(n195));
   INV_X1 U119 (.ZN(n194), 
	.A(n3132));
   OAI21_X1 AO21i6 (.ZN(n2307), 
	.B2(n189), 
	.B1(n188), 
	.A(n190));
   INV_X1 U36 (.ZN(n190), 
	.A(n2828));
   INV_X1 U213 (.ZN(n189), 
	.A(FE_OFN58_n3132));
   INV_X1 U120 (.ZN(n188), 
	.A(FE_OFN55_n3116));
   NAND2_X1 OR_NOTi7 (.ZN(n2827), 
	.A2(a[15]), 
	.A1(n263));
   NAND2_X1 AND_NOTi7 (.ZN(n179), 
	.A2(n178), 
	.A1(b[0]));
   INV_X1 U214 (.ZN(n2306), 
	.A(n179));
   INV_X1 U122 (.ZN(n178), 
	.A(n3131));
   OAI21_X1 AO21i7 (.ZN(n2275), 
	.B2(n173), 
	.B1(n172), 
	.A(n174));
   INV_X1 U37 (.ZN(n174), 
	.A(n2795));
   INV_X1 U215 (.ZN(n173), 
	.A(FE_OFN52_n3131));
   INV_X1 U123 (.ZN(n172), 
	.A(FE_OFN51_n3115));
   NAND2_X1 OR_NOTi8 (.ZN(n2794), 
	.A2(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A1(n167));
   INV_X1 U124 (.ZN(n167), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   NAND2_X1 AND_NOTi8 (.ZN(n163), 
	.A2(n162), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U216 (.ZN(n2274), 
	.A(n163));
   INV_X1 U125 (.ZN(n162), 
	.A(FE_OFN48_n3130));
   OAI21_X1 AO21i8 (.ZN(n2243), 
	.B2(n162), 
	.B1(n156), 
	.A(n158));
   INV_X1 U38 (.ZN(n158), 
	.A(n2762));
   INV_X1 U126 (.ZN(n156), 
	.A(FE_OFN47_n3114));
   NAND2_X1 OR_NOTi9 (.ZN(n2761), 
	.A2(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A1(n167));
   NAND2_X1 AND_NOTi9 (.ZN(n147), 
	.A2(n146), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U218 (.ZN(n2242), 
	.A(n147));
   INV_X1 U128 (.ZN(n146), 
	.A(FE_OFN46_n3129));
   OAI21_X1 AO21i9 (.ZN(n2211), 
	.B2(n146), 
	.B1(n140), 
	.A(n142));
   INV_X1 U39 (.ZN(n142), 
	.A(n2729));
   INV_X1 U129 (.ZN(n140), 
	.A(FE_OFN45_n3113));
   NAND2_X1 OR_NOTi10 (.ZN(n2728), 
	.A2(a[21]), 
	.A1(n167));
   NAND2_X1 AND_NOTi10 (.ZN(n131), 
	.A2(n130), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U220 (.ZN(n2210), 
	.A(n131));
   INV_X1 U131 (.ZN(n130), 
	.A(FE_OFN44_n3128));
   OAI21_X1 AO21i10 (.ZN(n2179), 
	.B2(n130), 
	.B1(n124), 
	.A(n126));
   INV_X1 U310 (.ZN(n126), 
	.A(n2696));
   INV_X1 U132 (.ZN(n124), 
	.A(FE_OFN43_n3112));
   NAND2_X1 OR_NOTi11 (.ZN(n2695), 
	.A2(a[23]), 
	.A1(n167));
   NAND2_X1 AND_NOTi11 (.ZN(n115), 
	.A2(n114), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U222 (.ZN(n2178), 
	.A(n115));
   INV_X1 U134 (.ZN(n114), 
	.A(FE_OFN42_n3127));
   OAI21_X1 AO21i11 (.ZN(n2147), 
	.B2(n114), 
	.B1(n108), 
	.A(n110));
   INV_X1 U311 (.ZN(n110), 
	.A(n2663));
   INV_X1 U135 (.ZN(n108), 
	.A(FE_OFN41_n3111));
   NAND2_X1 OR_NOTi12 (.ZN(n2662), 
	.A2(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A1(n167));
   NAND2_X1 AND_NOTi12 (.ZN(n99), 
	.A2(n98), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U224 (.ZN(n2146), 
	.A(n99));
   INV_X1 U137 (.ZN(n98), 
	.A(FE_OFN40_n3126));
   OAI21_X1 AO21i12 (.ZN(n2115), 
	.B2(n98), 
	.B1(n92), 
	.A(n94));
   INV_X1 U312 (.ZN(n94), 
	.A(n2630));
   INV_X1 U138 (.ZN(n92), 
	.A(FE_OFN39_n3110));
   NAND2_X1 OR_NOTi13 (.ZN(n2629), 
	.A2(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A1(n167));
   NAND2_X1 AND_NOTi13 (.ZN(n83), 
	.A2(n82), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U226 (.ZN(n2114), 
	.A(n83));
   INV_X1 U140 (.ZN(n82), 
	.A(FE_OFN38_n3125));
   OAI21_X1 AO21i13 (.ZN(n2083), 
	.B2(n82), 
	.B1(n40), 
	.A(n60));
   INV_X1 U313 (.ZN(n60), 
	.A(n2597));
   INV_X1 U141 (.ZN(n40), 
	.A(FE_OFN37_n3109));
   NAND2_X1 OR_NOTi14 (.ZN(n2596), 
	.A2(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A1(n167));
   NAND2_X1 AND_NOTi14 (.ZN(n31), 
	.A2(n30), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U228 (.ZN(n2082), 
	.A(n31));
   INV_X1 U143 (.ZN(n30), 
	.A(FE_OFN36_n3124));
   OAI21_X1 AO21i14 (.ZN(n2051), 
	.B2(n30), 
	.B1(n24), 
	.A(n26));
   INV_X1 U314 (.ZN(n26), 
	.A(n2564));
   INV_X1 U144 (.ZN(n24), 
	.A(FE_OFN33_n3108));
   NAND2_X1 OR_NOTi15 (.ZN(n2563), 
	.A2(a[31]), 
	.A1(n263));
   NAND2_X1 AND_NOTi15 (.ZN(n15), 
	.A2(n14), 
	.A1(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   INV_X1 U230 (.ZN(n2050), 
	.A(n15));
   INV_X1 U146 (.ZN(n14), 
	.A(FE_OFN35_n3123));
   OAI21_X1 AO21i15 (.ZN(n2019), 
	.B2(n14), 
	.B1(n8), 
	.A(n10));
   INV_X1 U315 (.ZN(n10), 
	.A(n2531));
   INV_X1 U147 (.ZN(n8), 
	.A(FE_OFN34_n3107));
   INV_X1 U242 (.ZN(product[63]), 
	.A(n510));
   XNOR2_X1 U243 (.ZN(product[62]), 
	.B(n448), 
	.A(n517));
   OAI21_X1 U244 (.ZN(n510), 
	.B2(n511), 
	.B1(FE_OFN32_n765), 
	.A(n512));
   NAND2_X1 U245 (.ZN(n511), 
	.A2(n513), 
	.A1(n520));
   AOI21_X1 U246 (.ZN(n512), 
	.B2(n513), 
	.B1(n521), 
	.A(n514));
   INV_X1 U247 (.ZN(n513), 
	.A(n515));
   INV_X1 U248 (.ZN(n514), 
	.A(n516));
   NAND2_X1 U249 (.ZN(n448), 
	.A2(n516), 
	.A1(n513));
   NOR2_X1 U251 (.ZN(n515), 
	.A2(n1073), 
	.A1(n2019));
   NAND2_X1 U252 (.ZN(n516), 
	.A2(n1073), 
	.A1(n2019));
   XNOR2_X1 U253 (.ZN(product[61]), 
	.B(n449), 
	.A(n528));
   OAI21_X1 U254 (.ZN(n517), 
	.B2(n518), 
	.B1(FE_OFN32_n765), 
	.A(n519));
   INV_X1 U255 (.ZN(n518), 
	.A(n520));
   INV_X1 U256 (.ZN(n519), 
	.A(n521));
   NOR2_X1 U257 (.ZN(n520), 
	.A2(n522), 
	.A1(n682));
   OAI21_X1 U258 (.ZN(n521), 
	.B2(n522), 
	.B1(n683), 
	.A(n523));
   NAND2_X1 U259 (.ZN(n522), 
	.A2(n524), 
	.A1(n533));
   AOI21_X1 U260 (.ZN(n523), 
	.B2(n524), 
	.B1(n534), 
	.A(n525));
   INV_X1 U261 (.ZN(n524), 
	.A(n526));
   INV_X1 U262 (.ZN(n525), 
	.A(n527));
   NAND2_X1 U263 (.ZN(n449), 
	.A2(n527), 
	.A1(n524));
   NOR2_X1 U265 (.ZN(n526), 
	.A2(n1074), 
	.A1(n1075));
   NAND2_X1 U266 (.ZN(n527), 
	.A2(n1074), 
	.A1(n1075));
   XNOR2_X1 U267 (.ZN(product[60]), 
	.B(n450), 
	.A(n537));
   OAI21_X1 U268 (.ZN(n528), 
	.B2(n529), 
	.B1(FE_OFN32_n765), 
	.A(n530));
   NAND2_X1 U269 (.ZN(n529), 
	.A2(n533), 
	.A1(n680));
   AOI21_X1 U270 (.ZN(n530), 
	.B2(n533), 
	.B1(n681), 
	.A(n534));
   NOR2_X1 U273 (.ZN(n533), 
	.A2(n535), 
	.A1(n542));
   OAI21_X1 U274 (.ZN(n534), 
	.B2(n535), 
	.B1(n543), 
	.A(n536));
   NAND2_X1 U275 (.ZN(n450), 
	.A2(n536), 
	.A1(n1013));
   INV_X1 U276 (.ZN(n1013), 
	.A(n535));
   NOR2_X1 U277 (.ZN(n535), 
	.A2(n1076), 
	.A1(n1077));
   NAND2_X1 U278 (.ZN(n536), 
	.A2(n1076), 
	.A1(n1077));
   XNOR2_X1 U279 (.ZN(product[59]), 
	.B(n451), 
	.A(n552));
   OAI21_X1 U280 (.ZN(n537), 
	.B2(n538), 
	.B1(FE_OFN32_n765), 
	.A(n539));
   NAND2_X1 U281 (.ZN(n538), 
	.A2(n540), 
	.A1(n680));
   AOI21_X1 U282 (.ZN(n539), 
	.B2(n540), 
	.B1(n681), 
	.A(n541));
   INV_X1 U283 (.ZN(n540), 
	.A(n542));
   INV_X1 U284 (.ZN(n541), 
	.A(n543));
   NAND2_X1 U285 (.ZN(n542), 
	.A2(n544), 
	.A1(n651));
   AOI21_X1 U286 (.ZN(n543), 
	.B2(n652), 
	.B1(n544), 
	.A(n545));
   NOR2_X1 U287 (.ZN(n544), 
	.A2(n546), 
	.A1(n616));
   OAI21_X1 U288 (.ZN(n545), 
	.B2(n546), 
	.B1(n617), 
	.A(n547));
   NAND2_X1 U289 (.ZN(n546), 
	.A2(n548), 
	.A1(n557));
   AOI21_X1 U290 (.ZN(n547), 
	.B2(n548), 
	.B1(n558), 
	.A(n549));
   INV_X1 U291 (.ZN(n548), 
	.A(n550));
   INV_X1 U292 (.ZN(n549), 
	.A(n551));
   NAND2_X1 U293 (.ZN(n451), 
	.A2(n551), 
	.A1(n548));
   NOR2_X1 U295 (.ZN(n550), 
	.A2(n1081), 
	.A1(n1078));
   NAND2_X1 U296 (.ZN(n551), 
	.A2(n1081), 
	.A1(n1078));
   XNOR2_X1 U297 (.ZN(product[58]), 
	.B(n452), 
	.A(n565));
   OAI21_X1 U298 (.ZN(n552), 
	.B2(n553), 
	.B1(FE_OFN32_n765), 
	.A(n554));
   NAND2_X1 U299 (.ZN(n553), 
	.A2(n557), 
	.A1(n608));
   AOI21_X1 U300 (.ZN(n554), 
	.B2(n557), 
	.B1(n609), 
	.A(n558));
   NOR2_X1 U303 (.ZN(n557), 
	.A2(n559), 
	.A1(n590));
   OAI21_X1 U304 (.ZN(n558), 
	.B2(n559), 
	.B1(n591), 
	.A(n560));
   NAND2_X1 U305 (.ZN(n559), 
	.A2(n561), 
	.A1(n570));
   AOI21_X1 U306 (.ZN(n560), 
	.B2(n561), 
	.B1(n571), 
	.A(n562));
   INV_X1 U307 (.ZN(n561), 
	.A(n563));
   INV_X1 U308 (.ZN(n562), 
	.A(n564));
   NAND2_X1 U309 (.ZN(n452), 
	.A2(n564), 
	.A1(n561));
   NOR2_X1 U317 (.ZN(n563), 
	.A2(n1082), 
	.A1(n1085));
   NAND2_X1 U318 (.ZN(n564), 
	.A2(n1082), 
	.A1(n1085));
   XNOR2_X1 U319 (.ZN(product[57]), 
	.B(n453), 
	.A(n574));
   OAI21_X1 U320 (.ZN(n565), 
	.B2(n566), 
	.B1(n765), 
	.A(n567));
   NAND2_X1 U321 (.ZN(n566), 
	.A2(n570), 
	.A1(n584));
   AOI21_X1 U322 (.ZN(n567), 
	.B2(n570), 
	.B1(n585), 
	.A(n571));
   NOR2_X1 U325 (.ZN(n570), 
	.A2(n572), 
	.A1(n579));
   OAI21_X1 U326 (.ZN(n571), 
	.B2(n572), 
	.B1(n580), 
	.A(n573));
   NAND2_X1 U327 (.ZN(n453), 
	.A2(n573), 
	.A1(n1016));
   INV_X1 U328 (.ZN(n1016), 
	.A(n572));
   NOR2_X1 U329 (.ZN(n572), 
	.A2(n1091), 
	.A1(n1086));
   NAND2_X1 U330 (.ZN(n573), 
	.A2(n1091), 
	.A1(n1086));
   XNOR2_X1 U331 (.ZN(product[56]), 
	.B(n454), 
	.A(n581));
   OAI21_X1 U332 (.ZN(n574), 
	.B2(n575), 
	.B1(n765), 
	.A(n576));
   NAND2_X1 U333 (.ZN(n575), 
	.A2(n577), 
	.A1(n584));
   AOI21_X1 U334 (.ZN(n576), 
	.B2(n577), 
	.B1(n585), 
	.A(n578));
   INV_X1 U335 (.ZN(n577), 
	.A(n579));
   INV_X1 U336 (.ZN(n578), 
	.A(n580));
   NAND2_X1 U337 (.ZN(n454), 
	.A2(n580), 
	.A1(n577));
   NOR2_X1 U339 (.ZN(n579), 
	.A2(n1097), 
	.A1(n1092));
   NAND2_X1 U340 (.ZN(n580), 
	.A2(n1097), 
	.A1(n1092));
   XNOR2_X1 U341 (.ZN(product[55]), 
	.B(n455), 
	.A(n596));
   OAI21_X1 U342 (.ZN(n581), 
	.B2(n582), 
	.B1(n765), 
	.A(n583));
   INV_X1 U343 (.ZN(n582), 
	.A(n584));
   INV_X1 U344 (.ZN(n583), 
	.A(n585));
   NOR2_X1 U345 (.ZN(n584), 
	.A2(n586), 
	.A1(n682));
   OAI21_X1 U346 (.ZN(n585), 
	.B2(n586), 
	.B1(n683), 
	.A(n587));
   NAND2_X1 U347 (.ZN(n586), 
	.A2(n588), 
	.A1(n612));
   AOI21_X1 U348 (.ZN(n587), 
	.B2(n588), 
	.B1(n613), 
	.A(n589));
   INV_X1 U349 (.ZN(n588), 
	.A(n590));
   INV_X1 U350 (.ZN(n589), 
	.A(n591));
   NAND2_X1 U351 (.ZN(n590), 
	.A2(n592), 
	.A1(n601));
   AOI21_X1 U352 (.ZN(n591), 
	.B2(n592), 
	.B1(n602), 
	.A(n593));
   INV_X1 U353 (.ZN(n592), 
	.A(n594));
   INV_X1 U354 (.ZN(n593), 
	.A(n595));
   NAND2_X1 U355 (.ZN(n455), 
	.A2(n595), 
	.A1(n592));
   NOR2_X1 U357 (.ZN(n594), 
	.A2(n1105), 
	.A1(n1098));
   NAND2_X1 U358 (.ZN(n595), 
	.A2(n1105), 
	.A1(n1098));
   XNOR2_X1 U359 (.ZN(product[54]), 
	.B(n456), 
	.A(n605));
   OAI21_X1 U360 (.ZN(n596), 
	.B2(n597), 
	.B1(FE_OFN32_n765), 
	.A(n598));
   NAND2_X1 U361 (.ZN(n597), 
	.A2(n601), 
	.A1(n608));
   AOI21_X1 U362 (.ZN(n598), 
	.B2(n601), 
	.B1(n609), 
	.A(n602));
   INV_X1 U365 (.ZN(n601), 
	.A(n603));
   INV_X1 U366 (.ZN(n602), 
	.A(n604));
   NAND2_X1 U367 (.ZN(n456), 
	.A2(n604), 
	.A1(n601));
   NOR2_X1 U369 (.ZN(n603), 
	.A2(n1113), 
	.A1(n1106));
   NAND2_X1 U370 (.ZN(n604), 
	.A2(n1113), 
	.A1(n1106));
   XNOR2_X1 U371 (.ZN(product[53]), 
	.B(n457), 
	.A(n622));
   OAI21_X1 U372 (.ZN(n605), 
	.B2(n606), 
	.B1(FE_OFN32_n765), 
	.A(n607));
   INV_X1 U373 (.ZN(n606), 
	.A(n608));
   INV_X1 U374 (.ZN(n607), 
	.A(n609));
   NOR2_X1 U375 (.ZN(n608), 
	.A2(n610), 
	.A1(n682));
   OAI21_X1 U376 (.ZN(n609), 
	.B2(n610), 
	.B1(n683), 
	.A(n611));
   INV_X1 U377 (.ZN(n610), 
	.A(n612));
   INV_X1 U378 (.ZN(n611), 
	.A(n613));
   NOR2_X1 U379 (.ZN(n612), 
	.A2(n616), 
	.A1(n649));
   OAI21_X1 U380 (.ZN(n613), 
	.B2(n616), 
	.B1(n650), 
	.A(n617));
   NAND2_X1 U383 (.ZN(n616), 
	.A2(n638), 
	.A1(n618));
   AOI21_X1 U384 (.ZN(n617), 
	.B2(n639), 
	.B1(n618), 
	.A(n619));
   NOR2_X1 U385 (.ZN(n618), 
	.A2(n620), 
	.A1(n627));
   OAI21_X1 U386 (.ZN(n619), 
	.B2(n620), 
	.B1(n628), 
	.A(n621));
   NAND2_X1 U387 (.ZN(n457), 
	.A2(n621), 
	.A1(n1020));
   INV_X1 U388 (.ZN(n1020), 
	.A(n620));
   NOR2_X1 U389 (.ZN(n620), 
	.A2(n1123), 
	.A1(n1114));
   NAND2_X1 U390 (.ZN(n621), 
	.A2(n1123), 
	.A1(n1114));
   XNOR2_X1 U391 (.ZN(product[52]), 
	.B(n458), 
	.A(n629));
   OAI21_X1 U392 (.ZN(n622), 
	.B2(n623), 
	.B1(FE_OFN32_n765), 
	.A(n624));
   NAND2_X1 U393 (.ZN(n623), 
	.A2(n625), 
	.A1(n632));
   AOI21_X1 U394 (.ZN(n624), 
	.B2(n625), 
	.B1(n633), 
	.A(n626));
   INV_X1 U395 (.ZN(n625), 
	.A(n627));
   INV_X1 U396 (.ZN(n626), 
	.A(n628));
   NAND2_X1 U397 (.ZN(n458), 
	.A2(n628), 
	.A1(n625));
   NOR2_X1 U399 (.ZN(n627), 
	.A2(n1133), 
	.A1(n1124));
   NAND2_X1 U400 (.ZN(n628), 
	.A2(n1133), 
	.A1(n1124));
   XNOR2_X1 U401 (.ZN(product[51]), 
	.B(n459), 
	.A(n642));
   OAI21_X1 U402 (.ZN(n629), 
	.B2(n630), 
	.B1(FE_OFN32_n765), 
	.A(n631));
   INV_X1 U403 (.ZN(n630), 
	.A(n632));
   INV_X1 U404 (.ZN(n631), 
	.A(n633));
   NOR2_X1 U405 (.ZN(n632), 
	.A2(n634), 
	.A1(n682));
   OAI21_X1 U406 (.ZN(n633), 
	.B2(n634), 
	.B1(n683), 
	.A(n635));
   NAND2_X1 U407 (.ZN(n634), 
	.A2(n638), 
	.A1(n647));
   AOI21_X1 U408 (.ZN(n635), 
	.B2(n638), 
	.B1(n648), 
	.A(n639));
   INV_X1 U411 (.ZN(n638), 
	.A(n640));
   INV_X1 U412 (.ZN(n639), 
	.A(n641));
   NAND2_X1 U413 (.ZN(n459), 
	.A2(n641), 
	.A1(n638));
   NOR2_X1 U415 (.ZN(n640), 
	.A2(n1145), 
	.A1(n1134));
   NAND2_X1 U416 (.ZN(n641), 
	.A2(n1145), 
	.A1(n1134));
   XNOR2_X1 U417 (.ZN(product[50]), 
	.B(n460), 
	.A(n659));
   OAI21_X1 U418 (.ZN(n642), 
	.B2(n643), 
	.B1(FE_OFN32_n765), 
	.A(n644));
   NAND2_X1 U419 (.ZN(n643), 
	.A2(n647), 
	.A1(n680));
   AOI21_X1 U420 (.ZN(n644), 
	.B2(n647), 
	.B1(n681), 
	.A(n648));
   INV_X1 U423 (.ZN(n647), 
	.A(n649));
   INV_X1 U424 (.ZN(n648), 
	.A(n650));
   INV_X1 U425 (.ZN(n649), 
	.A(n651));
   INV_X1 U426 (.ZN(n650), 
	.A(n652));
   NOR2_X1 U427 (.ZN(n651), 
	.A2(n653), 
	.A1(n675));
   OAI21_X1 U428 (.ZN(n652), 
	.B2(n676), 
	.B1(n653), 
	.A(n654));
   NAND2_X1 U429 (.ZN(n653), 
	.A2(n655), 
	.A1(n664));
   AOI21_X1 U430 (.ZN(n654), 
	.B2(n655), 
	.B1(n665), 
	.A(n656));
   INV_X1 U431 (.ZN(n655), 
	.A(n657));
   INV_X1 U432 (.ZN(n656), 
	.A(n658));
   NAND2_X1 U433 (.ZN(n460), 
	.A2(n658), 
	.A1(n655));
   NOR2_X1 U435 (.ZN(n657), 
	.A2(n1146), 
	.A1(n1157));
   NAND2_X1 U436 (.ZN(n658), 
	.A2(n1146), 
	.A1(n1157));
   XNOR2_X1 U437 (.ZN(product[49]), 
	.B(n461), 
	.A(n668));
   OAI21_X1 U438 (.ZN(n659), 
	.B2(n660), 
	.B1(FE_OFN32_n765), 
	.A(n661));
   NAND2_X1 U439 (.ZN(n660), 
	.A2(n664), 
	.A1(n671));
   AOI21_X1 U440 (.ZN(n661), 
	.B2(n664), 
	.B1(n672), 
	.A(n665));
   INV_X1 U443 (.ZN(n664), 
	.A(n666));
   INV_X1 U444 (.ZN(n665), 
	.A(n667));
   NAND2_X1 U445 (.ZN(n461), 
	.A2(n667), 
	.A1(n664));
   NOR2_X1 U447 (.ZN(n666), 
	.A2(n1171), 
	.A1(n1158));
   NAND2_X1 U448 (.ZN(n667), 
	.A2(n1171), 
	.A1(n1158));
   XNOR2_X1 U449 (.ZN(product[48]), 
	.B(n462), 
	.A(n677));
   OAI21_X1 U450 (.ZN(n668), 
	.B2(n669), 
	.B1(FE_OFN32_n765), 
	.A(n670));
   INV_X1 U451 (.ZN(n669), 
	.A(n671));
   INV_X1 U452 (.ZN(n670), 
	.A(n672));
   NOR2_X1 U453 (.ZN(n671), 
	.A2(n675), 
	.A1(n682));
   OAI21_X1 U454 (.ZN(n672), 
	.B2(n675), 
	.B1(n683), 
	.A(n676));
   NAND2_X1 U457 (.ZN(n462), 
	.A2(n676), 
	.A1(n1025));
   INV_X1 U458 (.ZN(n1025), 
	.A(n675));
   NOR2_X1 U459 (.ZN(n675), 
	.A2(n1185), 
	.A1(n1172));
   NAND2_X1 U460 (.ZN(n676), 
	.A2(n1185), 
	.A1(n1172));
   XNOR2_X1 U461 (.ZN(product[47]), 
	.B(n463), 
	.A(n692));
   OAI21_X1 U462 (.ZN(n677), 
	.B2(n678), 
	.B1(FE_OFN32_n765), 
	.A(n679));
   INV_X1 U463 (.ZN(n678), 
	.A(n680));
   INV_X1 U464 (.ZN(n679), 
	.A(n681));
   INV_X1 U465 (.ZN(n680), 
	.A(n682));
   INV_X1 U466 (.ZN(n681), 
	.A(n683));
   NAND2_X1 U467 (.ZN(n682), 
	.A2(n684), 
	.A1(n741));
   AOI21_X1 U468 (.ZN(n683), 
	.B2(n742), 
	.B1(n684), 
	.A(n685));
   NOR2_X1 U469 (.ZN(n684), 
	.A2(n719), 
	.A1(n686));
   OAI21_X1 U470 (.ZN(n685), 
	.B2(n720), 
	.B1(n686), 
	.A(n687));
   NAND2_X1 U471 (.ZN(n686), 
	.A2(n708), 
	.A1(n688));
   AOI21_X1 U472 (.ZN(n687), 
	.B2(n709), 
	.B1(n688), 
	.A(n689));
   NOR2_X1 U473 (.ZN(n688), 
	.A2(n690), 
	.A1(n697));
   OAI21_X1 U474 (.ZN(n689), 
	.B2(n698), 
	.B1(n690), 
	.A(n691));
   NAND2_X1 U475 (.ZN(n463), 
	.A2(n691), 
	.A1(n1026));
   INV_X1 U476 (.ZN(n1026), 
	.A(n690));
   NOR2_X1 U477 (.ZN(n690), 
	.A2(n1201), 
	.A1(n1186));
   NAND2_X1 U478 (.ZN(n691), 
	.A2(n1201), 
	.A1(n1186));
   XNOR2_X1 U479 (.ZN(product[46]), 
	.B(n464), 
	.A(n699));
   OAI21_X1 U480 (.ZN(n692), 
	.B2(n693), 
	.B1(FE_OFN32_n765), 
	.A(n694));
   NAND2_X1 U481 (.ZN(n693), 
	.A2(n695), 
	.A1(n702));
   AOI21_X1 U482 (.ZN(n694), 
	.B2(n695), 
	.B1(n703), 
	.A(n696));
   INV_X1 U483 (.ZN(n695), 
	.A(n697));
   INV_X1 U484 (.ZN(n696), 
	.A(n698));
   NAND2_X1 U485 (.ZN(n464), 
	.A2(n698), 
	.A1(n695));
   NOR2_X1 U487 (.ZN(n697), 
	.A2(n1217), 
	.A1(n1202));
   NAND2_X1 U488 (.ZN(n698), 
	.A2(n1217), 
	.A1(n1202));
   XNOR2_X1 U489 (.ZN(product[45]), 
	.B(n465), 
	.A(n712));
   OAI21_X1 U490 (.ZN(n699), 
	.B2(n700), 
	.B1(FE_OFN32_n765), 
	.A(n701));
   INV_X1 U491 (.ZN(n700), 
	.A(n702));
   INV_X1 U492 (.ZN(n701), 
	.A(n703));
   NOR2_X1 U493 (.ZN(n702), 
	.A2(n704), 
	.A1(n739));
   OAI21_X1 U494 (.ZN(n703), 
	.B2(n704), 
	.B1(n740), 
	.A(n705));
   NAND2_X1 U495 (.ZN(n704), 
	.A2(n708), 
	.A1(n717));
   AOI21_X1 U496 (.ZN(n705), 
	.B2(n708), 
	.B1(n718), 
	.A(n709));
   INV_X1 U499 (.ZN(n708), 
	.A(n710));
   INV_X1 U500 (.ZN(n709), 
	.A(n711));
   NAND2_X1 U501 (.ZN(n465), 
	.A2(n711), 
	.A1(n708));
   NOR2_X1 U503 (.ZN(n710), 
	.A2(n1235), 
	.A1(n1218));
   NAND2_X1 U504 (.ZN(n711), 
	.A2(n1235), 
	.A1(n1218));
   XNOR2_X1 U505 (.ZN(product[44]), 
	.B(n466), 
	.A(n725));
   OAI21_X1 U506 (.ZN(n712), 
	.B2(n713), 
	.B1(FE_OFN32_n765), 
	.A(n714));
   NAND2_X1 U507 (.ZN(n713), 
	.A2(n717), 
	.A1(n737));
   AOI21_X1 U508 (.ZN(n714), 
	.B2(n717), 
	.B1(n738), 
	.A(n718));
   INV_X1 U511 (.ZN(n717), 
	.A(n719));
   INV_X1 U512 (.ZN(n718), 
	.A(n720));
   NAND2_X1 U513 (.ZN(n719), 
	.A2(n721), 
	.A1(n730));
   AOI21_X1 U514 (.ZN(n720), 
	.B2(n731), 
	.B1(n721), 
	.A(n722));
   INV_X1 U515 (.ZN(n721), 
	.A(n723));
   INV_X1 U516 (.ZN(n722), 
	.A(n724));
   NAND2_X1 U517 (.ZN(n466), 
	.A2(n724), 
	.A1(n721));
   NOR2_X1 U519 (.ZN(n723), 
	.A2(n1253), 
	.A1(n1236));
   NAND2_X1 U520 (.ZN(n724), 
	.A2(n1253), 
	.A1(n1236));
   XNOR2_X1 U521 (.ZN(product[43]), 
	.B(n467), 
	.A(n734));
   OAI21_X1 U522 (.ZN(n725), 
	.B2(n726), 
	.B1(FE_OFN32_n765), 
	.A(n727));
   NAND2_X1 U523 (.ZN(n726), 
	.A2(n730), 
	.A1(n737));
   AOI21_X1 U524 (.ZN(n727), 
	.B2(n730), 
	.B1(n738), 
	.A(n731));
   INV_X1 U527 (.ZN(n730), 
	.A(n732));
   INV_X1 U528 (.ZN(n731), 
	.A(n733));
   NAND2_X1 U529 (.ZN(n467), 
	.A2(n733), 
	.A1(n730));
   NOR2_X1 U531 (.ZN(n732), 
	.A2(n1273), 
	.A1(n1254));
   NAND2_X1 U532 (.ZN(n733), 
	.A2(n1273), 
	.A1(n1254));
   XNOR2_X1 U533 (.ZN(product[42]), 
	.B(n468), 
	.A(n749));
   OAI21_X1 U534 (.ZN(n734), 
	.B2(n735), 
	.B1(FE_OFN32_n765), 
	.A(n736));
   INV_X1 U535 (.ZN(n735), 
	.A(n737));
   INV_X1 U536 (.ZN(n736), 
	.A(n738));
   INV_X1 U537 (.ZN(n737), 
	.A(n739));
   INV_X1 U538 (.ZN(n738), 
	.A(n740));
   INV_X1 U539 (.ZN(n739), 
	.A(n741));
   INV_X1 U540 (.ZN(n740), 
	.A(n742));
   NOR2_X1 U541 (.ZN(n741), 
	.A2(n743), 
	.A1(n763));
   OAI21_X1 U542 (.ZN(n742), 
	.B2(n764), 
	.B1(n743), 
	.A(n744));
   NAND2_X1 U543 (.ZN(n743), 
	.A2(n745), 
	.A1(n754));
   AOI21_X1 U544 (.ZN(n744), 
	.B2(n755), 
	.B1(n745), 
	.A(n746));
   INV_X1 U545 (.ZN(n745), 
	.A(n747));
   INV_X1 U546 (.ZN(n746), 
	.A(n748));
   NAND2_X1 U547 (.ZN(n468), 
	.A2(n748), 
	.A1(n745));
   NOR2_X1 U549 (.ZN(n747), 
	.A2(n1293), 
	.A1(n1274));
   NAND2_X1 U550 (.ZN(n748), 
	.A2(n1293), 
	.A1(n1274));
   XNOR2_X1 U551 (.ZN(product[41]), 
	.B(n469), 
	.A(n758));
   OAI21_X1 U552 (.ZN(n749), 
	.B2(n750), 
	.B1(FE_OFN32_n765), 
	.A(n751));
   NAND2_X1 U553 (.ZN(n750), 
	.A2(n754), 
	.A1(n761));
   AOI21_X1 U554 (.ZN(n751), 
	.B2(n754), 
	.B1(n762), 
	.A(n755));
   INV_X1 U557 (.ZN(n754), 
	.A(n756));
   INV_X1 U558 (.ZN(n755), 
	.A(n757));
   NAND2_X1 U559 (.ZN(n469), 
	.A2(n757), 
	.A1(n754));
   NOR2_X1 U561 (.ZN(n756), 
	.A2(n1315), 
	.A1(n1294));
   NAND2_X1 U562 (.ZN(n757), 
	.A2(n1315), 
	.A1(n1294));
   XOR2_X1 U563 (.Z(product[40]), 
	.B(n470), 
	.A(FE_OFN32_n765));
   OAI21_X1 U564 (.ZN(n758), 
	.B2(n759), 
	.B1(FE_OFN32_n765), 
	.A(n760));
   INV_X1 U565 (.ZN(n759), 
	.A(n761));
   INV_X1 U566 (.ZN(n760), 
	.A(n762));
   INV_X1 U567 (.ZN(n761), 
	.A(n763));
   INV_X1 U568 (.ZN(n762), 
	.A(n764));
   NAND2_X1 U569 (.ZN(n470), 
	.A2(n764), 
	.A1(n761));
   NOR2_X1 U571 (.ZN(n763), 
	.A2(n1337), 
	.A1(n1316));
   NAND2_X1 U572 (.ZN(n764), 
	.A2(n1337), 
	.A1(n1316));
   XNOR2_X1 U573 (.ZN(product[39]), 
	.B(n471), 
	.A(n774));
   AOI21_X1 U574 (.ZN(n765), 
	.B2(n834), 
	.B1(n766), 
	.A(n767));
   NOR2_X1 U575 (.ZN(n766), 
	.A2(n768), 
	.A1(n806));
   OAI21_X1 U576 (.ZN(n767), 
	.B2(n768), 
	.B1(n807), 
	.A(n769));
   NAND2_X1 U577 (.ZN(n768), 
	.A2(n770), 
	.A1(n790));
   AOI21_X1 U578 (.ZN(n769), 
	.B2(n791), 
	.B1(n770), 
	.A(n771));
   NOR2_X1 U579 (.ZN(n770), 
	.A2(n772), 
	.A1(n781));
   OAI21_X1 U580 (.ZN(n771), 
	.B2(n772), 
	.B1(n782), 
	.A(n773));
   NAND2_X1 U581 (.ZN(n471), 
	.A2(n773), 
	.A1(n1034));
   INV_X1 U582 (.ZN(n1034), 
	.A(n772));
   NOR2_X1 U583 (.ZN(n772), 
	.A2(n1361), 
	.A1(n1338));
   NAND2_X1 U584 (.ZN(n773), 
	.A2(n1361), 
	.A1(n1338));
   XNOR2_X1 U585 (.ZN(product[38]), 
	.B(n472), 
	.A(n783));
   OAI21_X1 U586 (.ZN(n774), 
	.B2(n833), 
	.B1(n775), 
	.A(n776));
   NAND2_X1 U587 (.ZN(n775), 
	.A2(n804), 
	.A1(n777));
   AOI21_X1 U588 (.ZN(n776), 
	.B2(n777), 
	.B1(n805), 
	.A(n778));
   NOR2_X1 U589 (.ZN(n777), 
	.A2(n781), 
	.A1(n788));
   OAI21_X1 U590 (.ZN(n778), 
	.B2(n781), 
	.B1(n789), 
	.A(n782));
   NAND2_X1 U593 (.ZN(n472), 
	.A2(n782), 
	.A1(n1035));
   INV_X1 U594 (.ZN(n1035), 
	.A(n781));
   NOR2_X1 U595 (.ZN(n781), 
	.A2(n1385), 
	.A1(n1362));
   NAND2_X1 U596 (.ZN(n782), 
	.A2(n1385), 
	.A1(n1362));
   XNOR2_X1 U597 (.ZN(product[37]), 
	.B(n473), 
	.A(n794));
   OAI21_X1 U598 (.ZN(n783), 
	.B2(n784), 
	.B1(n833), 
	.A(n785));
   NAND2_X1 U599 (.ZN(n784), 
	.A2(n786), 
	.A1(n804));
   AOI21_X1 U600 (.ZN(n785), 
	.B2(n786), 
	.B1(n805), 
	.A(n787));
   INV_X1 U601 (.ZN(n786), 
	.A(n788));
   INV_X1 U602 (.ZN(n787), 
	.A(n789));
   INV_X1 U603 (.ZN(n788), 
	.A(n790));
   INV_X1 U604 (.ZN(n789), 
	.A(n791));
   NOR2_X1 U605 (.ZN(n790), 
	.A2(n792), 
	.A1(n799));
   OAI21_X1 U606 (.ZN(n791), 
	.B2(n800), 
	.B1(n792), 
	.A(n793));
   NAND2_X1 U607 (.ZN(n473), 
	.A2(n793), 
	.A1(n1036));
   INV_X1 U608 (.ZN(n1036), 
	.A(n792));
   NOR2_X1 U609 (.ZN(n792), 
	.A2(n1411), 
	.A1(n1386));
   NAND2_X1 U610 (.ZN(n793), 
	.A2(n1411), 
	.A1(n1386));
   XNOR2_X1 U611 (.ZN(product[36]), 
	.B(n474), 
	.A(n801));
   OAI21_X1 U612 (.ZN(n794), 
	.B2(n795), 
	.B1(n833), 
	.A(n796));
   NAND2_X1 U613 (.ZN(n795), 
	.A2(n797), 
	.A1(n804));
   AOI21_X1 U614 (.ZN(n796), 
	.B2(n797), 
	.B1(n805), 
	.A(n798));
   INV_X1 U615 (.ZN(n797), 
	.A(n799));
   INV_X1 U616 (.ZN(n798), 
	.A(n800));
   NAND2_X1 U617 (.ZN(n474), 
	.A2(n800), 
	.A1(n797));
   NOR2_X1 U619 (.ZN(n799), 
	.A2(n1437), 
	.A1(n1412));
   NAND2_X1 U620 (.ZN(n800), 
	.A2(n1437), 
	.A1(n1412));
   XNOR2_X1 U621 (.ZN(product[35]), 
	.B(n475), 
	.A(n812));
   OAI21_X1 U622 (.ZN(n801), 
	.B2(n802), 
	.B1(n833), 
	.A(n803));
   INV_X1 U623 (.ZN(n802), 
	.A(n804));
   INV_X1 U624 (.ZN(n803), 
	.A(n805));
   INV_X1 U625 (.ZN(n804), 
	.A(n806));
   INV_X1 U626 (.ZN(n805), 
	.A(n807));
   NAND2_X1 U627 (.ZN(n806), 
	.A2(n808), 
	.A1(n826));
   AOI21_X1 U628 (.ZN(n807), 
	.B2(n827), 
	.B1(n808), 
	.A(n809));
   NOR2_X1 U629 (.ZN(n808), 
	.A2(n817), 
	.A1(n810));
   OAI21_X1 U630 (.ZN(n809), 
	.B2(n818), 
	.B1(n810), 
	.A(n811));
   NAND2_X1 U631 (.ZN(n475), 
	.A2(n811), 
	.A1(n1038));
   INV_X1 U632 (.ZN(n1038), 
	.A(n810));
   NOR2_X1 U633 (.ZN(n810), 
	.A2(n1465), 
	.A1(n1438));
   NAND2_X1 U634 (.ZN(n811), 
	.A2(n1465), 
	.A1(n1438));
   XNOR2_X1 U635 (.ZN(product[34]), 
	.B(n476), 
	.A(n819));
   OAI21_X1 U636 (.ZN(n812), 
	.B2(n813), 
	.B1(n833), 
	.A(n814));
   NAND2_X1 U637 (.ZN(n813), 
	.A2(n815), 
	.A1(n826));
   AOI21_X1 U638 (.ZN(n814), 
	.B2(n815), 
	.B1(n827), 
	.A(n816));
   INV_X1 U639 (.ZN(n815), 
	.A(n817));
   INV_X1 U640 (.ZN(n816), 
	.A(n818));
   NAND2_X1 U641 (.ZN(n476), 
	.A2(n818), 
	.A1(n815));
   NOR2_X1 U643 (.ZN(n817), 
	.A2(n1493), 
	.A1(n1466));
   NAND2_X1 U644 (.ZN(n818), 
	.A2(n1493), 
	.A1(n1466));
   XNOR2_X1 U645 (.ZN(product[33]), 
	.B(n477), 
	.A(n830));
   OAI21_X1 U646 (.ZN(n819), 
	.B2(n820), 
	.B1(n833), 
	.A(n821));
   INV_X1 U647 (.ZN(n820), 
	.A(n826));
   INV_X1 U648 (.ZN(n821), 
	.A(n827));
   NOR2_X1 U653 (.ZN(n826), 
	.A2(n828), 
	.A1(n831));
   OAI21_X1 U654 (.ZN(n827), 
	.B2(n832), 
	.B1(n828), 
	.A(n829));
   NAND2_X1 U655 (.ZN(n477), 
	.A2(n829), 
	.A1(n1040));
   INV_X1 U656 (.ZN(n1040), 
	.A(n828));
   NOR2_X1 U657 (.ZN(n828), 
	.A2(n1523), 
	.A1(n1494));
   NAND2_X1 U658 (.ZN(n829), 
	.A2(n1523), 
	.A1(n1494));
   XOR2_X1 U659 (.Z(product[32]), 
	.B(n478), 
	.A(n833));
   OAI21_X1 U660 (.ZN(n830), 
	.B2(n831), 
	.B1(n833), 
	.A(n832));
   NAND2_X1 U661 (.ZN(n478), 
	.A2(n832), 
	.A1(n1041));
   INV_X1 U662 (.ZN(n1041), 
	.A(n831));
   NOR2_X1 U663 (.ZN(n831), 
	.A2(n1553), 
	.A1(n1524));
   NAND2_X1 U664 (.ZN(n832), 
	.A2(n1553), 
	.A1(n1524));
   XNOR2_X1 U665 (.ZN(product[31]), 
	.B(n479), 
	.A(n841));
   INV_X1 U666 (.ZN(n833), 
	.A(n834));
   OAI21_X1 U667 (.ZN(n834), 
	.B2(n855), 
	.B1(n835), 
	.A(n836));
   NAND2_X1 U668 (.ZN(n835), 
	.A2(n845), 
	.A1(n837));
   AOI21_X1 U669 (.ZN(n836), 
	.B2(n846), 
	.B1(n837), 
	.A(n838));
   NOR2_X1 U670 (.ZN(n837), 
	.A2(n839), 
	.A1(n842));
   OAI21_X1 U671 (.ZN(n838), 
	.B2(n843), 
	.B1(n839), 
	.A(n840));
   NAND2_X1 U672 (.ZN(n479), 
	.A2(n840), 
	.A1(n1042));
   INV_X1 U673 (.ZN(n1042), 
	.A(n839));
   NOR2_X1 U674 (.ZN(n839), 
	.A2(n1583), 
	.A1(n1554));
   NAND2_X1 U675 (.ZN(n840), 
	.A2(n1583), 
	.A1(n1554));
   XOR2_X1 U676 (.Z(product[30]), 
	.B(n480), 
	.A(n844));
   OAI21_X1 U677 (.ZN(n841), 
	.B2(n842), 
	.B1(n844), 
	.A(n843));
   NAND2_X1 U678 (.ZN(n480), 
	.A2(n843), 
	.A1(n1043));
   INV_X1 U679 (.ZN(n1043), 
	.A(n842));
   NOR2_X1 U680 (.ZN(n842), 
	.A2(n1611), 
	.A1(n1584));
   NAND2_X1 U681 (.ZN(n843), 
	.A2(n1611), 
	.A1(n1584));
   XOR2_X1 U682 (.Z(product[29]), 
	.B(n481), 
	.A(n849));
   AOI21_X1 U683 (.ZN(n844), 
	.B2(n845), 
	.B1(n854), 
	.A(n846));
   NOR2_X1 U684 (.ZN(n845), 
	.A2(n852), 
	.A1(n847));
   OAI21_X1 U685 (.ZN(n846), 
	.B2(n853), 
	.B1(n847), 
	.A(n848));
   NAND2_X1 U686 (.ZN(n481), 
	.A2(n848), 
	.A1(n1044));
   INV_X1 U687 (.ZN(n1044), 
	.A(n847));
   NOR2_X1 U688 (.ZN(n847), 
	.A2(n1639), 
	.A1(n1612));
   NAND2_X1 U689 (.ZN(n848), 
	.A2(n1639), 
	.A1(n1612));
   XNOR2_X1 U690 (.ZN(product[28]), 
	.B(n482), 
	.A(n854));
   AOI21_X1 U691 (.ZN(n849), 
	.B2(n850), 
	.B1(n854), 
	.A(n851));
   INV_X1 U692 (.ZN(n850), 
	.A(n852));
   INV_X1 U693 (.ZN(n851), 
	.A(n853));
   NAND2_X1 U694 (.ZN(n482), 
	.A2(n853), 
	.A1(n850));
   NOR2_X1 U696 (.ZN(n852), 
	.A2(n1665), 
	.A1(n1640));
   NAND2_X1 U697 (.ZN(n853), 
	.A2(n1665), 
	.A1(n1640));
   XOR2_X1 U698 (.Z(product[27]), 
	.B(n483), 
	.A(n864));
   INV_X1 U699 (.ZN(n854), 
	.A(n855));
   AOI21_X1 U700 (.ZN(n855), 
	.B2(n856), 
	.B1(n884), 
	.A(n857));
   NOR2_X1 U701 (.ZN(n856), 
	.A2(n870), 
	.A1(n858));
   OAI21_X1 U702 (.ZN(n857), 
	.B2(n858), 
	.B1(n871), 
	.A(n859));
   NAND2_X1 U703 (.ZN(n858), 
	.A2(n865), 
	.A1(n860));
   AOI21_X1 U704 (.ZN(n859), 
	.B2(n866), 
	.B1(n860), 
	.A(n861));
   INV_X1 U705 (.ZN(n860), 
	.A(n862));
   INV_X1 U706 (.ZN(n861), 
	.A(n863));
   NAND2_X1 U707 (.ZN(n483), 
	.A2(n863), 
	.A1(n860));
   NOR2_X1 U709 (.ZN(n862), 
	.A2(n1691), 
	.A1(n1666));
   NAND2_X1 U710 (.ZN(n863), 
	.A2(n1691), 
	.A1(n1666));
   XNOR2_X1 U711 (.ZN(product[26]), 
	.B(n484), 
	.A(n869));
   AOI21_X1 U712 (.ZN(n864), 
	.B2(n865), 
	.B1(n869), 
	.A(n866));
   INV_X1 U713 (.ZN(n865), 
	.A(n867));
   INV_X1 U714 (.ZN(n866), 
	.A(n868));
   NAND2_X1 U715 (.ZN(n484), 
	.A2(n868), 
	.A1(n865));
   NOR2_X1 U717 (.ZN(n867), 
	.A2(n1715), 
	.A1(n1692));
   NAND2_X1 U718 (.ZN(n868), 
	.A2(n1715), 
	.A1(n1692));
   XNOR2_X1 U719 (.ZN(product[25]), 
	.B(n485), 
	.A(n876));
   OAI21_X1 U720 (.ZN(n869), 
	.B2(n870), 
	.B1(n883), 
	.A(n871));
   NAND2_X1 U721 (.ZN(n870), 
	.A2(n879), 
	.A1(n872));
   AOI21_X1 U722 (.ZN(n871), 
	.B2(n880), 
	.B1(n872), 
	.A(n873));
   INV_X1 U723 (.ZN(n872), 
	.A(n874));
   INV_X1 U724 (.ZN(n873), 
	.A(n875));
   NAND2_X1 U725 (.ZN(n485), 
	.A2(n875), 
	.A1(n872));
   NOR2_X1 U727 (.ZN(n874), 
	.A2(n1739), 
	.A1(n1716));
   NAND2_X1 U728 (.ZN(n875), 
	.A2(n1739), 
	.A1(n1716));
   XOR2_X1 U729 (.Z(product[24]), 
	.B(n486), 
	.A(n883));
   OAI21_X1 U730 (.ZN(n876), 
	.B2(n877), 
	.B1(n883), 
	.A(n878));
   INV_X1 U731 (.ZN(n877), 
	.A(n879));
   INV_X1 U732 (.ZN(n878), 
	.A(n880));
   INV_X1 U733 (.ZN(n879), 
	.A(n881));
   INV_X1 U734 (.ZN(n880), 
	.A(n882));
   NAND2_X1 U735 (.ZN(n486), 
	.A2(n882), 
	.A1(n879));
   NOR2_X1 U737 (.ZN(n881), 
	.A2(n1761), 
	.A1(n1740));
   NAND2_X1 U738 (.ZN(n882), 
	.A2(n1761), 
	.A1(n1740));
   XNOR2_X1 U739 (.ZN(product[23]), 
	.B(n487), 
	.A(n891));
   INV_X1 U740 (.ZN(n883), 
	.A(n884));
   OAI21_X1 U741 (.ZN(n884), 
	.B2(n905), 
	.B1(n885), 
	.A(n886));
   NAND2_X1 U742 (.ZN(n885), 
	.A2(n895), 
	.A1(n887));
   AOI21_X1 U743 (.ZN(n886), 
	.B2(n896), 
	.B1(n887), 
	.A(n888));
   NOR2_X1 U744 (.ZN(n887), 
	.A2(n892), 
	.A1(n889));
   OAI21_X1 U745 (.ZN(n888), 
	.B2(n893), 
	.B1(n889), 
	.A(n890));
   NAND2_X1 U746 (.ZN(n487), 
	.A2(n890), 
	.A1(n1050));
   INV_X1 U747 (.ZN(n1050), 
	.A(n889));
   NOR2_X1 U748 (.ZN(n889), 
	.A2(n1783), 
	.A1(n1762));
   NAND2_X1 U749 (.ZN(n890), 
	.A2(n1783), 
	.A1(n1762));
   XOR2_X1 U750 (.Z(product[22]), 
	.B(n488), 
	.A(n894));
   OAI21_X1 U751 (.ZN(n891), 
	.B2(n892), 
	.B1(n894), 
	.A(n893));
   NAND2_X1 U752 (.ZN(n488), 
	.A2(n893), 
	.A1(n1051));
   INV_X1 U753 (.ZN(n1051), 
	.A(n892));
   NOR2_X1 U754 (.ZN(n892), 
	.A2(n1803), 
	.A1(n1784));
   NAND2_X1 U755 (.ZN(n893), 
	.A2(n1803), 
	.A1(n1784));
   XOR2_X1 U756 (.Z(product[21]), 
	.B(n489), 
	.A(n899));
   AOI21_X1 U757 (.ZN(n894), 
	.B2(n895), 
	.B1(n904), 
	.A(n896));
   NOR2_X1 U758 (.ZN(n895), 
	.A2(n902), 
	.A1(n897));
   OAI21_X1 U759 (.ZN(n896), 
	.B2(n903), 
	.B1(n897), 
	.A(n898));
   NAND2_X1 U760 (.ZN(n489), 
	.A2(n898), 
	.A1(n1052));
   INV_X1 U761 (.ZN(n1052), 
	.A(n897));
   NOR2_X1 U762 (.ZN(n897), 
	.A2(n1823), 
	.A1(n1804));
   NAND2_X1 U763 (.ZN(n898), 
	.A2(n1823), 
	.A1(n1804));
   XNOR2_X1 U764 (.ZN(product[20]), 
	.B(n490), 
	.A(n904));
   AOI21_X1 U765 (.ZN(n899), 
	.B2(n900), 
	.B1(n904), 
	.A(n901));
   INV_X1 U766 (.ZN(n900), 
	.A(n902));
   INV_X1 U767 (.ZN(n901), 
	.A(n903));
   NAND2_X1 U768 (.ZN(n490), 
	.A2(n903), 
	.A1(n900));
   NOR2_X1 U770 (.ZN(n902), 
	.A2(n1841), 
	.A1(n1824));
   NAND2_X1 U771 (.ZN(n903), 
	.A2(n1841), 
	.A1(n1824));
   XOR2_X1 U772 (.Z(product[19]), 
	.B(n491), 
	.A(n914));
   INV_X1 U773 (.ZN(n904), 
	.A(n905));
   AOI21_X1 U774 (.ZN(n905), 
	.B2(n934), 
	.B1(n906), 
	.A(n907));
   NOR2_X1 U775 (.ZN(n906), 
	.A2(n920), 
	.A1(n908));
   OAI21_X1 U776 (.ZN(n907), 
	.B2(n921), 
	.B1(n908), 
	.A(n909));
   NAND2_X1 U777 (.ZN(n908), 
	.A2(n915), 
	.A1(n910));
   AOI21_X1 U778 (.ZN(n909), 
	.B2(n916), 
	.B1(n910), 
	.A(n911));
   INV_X1 U779 (.ZN(n910), 
	.A(n912));
   INV_X1 U780 (.ZN(n911), 
	.A(n913));
   NAND2_X1 U781 (.ZN(n491), 
	.A2(n913), 
	.A1(n910));
   NOR2_X1 U783 (.ZN(n912), 
	.A2(n1859), 
	.A1(n1842));
   NAND2_X1 U784 (.ZN(n913), 
	.A2(n1859), 
	.A1(n1842));
   XNOR2_X1 U785 (.ZN(product[18]), 
	.B(n492), 
	.A(n919));
   AOI21_X1 U786 (.ZN(n914), 
	.B2(n915), 
	.B1(n919), 
	.A(n916));
   INV_X1 U787 (.ZN(n915), 
	.A(n917));
   INV_X1 U788 (.ZN(n916), 
	.A(n918));
   NAND2_X1 U789 (.ZN(n492), 
	.A2(n918), 
	.A1(n915));
   NOR2_X1 U791 (.ZN(n917), 
	.A2(n1875), 
	.A1(n1860));
   NAND2_X1 U792 (.ZN(n918), 
	.A2(n1875), 
	.A1(n1860));
   XNOR2_X1 U793 (.ZN(product[17]), 
	.B(n493), 
	.A(n926));
   OAI21_X1 U794 (.ZN(n919), 
	.B2(n920), 
	.B1(n933), 
	.A(n921));
   NAND2_X1 U795 (.ZN(n920), 
	.A2(n929), 
	.A1(n922));
   AOI21_X1 U796 (.ZN(n921), 
	.B2(n930), 
	.B1(n922), 
	.A(n923));
   INV_X1 U797 (.ZN(n922), 
	.A(n924));
   INV_X1 U798 (.ZN(n923), 
	.A(n925));
   NAND2_X1 U799 (.ZN(n493), 
	.A2(n925), 
	.A1(n922));
   NOR2_X1 U801 (.ZN(n924), 
	.A2(n1891), 
	.A1(n1876));
   NAND2_X1 U802 (.ZN(n925), 
	.A2(n1891), 
	.A1(n1876));
   XOR2_X1 U803 (.Z(product[16]), 
	.B(n494), 
	.A(n933));
   OAI21_X1 U804 (.ZN(n926), 
	.B2(n927), 
	.B1(n933), 
	.A(n928));
   INV_X1 U805 (.ZN(n927), 
	.A(n929));
   INV_X1 U806 (.ZN(n928), 
	.A(n930));
   INV_X1 U807 (.ZN(n929), 
	.A(n931));
   INV_X1 U808 (.ZN(n930), 
	.A(n932));
   NAND2_X1 U809 (.ZN(n494), 
	.A2(n932), 
	.A1(n929));
   NOR2_X1 U811 (.ZN(n931), 
	.A2(n1905), 
	.A1(n1892));
   NAND2_X1 U812 (.ZN(n932), 
	.A2(n1905), 
	.A1(n1892));
   XOR2_X1 U813 (.Z(product[15]), 
	.B(n495), 
	.A(n941));
   INV_X1 U814 (.ZN(n933), 
	.A(n934));
   OAI21_X1 U815 (.ZN(n934), 
	.B2(n935), 
	.B1(n947), 
	.A(n936));
   NAND2_X1 U816 (.ZN(n935), 
	.A2(n942), 
	.A1(n937));
   AOI21_X1 U817 (.ZN(n936), 
	.B2(n943), 
	.B1(n937), 
	.A(n938));
   INV_X1 U818 (.ZN(n937), 
	.A(n939));
   INV_X1 U819 (.ZN(n938), 
	.A(n940));
   NAND2_X1 U820 (.ZN(n495), 
	.A2(n940), 
	.A1(n937));
   NOR2_X1 U822 (.ZN(n939), 
	.A2(n1919), 
	.A1(n1906));
   NAND2_X1 U823 (.ZN(n940), 
	.A2(n1919), 
	.A1(n1906));
   XNOR2_X1 U824 (.ZN(product[14]), 
	.B(n496), 
	.A(n946));
   AOI21_X1 U825 (.ZN(n941), 
	.B2(n942), 
	.B1(n946), 
	.A(n943));
   INV_X1 U826 (.ZN(n942), 
	.A(n944));
   INV_X1 U827 (.ZN(n943), 
	.A(n945));
   NAND2_X1 U828 (.ZN(n496), 
	.A2(n945), 
	.A1(n942));
   NOR2_X1 U830 (.ZN(n944), 
	.A2(n1931), 
	.A1(n1920));
   NAND2_X1 U831 (.ZN(n945), 
	.A2(n1931), 
	.A1(n1920));
   XNOR2_X1 U832 (.ZN(product[13]), 
	.B(n497), 
	.A(n952));
   INV_X1 U833 (.ZN(n946), 
	.A(n947));
   AOI21_X1 U834 (.ZN(n947), 
	.B2(n956), 
	.B1(n948), 
	.A(n949));
   NOR2_X1 U835 (.ZN(n948), 
	.A2(n953), 
	.A1(n950));
   OAI21_X1 U836 (.ZN(n949), 
	.B2(n954), 
	.B1(n950), 
	.A(n951));
   NAND2_X1 U837 (.ZN(n497), 
	.A2(n951), 
	.A1(n1060));
   INV_X1 U838 (.ZN(n1060), 
	.A(n950));
   NOR2_X1 U839 (.ZN(n950), 
	.A2(n1943), 
	.A1(n1932));
   NAND2_X1 U840 (.ZN(n951), 
	.A2(n1943), 
	.A1(n1932));
   XOR2_X1 U841 (.Z(product[12]), 
	.B(n498), 
	.A(n955));
   OAI21_X1 U842 (.ZN(n952), 
	.B2(n953), 
	.B1(n955), 
	.A(n954));
   NAND2_X1 U843 (.ZN(n498), 
	.A2(n954), 
	.A1(n1061));
   INV_X1 U844 (.ZN(n1061), 
	.A(n953));
   NOR2_X1 U845 (.ZN(n953), 
	.A2(n1953), 
	.A1(n1944));
   NAND2_X1 U846 (.ZN(n954), 
	.A2(n1953), 
	.A1(n1944));
   XOR2_X1 U847 (.Z(product[11]), 
	.B(n499), 
	.A(n963));
   INV_X1 U848 (.ZN(n955), 
	.A(n956));
   OAI21_X1 U849 (.ZN(n956), 
	.B2(n969), 
	.B1(n957), 
	.A(n958));
   NAND2_X1 U850 (.ZN(n957), 
	.A2(n959), 
	.A1(n964));
   AOI21_X1 U851 (.ZN(n958), 
	.B2(n965), 
	.B1(n959), 
	.A(n960));
   INV_X1 U852 (.ZN(n959), 
	.A(n961));
   INV_X1 U853 (.ZN(n960), 
	.A(n962));
   NAND2_X1 U854 (.ZN(n499), 
	.A2(n962), 
	.A1(n959));
   NOR2_X1 U856 (.ZN(n961), 
	.A2(n1963), 
	.A1(n1954));
   NAND2_X1 U857 (.ZN(n962), 
	.A2(n1963), 
	.A1(n1954));
   XNOR2_X1 U858 (.ZN(product[10]), 
	.B(n968), 
	.A(n500));
   AOI21_X1 U859 (.ZN(n963), 
	.B2(n964), 
	.B1(n968), 
	.A(n965));
   INV_X1 U860 (.ZN(n964), 
	.A(n966));
   INV_X1 U861 (.ZN(n965), 
	.A(n967));
   NAND2_X1 U862 (.ZN(n500), 
	.A2(n967), 
	.A1(n964));
   NOR2_X1 U864 (.ZN(n966), 
	.A2(n1971), 
	.A1(n1964));
   NAND2_X1 U865 (.ZN(n967), 
	.A2(n1971), 
	.A1(n1964));
   XNOR2_X1 U866 (.ZN(product[9]), 
	.B(n974), 
	.A(n501));
   INV_X1 U867 (.ZN(n968), 
	.A(n969));
   AOI21_X1 U868 (.ZN(n969), 
	.B2(n970), 
	.B1(n974), 
	.A(n971));
   INV_X1 U869 (.ZN(n970), 
	.A(n972));
   INV_X1 U870 (.ZN(n971), 
	.A(n973));
   NAND2_X1 U871 (.ZN(n501), 
	.A2(n973), 
	.A1(n970));
   NOR2_X1 U873 (.ZN(n972), 
	.A2(n1979), 
	.A1(n1972));
   NAND2_X1 U874 (.ZN(n973), 
	.A2(n1979), 
	.A1(n1972));
   XOR2_X1 U875 (.Z(product[8]), 
	.B(n502), 
	.A(n981));
   OAI21_X1 U876 (.ZN(n974), 
	.B2(n987), 
	.B1(n975), 
	.A(n976));
   NAND2_X1 U877 (.ZN(n975), 
	.A2(n982), 
	.A1(n977));
   AOI21_X1 U878 (.ZN(n976), 
	.B2(n983), 
	.B1(n977), 
	.A(n978));
   INV_X1 U879 (.ZN(n977), 
	.A(n979));
   INV_X1 U880 (.ZN(n978), 
	.A(n980));
   NAND2_X1 U881 (.ZN(n502), 
	.A2(n980), 
	.A1(n977));
   NOR2_X1 U883 (.ZN(n979), 
	.A2(n1985), 
	.A1(n1980));
   NAND2_X1 U884 (.ZN(n980), 
	.A2(n1985), 
	.A1(n1980));
   XNOR2_X1 U885 (.ZN(product[7]), 
	.B(n503), 
	.A(n986));
   AOI21_X1 U886 (.ZN(n981), 
	.B2(n982), 
	.B1(n986), 
	.A(n983));
   INV_X1 U887 (.ZN(n982), 
	.A(n984));
   INV_X1 U888 (.ZN(n983), 
	.A(n985));
   NAND2_X1 U889 (.ZN(n503), 
	.A2(n985), 
	.A1(n982));
   NOR2_X1 U891 (.ZN(n984), 
	.A2(n1991), 
	.A1(n1986));
   NAND2_X1 U892 (.ZN(n985), 
	.A2(n1991), 
	.A1(n1986));
   XNOR2_X1 U893 (.ZN(product[6]), 
	.B(n992), 
	.A(n504));
   INV_X1 U894 (.ZN(n986), 
	.A(n987));
   AOI21_X1 U895 (.ZN(n987), 
	.B2(n992), 
	.B1(n988), 
	.A(n989));
   INV_X1 U896 (.ZN(n988), 
	.A(n990));
   INV_X1 U897 (.ZN(n989), 
	.A(n991));
   NAND2_X1 U898 (.ZN(n504), 
	.A2(n991), 
	.A1(n988));
   NOR2_X1 U900 (.ZN(n990), 
	.A2(n1995), 
	.A1(n1992));
   NAND2_X1 U901 (.ZN(n991), 
	.A2(n1995), 
	.A1(n1992));
   XNOR2_X1 U902 (.ZN(product[5]), 
	.B(n998), 
	.A(n505));
   INV_X1 U903 (.ZN(n992), 
	.A(n993));
   AOI21_X1 U904 (.ZN(n993), 
	.B2(n998), 
	.B1(n994), 
	.A(n995));
   INV_X1 U905 (.ZN(n994), 
	.A(n996));
   INV_X1 U906 (.ZN(n995), 
	.A(n997));
   NAND2_X1 U907 (.ZN(n505), 
	.A2(n997), 
	.A1(n994));
   NOR2_X1 U909 (.ZN(n996), 
	.A2(n1999), 
	.A1(n1996));
   NAND2_X1 U910 (.ZN(n997), 
	.A2(n1999), 
	.A1(n1996));
   XOR2_X1 U911 (.Z(product[4]), 
	.B(n1001), 
	.A(n506));
   OAI21_X1 U912 (.ZN(n998), 
	.B2(n1001), 
	.B1(n999), 
	.A(n1000));
   NAND2_X1 U913 (.ZN(n506), 
	.A2(n1000), 
	.A1(n1069));
   INV_X1 U914 (.ZN(n1069), 
	.A(n999));
   NOR2_X1 U915 (.ZN(n999), 
	.A2(n2001), 
	.A1(n2000));
   NAND2_X1 U916 (.ZN(n1000), 
	.A2(n2001), 
	.A1(n2000));
   XNOR2_X1 U917 (.ZN(product[3]), 
	.B(n1006), 
	.A(n507));
   AOI21_X1 U918 (.ZN(n1001), 
	.B2(n1006), 
	.B1(n1002), 
	.A(n1003));
   INV_X1 U919 (.ZN(n1002), 
	.A(n1004));
   INV_X1 U920 (.ZN(n1003), 
	.A(n1005));
   NAND2_X1 U921 (.ZN(n507), 
	.A2(n1005), 
	.A1(n1002));
   NOR2_X1 U923 (.ZN(n1004), 
	.A2(n2017), 
	.A1(n2002));
   NAND2_X1 U924 (.ZN(n1005), 
	.A2(n2017), 
	.A1(n2002));
   XOR2_X1 U925 (.Z(product[2]), 
	.B(n1010), 
	.A(n508));
   OAI21_X1 U926 (.ZN(n1006), 
	.B2(n1010), 
	.B1(n1007), 
	.A(n1008));
   NAND2_X1 U927 (.ZN(n508), 
	.A2(n1008), 
	.A1(n1071));
   INV_X1 U928 (.ZN(n1071), 
	.A(n1007));
   NOR2_X1 U929 (.ZN(n1007), 
	.A2(n2529), 
	.A1(n2498));
   NAND2_X1 U930 (.ZN(n1008), 
	.A2(n2529), 
	.A1(n2498));
   INV_X1 U931 (.ZN(product[1]), 
	.A(n509));
   NAND2_X1 U932 (.ZN(n509), 
	.A2(n1010), 
	.A1(n1072));
   INV_X1 U933 (.ZN(n1072), 
	.A(n1009));
   NOR2_X1 U934 (.ZN(n1009), 
	.A2(n2018), 
	.A1(n2530));
   NAND2_X1 U935 (.ZN(n1010), 
	.A2(n2018), 
	.A1(n2530));
   INV_X1 U936 (.ZN(n1074), 
	.A(n1073));
   FA_X1 U937 (.S(n1076), 
	.CO(n1075), 
	.CI(n2051), 
	.B(n1079), 
	.A(n2020));
   FA_X1 U938 (.S(n1078), 
	.CO(n1077), 
	.CI(n1083), 
	.B(n2021), 
	.A(n1080));
   INV_X1 U939 (.ZN(n1080), 
	.A(n1079));
   FA_X1 U940 (.S(n1082), 
	.CO(n1081), 
	.CI(n1084), 
	.B(n2083), 
	.A(n1087));
   FA_X1 U941 (.S(n1084), 
	.CO(n1083), 
	.CI(n2022), 
	.B(n1089), 
	.A(n2052));
   FA_X1 U942 (.S(n1086), 
	.CO(n1085), 
	.CI(n1093), 
	.B(n1095), 
	.A(n1088));
   FA_X1 U943 (.S(n1088), 
	.CO(n1087), 
	.CI(n1090), 
	.B(n2053), 
	.A(n2023));
   INV_X1 U944 (.ZN(n1090), 
	.A(n1089));
   FA_X1 U945 (.S(n1092), 
	.CO(n1091), 
	.CI(n1094), 
	.B(n1096), 
	.A(n1099));
   FA_X1 U946 (.S(n1094), 
	.CO(n1093), 
	.CI(n1101), 
	.B(n2084), 
	.A(n2115));
   FA_X1 U947 (.S(n1096), 
	.CO(n1095), 
	.CI(n1103), 
	.B(n2024), 
	.A(n2054));
   FA_X1 U948 (.S(n1098), 
	.CO(n1097), 
	.CI(n1107), 
	.B(n1102), 
	.A(n1100));
   FA_X1 U949 (.S(n1100), 
	.CO(n1099), 
	.CI(n1109), 
	.B(n2085), 
	.A(n1111));
   FA_X1 U950 (.S(n1102), 
	.CO(n1101), 
	.CI(n1104), 
	.B(n2025), 
	.A(n2055));
   INV_X1 U951 (.ZN(n1104), 
	.A(n1103));
   FA_X1 U952 (.S(n1106), 
	.CO(n1105), 
	.CI(n1108), 
	.B(n1117), 
	.A(n1115));
   FA_X1 U953 (.S(n1108), 
	.CO(n1107), 
	.CI(n1110), 
	.B(n1119), 
	.A(n1112));
   FA_X1 U954 (.S(n1110), 
	.CO(n1109), 
	.CI(n2147), 
	.B(n2056), 
	.A(n2086));
   FA_X1 U955 (.S(n1112), 
	.CO(n1111), 
	.CI(n1121), 
	.B(n2026), 
	.A(n2116));
   FA_X1 U956 (.S(n1114), 
	.CO(n1113), 
	.CI(n1116), 
	.B(n1118), 
	.A(n1125));
   FA_X1 U957 (.S(n1116), 
	.CO(n1115), 
	.CI(n1127), 
	.B(n1129), 
	.A(n1120));
   FA_X1 U958 (.S(n1118), 
	.CO(n1117), 
	.CI(n1131), 
	.B(n2087), 
	.A(n2027));
   FA_X1 U959 (.S(n1120), 
	.CO(n1119), 
	.CI(n1122), 
	.B(n2057), 
	.A(n2117));
   INV_X1 U960 (.ZN(n1122), 
	.A(n1121));
   FA_X1 U961 (.S(n1124), 
	.CO(n1123), 
	.CI(n1126), 
	.B(n1128), 
	.A(n1135));
   FA_X1 U962 (.S(n1126), 
	.CO(n1125), 
	.CI(n1137), 
	.B(n1130), 
	.A(n1132));
   FA_X1 U963 (.S(n1128), 
	.CO(n1127), 
	.CI(n1139), 
	.B(n2179), 
	.A(n1141));
   FA_X1 U964 (.S(n1130), 
	.CO(n1129), 
	.CI(n2118), 
	.B(n2148), 
	.A(n2058));
   FA_X1 U965 (.S(n1132), 
	.CO(n1131), 
	.CI(n2088), 
	.B(n2028), 
	.A(n1143));
   FA_X1 U966 (.S(n1134), 
	.CO(n1133), 
	.CI(n1136), 
	.B(n1138), 
	.A(n1147));
   FA_X1 U967 (.S(n1136), 
	.CO(n1135), 
	.CI(n1149), 
	.B(n1142), 
	.A(n1151));
   FA_X1 U968 (.S(n1138), 
	.CO(n1137), 
	.CI(n1140), 
	.B(n1155), 
	.A(n1153));
   FA_X1 U969 (.S(n1140), 
	.CO(n1139), 
	.CI(n2119), 
	.B(n2029), 
	.A(n2059));
   FA_X1 U970 (.S(n1142), 
	.CO(n1141), 
	.CI(n1144), 
	.B(n2089), 
	.A(n2149));
   INV_X1 U971 (.ZN(n1144), 
	.A(n1143));
   FA_X1 U972 (.S(n1146), 
	.CO(n1145), 
	.CI(n1148), 
	.B(n1150), 
	.A(n1159));
   FA_X1 U973 (.S(n1148), 
	.CO(n1147), 
	.CI(n1161), 
	.B(n1163), 
	.A(n1152));
   FA_X1 U974 (.S(n1150), 
	.CO(n1149), 
	.CI(n1156), 
	.B(n1165), 
	.A(n1154));
   FA_X1 U975 (.S(n1152), 
	.CO(n1151), 
	.CI(n1167), 
	.B(n2120), 
	.A(n2211));
   FA_X1 U976 (.S(n1154), 
	.CO(n1153), 
	.CI(n2180), 
	.B(n2150), 
	.A(n2090));
   FA_X1 U977 (.S(n1156), 
	.CO(n1155), 
	.CI(n2060), 
	.B(n2030), 
	.A(n1169));
   FA_X1 U978 (.S(n1158), 
	.CO(n1157), 
	.CI(n1160), 
	.B(n1162), 
	.A(n1173));
   FA_X1 U979 (.S(n1160), 
	.CO(n1159), 
	.CI(n1175), 
	.B(n1177), 
	.A(n1164));
   FA_X1 U980 (.S(n1162), 
	.CO(n1161), 
	.CI(n1168), 
	.B(n1179), 
	.A(n1166));
   FA_X1 U981 (.S(n1164), 
	.CO(n1163), 
	.CI(n1181), 
	.B(n2061), 
	.A(n1183));
   FA_X1 U982 (.S(n1166), 
	.CO(n1165), 
	.CI(n2121), 
	.B(n2151), 
	.A(n2031));
   FA_X1 U983 (.S(n1168), 
	.CO(n1167), 
	.CI(n1170), 
	.B(n2091), 
	.A(n2181));
   INV_X1 U984 (.ZN(n1170), 
	.A(n1169));
   FA_X1 U985 (.S(n1172), 
	.CO(n1171), 
	.CI(n1174), 
	.B(n1176), 
	.A(n1187));
   FA_X1 U986 (.S(n1174), 
	.CO(n1173), 
	.CI(n1189), 
	.B(n1191), 
	.A(n1178));
   FA_X1 U987 (.S(n1176), 
	.CO(n1175), 
	.CI(n1193), 
	.B(n1184), 
	.A(n1180));
   FA_X1 U988 (.S(n1178), 
	.CO(n1177), 
	.CI(n1182), 
	.B(n1197), 
	.A(n1195));
   FA_X1 U989 (.S(n1180), 
	.CO(n1179), 
	.CI(n2243), 
	.B(n2062), 
	.A(n2212));
   FA_X1 U990 (.S(n1182), 
	.CO(n1181), 
	.CI(n2152), 
	.B(n2182), 
	.A(n2122));
   FA_X1 U991 (.S(n1184), 
	.CO(n1183), 
	.CI(n2092), 
	.B(n2032), 
	.A(n1199));
   FA_X1 U992 (.S(n1186), 
	.CO(n1185), 
	.CI(n1188), 
	.B(n1190), 
	.A(n1203));
   FA_X1 U993 (.S(n1188), 
	.CO(n1187), 
	.CI(n1205), 
	.B(n1207), 
	.A(n1192));
   FA_X1 U994 (.S(n1190), 
	.CO(n1189), 
	.CI(n1194), 
	.B(n1198), 
	.A(n1209));
   FA_X1 U995 (.S(n1192), 
	.CO(n1191), 
	.CI(n1196), 
	.B(n1213), 
	.A(n1211));
   FA_X1 U996 (.S(n1194), 
	.CO(n1193), 
	.CI(n1215), 
	.B(n2153), 
	.A(n2123));
   FA_X1 U997 (.S(n1196), 
	.CO(n1195), 
	.CI(n2063), 
	.B(n2183), 
	.A(n2033));
   FA_X1 U998 (.S(n1198), 
	.CO(n1197), 
	.CI(n1200), 
	.B(n2093), 
	.A(n2213));
   INV_X1 U999 (.ZN(n1200), 
	.A(n1199));
   FA_X1 U1000 (.S(n1202), 
	.CO(n1201), 
	.CI(n1204), 
	.B(n1206), 
	.A(n1219));
   FA_X1 U1001 (.S(n1204), 
	.CO(n1203), 
	.CI(n1221), 
	.B(n1223), 
	.A(n1208));
   FA_X1 U1002 (.S(n1206), 
	.CO(n1205), 
	.CI(n1210), 
	.B(n1216), 
	.A(n1225));
   FA_X1 U1003 (.S(n1208), 
	.CO(n1207), 
	.CI(n1214), 
	.B(n1227), 
	.A(n1212));
   FA_X1 U1004 (.S(n1210), 
	.CO(n1209), 
	.CI(n1229), 
	.B(n2275), 
	.A(n1231));
   FA_X1 U1005 (.S(n1212), 
	.CO(n1211), 
	.CI(n2214), 
	.B(n2094), 
	.A(n2184));
   FA_X1 U1006 (.S(n1214), 
	.CO(n1213), 
	.CI(n2124), 
	.B(n2154), 
	.A(n2064));
   FA_X1 U1007 (.S(n1216), 
	.CO(n1215), 
	.CI(n1233), 
	.B(n2034), 
	.A(n2244));
   FA_X1 U1008 (.S(n1218), 
	.CO(n1217), 
	.CI(n1220), 
	.B(n1222), 
	.A(n1237));
   FA_X1 U1009 (.S(n1220), 
	.CO(n1219), 
	.CI(n1239), 
	.B(n1241), 
	.A(n1224));
   FA_X1 U1010 (.S(n1222), 
	.CO(n1221), 
	.CI(n1226), 
	.B(n1245), 
	.A(n1243));
   FA_X1 U1011 (.S(n1224), 
	.CO(n1223), 
	.CI(n1230), 
	.B(n1228), 
	.A(n1232));
   FA_X1 U1012 (.S(n1226), 
	.CO(n1225), 
	.CI(n1249), 
	.B(n1251), 
	.A(n1247));
   FA_X1 U1013 (.S(n1228), 
	.CO(n1227), 
	.CI(n2155), 
	.B(n2185), 
	.A(n2095));
   FA_X1 U1014 (.S(n1230), 
	.CO(n1229), 
	.CI(n2215), 
	.B(n2245), 
	.A(n2065));
   FA_X1 U1015 (.S(n1232), 
	.CO(n1231), 
	.CI(n1234), 
	.B(n2125), 
	.A(n2035));
   INV_X1 U1016 (.ZN(n1234), 
	.A(n1233));
   FA_X1 U1017 (.S(n1236), 
	.CO(n1235), 
	.CI(n1238), 
	.B(n1240), 
	.A(n1255));
   FA_X1 U1018 (.S(n1238), 
	.CO(n1237), 
	.CI(n1257), 
	.B(n1259), 
	.A(n1242));
   FA_X1 U1019 (.S(n1240), 
	.CO(n1239), 
	.CI(n1244), 
	.B(n1261), 
	.A(n1246));
   FA_X1 U1020 (.S(n1242), 
	.CO(n1241), 
	.CI(n1263), 
	.B(n1250), 
	.A(n1252));
   FA_X1 U1021 (.S(n1244), 
	.CO(n1243), 
	.CI(n1248), 
	.B(n1267), 
	.A(n1265));
   FA_X1 U1022 (.S(n1246), 
	.CO(n1245), 
	.CI(n1269), 
	.B(n2246), 
	.A(n2307));
   FA_X1 U1023 (.S(n1248), 
	.CO(n1247), 
	.CI(n2156), 
	.B(n2126), 
	.A(n2216));
   FA_X1 U1024 (.S(n1250), 
	.CO(n1249), 
	.CI(n1271), 
	.B(n2186), 
	.A(n2096));
   FA_X1 U1025 (.S(n1252), 
	.CO(n1251), 
	.CI(n2066), 
	.B(n2036), 
	.A(n2276));
   FA_X1 U1026 (.S(n1254), 
	.CO(n1253), 
	.CI(n1256), 
	.B(n1258), 
	.A(n1275));
   FA_X1 U1027 (.S(n1256), 
	.CO(n1255), 
	.CI(n1277), 
	.B(n1279), 
	.A(n1260));
   FA_X1 U1028 (.S(n1258), 
	.CO(n1257), 
	.CI(n1262), 
	.B(n1264), 
	.A(n1281));
   FA_X1 U1029 (.S(n1260), 
	.CO(n1259), 
	.CI(n1283), 
	.B(n1268), 
	.A(n1270));
   FA_X1 U1030 (.S(n1262), 
	.CO(n1261), 
	.CI(n1266), 
	.B(n1287), 
	.A(n1285));
   FA_X1 U1031 (.S(n1264), 
	.CO(n1263), 
	.CI(n1289), 
	.B(n2187), 
	.A(n1291));
   FA_X1 U1032 (.S(n1266), 
	.CO(n1265), 
	.CI(n2157), 
	.B(n2217), 
	.A(n2097));
   FA_X1 U1033 (.S(n1268), 
	.CO(n1267), 
	.CI(n2067), 
	.B(n2247), 
	.A(n2037));
   FA_X1 U1034 (.S(n1270), 
	.CO(n1269), 
	.CI(n1272), 
	.B(n2127), 
	.A(n2277));
   INV_X1 U1035 (.ZN(n1272), 
	.A(n1271));
   FA_X1 U1036 (.S(n1274), 
	.CO(n1273), 
	.CI(n1276), 
	.B(n1278), 
	.A(n1295));
   FA_X1 U1037 (.S(n1276), 
	.CO(n1275), 
	.CI(n1297), 
	.B(n1299), 
	.A(n1280));
   FA_X1 U1038 (.S(n1278), 
	.CO(n1277), 
	.CI(n1282), 
	.B(n1301), 
	.A(n1284));
   FA_X1 U1039 (.S(n1280), 
	.CO(n1279), 
	.CI(n1303), 
	.B(n1286), 
	.A(n1305));
   FA_X1 U1040 (.S(n1282), 
	.CO(n1281), 
	.CI(n1290), 
	.B(n1288), 
	.A(n1292));
   FA_X1 U1041 (.S(n1284), 
	.CO(n1283), 
	.CI(n1309), 
	.B(n1311), 
	.A(n1307));
   FA_X1 U1042 (.S(n1286), 
	.CO(n1285), 
	.CI(n2339), 
	.B(n2278), 
	.A(n2248));
   FA_X1 U1043 (.S(n1288), 
	.CO(n1287), 
	.CI(n2158), 
	.B(n2098), 
	.A(n2218));
   FA_X1 U1044 (.S(n1290), 
	.CO(n1289), 
	.CI(n2128), 
	.B(n2188), 
	.A(n1313));
   FA_X1 U1045 (.S(n1292), 
	.CO(n1291), 
	.CI(n2068), 
	.B(n2038), 
	.A(n2308));
   FA_X1 U1046 (.S(n1294), 
	.CO(n1293), 
	.CI(n1296), 
	.B(n1298), 
	.A(n1317));
   FA_X1 U1047 (.S(n1296), 
	.CO(n1295), 
	.CI(n1319), 
	.B(n1321), 
	.A(n1300));
   FA_X1 U1048 (.S(n1298), 
	.CO(n1297), 
	.CI(n1302), 
	.B(n1323), 
	.A(n1304));
   FA_X1 U1049 (.S(n1300), 
	.CO(n1299), 
	.CI(n1306), 
	.B(n1327), 
	.A(n1325));
   FA_X1 U1050 (.S(n1302), 
	.CO(n1301), 
	.CI(n1310), 
	.B(n1308), 
	.A(n1312));
   FA_X1 U1051 (.S(n1304), 
	.CO(n1303), 
	.CI(n1331), 
	.B(n1333), 
	.A(n1329));
   FA_X1 U1052 (.S(n1306), 
	.CO(n1305), 
	.CI(n1335), 
	.B(n2279), 
	.A(n2249));
   FA_X1 U1053 (.S(n1308), 
	.CO(n1307), 
	.CI(n2189), 
	.B(n2219), 
	.A(n2129));
   FA_X1 U1054 (.S(n1310), 
	.CO(n1309), 
	.CI(n2099), 
	.B(n2309), 
	.A(n2069));
   FA_X1 U1055 (.S(n1312), 
	.CO(n1311), 
	.CI(n1314), 
	.B(n2159), 
	.A(n2039));
   INV_X1 U1056 (.ZN(n1314), 
	.A(n1313));
   FA_X1 U1057 (.S(n1316), 
	.CO(n1315), 
	.CI(n1318), 
	.B(n1320), 
	.A(n1339));
   FA_X1 U1058 (.S(n1318), 
	.CO(n1317), 
	.CI(n1341), 
	.B(n1343), 
	.A(n1322));
   FA_X1 U1059 (.S(n1320), 
	.CO(n1319), 
	.CI(n1324), 
	.B(n1326), 
	.A(n1345));
   FA_X1 U1060 (.S(n1322), 
	.CO(n1321), 
	.CI(n1347), 
	.B(n1349), 
	.A(n1328));
   FA_X1 U1061 (.S(n1324), 
	.CO(n1323), 
	.CI(n1334), 
	.B(n1332), 
	.A(n1336));
   FA_X1 U1062 (.S(n1326), 
	.CO(n1325), 
	.CI(n1330), 
	.B(n1353), 
	.A(n1351));
   FA_X1 U1063 (.S(n1328), 
	.CO(n1327), 
	.CI(n1355), 
	.B(n2371), 
	.A(n1357));
   FA_X1 U1064 (.S(n1330), 
	.CO(n1329), 
	.CI(n2310), 
	.B(n2340), 
	.A(n2190));
   FA_X1 U1065 (.S(n1332), 
	.CO(n1331), 
	.CI(n2250), 
	.B(n2280), 
	.A(n2160));
   FA_X1 U1066 (.S(n1334), 
	.CO(n1333), 
	.CI(n2070), 
	.B(n2220), 
	.A(n2130));
   FA_X1 U1067 (.S(n1336), 
	.CO(n1335), 
	.CI(n2100), 
	.B(n2040), 
	.A(n1359));
   FA_X1 U1068 (.S(n1338), 
	.CO(n1337), 
	.CI(n1340), 
	.B(n1342), 
	.A(n1363));
   FA_X1 U1069 (.S(n1340), 
	.CO(n1339), 
	.CI(n1365), 
	.B(n1367), 
	.A(n1344));
   FA_X1 U1070 (.S(n1342), 
	.CO(n1341), 
	.CI(n1346), 
	.B(n1348), 
	.A(n1369));
   FA_X1 U1071 (.S(n1344), 
	.CO(n1343), 
	.CI(n1350), 
	.B(n1373), 
	.A(n1371));
   FA_X1 U1072 (.S(n1346), 
	.CO(n1345), 
	.CI(n1375), 
	.B(n1356), 
	.A(n1358));
   FA_X1 U1073 (.S(n1348), 
	.CO(n1347), 
	.CI(n1354), 
	.B(n1381), 
	.A(n1352));
   FA_X1 U1074 (.S(n1350), 
	.CO(n1349), 
	.CI(n1379), 
	.B(n1383), 
	.A(n1377));
   FA_X1 U1075 (.S(n1352), 
	.CO(n1351), 
	.CI(n2251), 
	.B(n2281), 
	.A(n2221));
   FA_X1 U1076 (.S(n1354), 
	.CO(n1353), 
	.CI(n2161), 
	.B(n2131), 
	.A(n2311));
   FA_X1 U1077 (.S(n1356), 
	.CO(n1355), 
	.CI(n2101), 
	.B(n2341), 
	.A(n2071));
   FA_X1 U1078 (.S(n1358), 
	.CO(n1357), 
	.CI(n1360), 
	.B(n2191), 
	.A(n2041));
   INV_X1 U1079 (.ZN(n1360), 
	.A(n1359));
   FA_X1 U1080 (.S(n1362), 
	.CO(n1361), 
	.CI(n1364), 
	.B(n1366), 
	.A(n1387));
   FA_X1 U1081 (.S(n1364), 
	.CO(n1363), 
	.CI(n1389), 
	.B(n1391), 
	.A(n1368));
   FA_X1 U1082 (.S(n1366), 
	.CO(n1365), 
	.CI(n1370), 
	.B(n1372), 
	.A(n1393));
   FA_X1 U1083 (.S(n1368), 
	.CO(n1367), 
	.CI(n1374), 
	.B(n1376), 
	.A(n1395));
   FA_X1 U1084 (.S(n1370), 
	.CO(n1369), 
	.CI(n1397), 
	.B(n1380), 
	.A(n1399));
   FA_X1 U1085 (.S(n1372), 
	.CO(n1371), 
	.CI(n1382), 
	.B(n1378), 
	.A(n1384));
   FA_X1 U1086 (.S(n1374), 
	.CO(n1373), 
	.CI(n1405), 
	.B(n1401), 
	.A(n1403));
   FA_X1 U1087 (.S(n1376), 
	.CO(n1375), 
	.CI(n1407), 
	.B(n2342), 
	.A(n2403));
   FA_X1 U1088 (.S(n1378), 
	.CO(n1377), 
	.CI(n2282), 
	.B(n2312), 
	.A(n2072));
   FA_X1 U1089 (.S(n1380), 
	.CO(n1379), 
	.CI(n2192), 
	.B(n2252), 
	.A(n2162));
   FA_X1 U1090 (.S(n1382), 
	.CO(n1381), 
	.CI(n2132), 
	.B(n2222), 
	.A(n2102));
   FA_X1 U1091 (.S(n1384), 
	.CO(n1383), 
	.CI(n1409), 
	.B(n2042), 
	.A(n2372));
   FA_X1 U1092 (.S(n1386), 
	.CO(n1385), 
	.CI(n1388), 
	.B(n1390), 
	.A(n1413));
   FA_X1 U1093 (.S(n1388), 
	.CO(n1387), 
	.CI(n1415), 
	.B(n1417), 
	.A(n1392));
   FA_X1 U1094 (.S(n1390), 
	.CO(n1389), 
	.CI(n1394), 
	.B(n1396), 
	.A(n1419));
   FA_X1 U1095 (.S(n1392), 
	.CO(n1391), 
	.CI(n1421), 
	.B(n1423), 
	.A(n1398));
   FA_X1 U1096 (.S(n1394), 
	.CO(n1393), 
	.CI(n1400), 
	.B(n1404), 
	.A(n1425));
   FA_X1 U1097 (.S(n1396), 
	.CO(n1395), 
	.CI(n1406), 
	.B(n1402), 
	.A(n1408));
   FA_X1 U1098 (.S(n1398), 
	.CO(n1397), 
	.CI(n1427), 
	.B(n1431), 
	.A(n1429));
   FA_X1 U1099 (.S(n1400), 
	.CO(n1399), 
	.CI(n1433), 
	.B(n2253), 
	.A(n1435));
   FA_X1 U1100 (.S(n1402), 
	.CO(n1401), 
	.CI(n2223), 
	.B(n2283), 
	.A(n2163));
   FA_X1 U1101 (.S(n1404), 
	.CO(n1403), 
	.CI(n2133), 
	.B(n2313), 
	.A(n2103));
   FA_X1 U1102 (.S(n1406), 
	.CO(n1405), 
	.CI(n2073), 
	.B(n2343), 
	.A(n2043));
   FA_X1 U1103 (.S(n1408), 
	.CO(n1407), 
	.CI(n1410), 
	.B(n2193), 
	.A(n2373));
   INV_X1 U1104 (.ZN(n1410), 
	.A(n1409));
   FA_X1 U1105 (.S(n1412), 
	.CO(n1411), 
	.CI(n1414), 
	.B(n1416), 
	.A(n1439));
   FA_X1 U1106 (.S(n1414), 
	.CO(n1413), 
	.CI(n1441), 
	.B(n1443), 
	.A(n1418));
   FA_X1 U1107 (.S(n1416), 
	.CO(n1415), 
	.CI(n1420), 
	.B(n1422), 
	.A(n1445));
   FA_X1 U1108 (.S(n1418), 
	.CO(n1417), 
	.CI(n1447), 
	.B(n1426), 
	.A(n1424));
   FA_X1 U1109 (.S(n1420), 
	.CO(n1419), 
	.CI(n1449), 
	.B(n1453), 
	.A(n1451));
   FA_X1 U1110 (.S(n1422), 
	.CO(n1421), 
	.CI(n1428), 
	.B(n1434), 
	.A(n1436));
   FA_X1 U1111 (.S(n1424), 
	.CO(n1423), 
	.CI(n1432), 
	.B(n1455), 
	.A(n1430));
   FA_X1 U1112 (.S(n1426), 
	.CO(n1425), 
	.CI(n1459), 
	.B(n1457), 
	.A(n1461));
   FA_X1 U1113 (.S(n1428), 
	.CO(n1427), 
	.CI(n2435), 
	.B(n2374), 
	.A(n2344));
   FA_X1 U1114 (.S(n1430), 
	.CO(n1429), 
	.CI(n2224), 
	.B(n2194), 
	.A(n2314));
   FA_X1 U1115 (.S(n1432), 
	.CO(n1431), 
	.CI(n2164), 
	.B(n2284), 
	.A(n1463));
   FA_X1 U1116 (.S(n1434), 
	.CO(n1433), 
	.CI(n2134), 
	.B(n2254), 
	.A(n2104));
   FA_X1 U1117 (.S(n1436), 
	.CO(n1435), 
	.CI(n2074), 
	.B(n2044), 
	.A(n2404));
   FA_X1 U1118 (.S(n1438), 
	.CO(n1437), 
	.CI(n1440), 
	.B(n1442), 
	.A(n1467));
   FA_X1 U1119 (.S(n1440), 
	.CO(n1439), 
	.CI(n1469), 
	.B(n1471), 
	.A(n1444));
   FA_X1 U1120 (.S(n1442), 
	.CO(n1441), 
	.CI(n1446), 
	.B(n1448), 
	.A(n1473));
   FA_X1 U1121 (.S(n1444), 
	.CO(n1443), 
	.CI(n1475), 
	.B(n1452), 
	.A(n1450));
   FA_X1 U1122 (.S(n1446), 
	.CO(n1445), 
	.CI(n1477), 
	.B(n1479), 
	.A(n1454));
   FA_X1 U1123 (.S(n1448), 
	.CO(n1447), 
	.CI(n1481), 
	.B(n1462), 
	.A(n1460));
   FA_X1 U1124 (.S(n1450), 
	.CO(n1449), 
	.CI(n1458), 
	.B(n1487), 
	.A(n1456));
   FA_X1 U1125 (.S(n1452), 
	.CO(n1451), 
	.CI(n1483), 
	.B(n1485), 
	.A(n1489));
   FA_X1 U1126 (.S(n1454), 
	.CO(n1453), 
	.CI(n1491), 
	.B(n2315), 
	.A(n2285));
   FA_X1 U1127 (.S(n1456), 
	.CO(n1455), 
	.CI(n2195), 
	.B(n2345), 
	.A(n2165));
   FA_X1 U1128 (.S(n1458), 
	.CO(n1457), 
	.CI(n2375), 
	.B(n2405), 
	.A(n2135));
   FA_X1 U1129 (.S(n1460), 
	.CO(n1459), 
	.CI(n2105), 
	.B(n2255), 
	.A(n2075));
   FA_X1 U1130 (.S(n1462), 
	.CO(n1461), 
	.CI(n1464), 
	.B(n2225), 
	.A(n2045));
   INV_X1 U1131 (.ZN(n1464), 
	.A(n1463));
   FA_X1 U1132 (.S(n1466), 
	.CO(n1465), 
	.CI(n1468), 
	.B(n1470), 
	.A(n1495));
   FA_X1 U1133 (.S(n1468), 
	.CO(n1467), 
	.CI(n1497), 
	.B(n1499), 
	.A(n1472));
   FA_X1 U1134 (.S(n1470), 
	.CO(n1469), 
	.CI(n1474), 
	.B(n1476), 
	.A(n1501));
   FA_X1 U1135 (.S(n1472), 
	.CO(n1471), 
	.CI(n1478), 
	.B(n1480), 
	.A(n1503));
   FA_X1 U1136 (.S(n1474), 
	.CO(n1473), 
	.CI(n1505), 
	.B(n1507), 
	.A(n1482));
   FA_X1 U1137 (.S(n1476), 
	.CO(n1475), 
	.CI(n1509), 
	.B(n1488), 
	.A(n1486));
   FA_X1 U1138 (.S(n1478), 
	.CO(n1477), 
	.CI(n1490), 
	.B(n1484), 
	.A(n1492));
   FA_X1 U1139 (.S(n1480), 
	.CO(n1479), 
	.CI(n1513), 
	.B(n1511), 
	.A(n1515));
   FA_X1 U1140 (.S(n1482), 
	.CO(n1481), 
	.CI(n1517), 
	.B(n2467), 
	.A(n1519));
   FA_X1 U1141 (.S(n1484), 
	.CO(n1483), 
	.CI(n2256), 
	.B(n2406), 
	.A(n2436));
   FA_X1 U1142 (.S(n1486), 
	.CO(n1485), 
	.CI(n2376), 
	.B(n2226), 
	.A(n2346));
   FA_X1 U1143 (.S(n1488), 
	.CO(n1487), 
	.CI(n2136), 
	.B(n2316), 
	.A(n2196));
   FA_X1 U1144 (.S(n1490), 
	.CO(n1489), 
	.CI(n2166), 
	.B(n2286), 
	.A(n2106));
   FA_X1 U1145 (.S(n1492), 
	.CO(n1491), 
	.CI(n2076), 
	.B(n2046), 
	.A(n1521));
   FA_X1 U1146 (.S(n1494), 
	.CO(n1493), 
	.CI(n1496), 
	.B(n1498), 
	.A(n1525));
   FA_X1 U1147 (.S(n1496), 
	.CO(n1495), 
	.CI(n1527), 
	.B(n1502), 
	.A(n1500));
   FA_X1 U1148 (.S(n1498), 
	.CO(n1497), 
	.CI(n1529), 
	.B(n1504), 
	.A(n1531));
   FA_X1 U1149 (.S(n1500), 
	.CO(n1499), 
	.CI(n1506), 
	.B(n1508), 
	.A(n1533));
   FA_X1 U1150 (.S(n1502), 
	.CO(n1501), 
	.CI(n1535), 
	.B(n1537), 
	.A(n1510));
   FA_X1 U1151 (.S(n1504), 
	.CO(n1503), 
	.CI(n1539), 
	.B(n1514), 
	.A(n1516));
   FA_X1 U1152 (.S(n1506), 
	.CO(n1505), 
	.CI(n1518), 
	.B(n1512), 
	.A(n1520));
   FA_X1 U1153 (.S(n1508), 
	.CO(n1507), 
	.CI(n1541), 
	.B(n1545), 
	.A(n1543));
   FA_X1 U1154 (.S(n1510), 
	.CO(n1509), 
	.CI(n1547), 
	.B(n1551), 
	.A(n1549));
   FA_X1 U1155 (.S(n1512), 
	.CO(n1511), 
	.CI(n2317), 
	.B(n2347), 
	.A(n2287));
   FA_X1 U1156 (.S(n1514), 
	.CO(n1513), 
	.CI(n2197), 
	.B(n2377), 
	.A(n2167));
   FA_X1 U1157 (.S(n1516), 
	.CO(n1515), 
	.CI(n2137), 
	.B(n2407), 
	.A(n2107));
   FA_X1 U1158 (.S(n1518), 
	.CO(n1517), 
	.CI(n2077), 
	.B(n2257), 
	.A(n2437));
   FA_X1 U1159 (.S(n1520), 
	.CO(n1519), 
	.CI(n1522), 
	.B(n2227), 
	.A(n2047));
   INV_X1 U1160 (.ZN(n1522), 
	.A(n1521));
   FA_X1 U1161 (.S(n1524), 
	.CO(n1523), 
	.CI(n1526), 
	.B(n1528), 
	.A(n1555));
   FA_X1 U1162 (.S(n1526), 
	.CO(n1525), 
	.CI(n1557), 
	.B(n1532), 
	.A(n1530));
   FA_X1 U1163 (.S(n1528), 
	.CO(n1527), 
	.CI(n1559), 
	.B(n1534), 
	.A(n1561));
   FA_X1 U1164 (.S(n1530), 
	.CO(n1529), 
	.CI(n1536), 
	.B(n1538), 
	.A(n1563));
   FA_X1 U1165 (.S(n1532), 
	.CO(n1531), 
	.CI(n1565), 
	.B(n1567), 
	.A(n1540));
   FA_X1 U1166 (.S(n1534), 
	.CO(n1533), 
	.CI(n1569), 
	.B(n1546), 
	.A(n1542));
   FA_X1 U1167 (.S(n1536), 
	.CO(n1535), 
	.CI(n1544), 
	.B(n1548), 
	.A(n1550));
   FA_X1 U1168 (.S(n1538), 
	.CO(n1537), 
	.CI(n1577), 
	.B(n1571), 
	.A(n1579));
   FA_X1 U1169 (.S(n1540), 
	.CO(n1539), 
	.CI(n1575), 
	.B(n1552), 
	.A(n1573));
   FA_X1 U1170 (.S(n1542), 
	.CO(n1541), 
	.CI(n1581), 
	.B(n2408), 
	.A(n2499));
   FA_X1 U1171 (.S(n1544), 
	.CO(n1543), 
	.CI(n2468), 
	.B(n2438), 
	.A(n2378));
   FA_X1 U1172 (.S(n1546), 
	.CO(n1545), 
	.CI(n2228), 
	.B(n2348), 
	.A(n2198));
   FA_X1 U1173 (.S(n1548), 
	.CO(n1547), 
	.CI(n2168), 
	.B(n2288), 
	.A(n2138));
   FA_X1 U1174 (.S(n1550), 
	.CO(n1549), 
	.CI(n2108), 
	.B(n2258), 
	.A(n2048));
   XNOR2_X1 U1175 (.ZN(n1552), 
	.B(n2078), 
	.A(n2318));
   OR2_X1 U1176 (.ZN(n1551), 
	.A2(n2078), 
	.A1(n2318));
   FA_X1 U1177 (.S(n1554), 
	.CO(n1553), 
	.CI(n1556), 
	.B(n1558), 
	.A(n1585));
   FA_X1 U1178 (.S(n1556), 
	.CO(n1555), 
	.CI(n1587), 
	.B(n1562), 
	.A(n1560));
   FA_X1 U1179 (.S(n1558), 
	.CO(n1557), 
	.CI(n1589), 
	.B(n1564), 
	.A(n1591));
   FA_X1 U1180 (.S(n1560), 
	.CO(n1559), 
	.CI(n1566), 
	.B(n1568), 
	.A(n1593));
   FA_X1 U1181 (.S(n1562), 
	.CO(n1561), 
	.CI(n1595), 
	.B(n1597), 
	.A(n1570));
   FA_X1 U1182 (.S(n1564), 
	.CO(n1563), 
	.CI(n1599), 
	.B(n1576), 
	.A(n1574));
   FA_X1 U1183 (.S(n1566), 
	.CO(n1565), 
	.CI(n1578), 
	.B(n1572), 
	.A(n1580));
   FA_X1 U1184 (.S(n1568), 
	.CO(n1567), 
	.CI(n1603), 
	.B(n1601), 
	.A(n1605));
   FA_X1 U1185 (.S(n1570), 
	.CO(n1569), 
	.CI(n1607), 
	.B(n1582), 
	.A(n1609));
   FA_X1 U1186 (.S(n1572), 
	.CO(n1571), 
	.CI(n2259), 
	.B(n2199), 
	.A(n2319));
   FA_X1 U1187 (.S(n1574), 
	.CO(n1573), 
	.CI(n2139), 
	.B(n2349), 
	.A(n2109));
   FA_X1 U1188 (.S(n1576), 
	.CO(n1575), 
	.CI(n2379), 
	.B(n2169), 
	.A(n2079));
   FA_X1 U1189 (.S(n1578), 
	.CO(n1577), 
	.CI(n2409), 
	.B(n2229), 
	.A(n2439));
   FA_X1 U1190 (.S(n1580), 
	.CO(n1579), 
	.CI(n2469), 
	.B(n2289), 
	.A(n2500));
   HA_X1 U1191 (.S(n1582), 
	.CO(n1581), 
	.B(n2003), 
	.A(n2049));
   FA_X1 U1192 (.S(n1584), 
	.CO(n1583), 
	.CI(n1586), 
	.B(n1588), 
	.A(n1613));
   FA_X1 U1193 (.S(n1586), 
	.CO(n1585), 
	.CI(n1615), 
	.B(n1592), 
	.A(n1590));
   FA_X1 U1194 (.S(n1588), 
	.CO(n1587), 
	.CI(n1617), 
	.B(n1594), 
	.A(n1619));
   FA_X1 U1195 (.S(n1590), 
	.CO(n1589), 
	.CI(n1596), 
	.B(n1621), 
	.A(n1598));
   FA_X1 U1196 (.S(n1592), 
	.CO(n1591), 
	.CI(n1600), 
	.B(n1625), 
	.A(n1623));
   FA_X1 U1197 (.S(n1594), 
	.CO(n1593), 
	.CI(n1627), 
	.B(n1604), 
	.A(n1606));
   FA_X1 U1198 (.S(n1596), 
	.CO(n1595), 
	.CI(n1608), 
	.B(n1602), 
	.A(n1610));
   FA_X1 U1199 (.S(n1598), 
	.CO(n1597), 
	.CI(n1631), 
	.B(n1629), 
	.A(n1633));
   FA_X1 U1200 (.S(n1600), 
	.CO(n1599), 
	.CI(n1635), 
	.B(n2350), 
	.A(n1637));
   FA_X1 U1201 (.S(n1602), 
	.CO(n1601), 
	.CI(n2320), 
	.B(n2380), 
	.A(n2290));
   FA_X1 U1202 (.S(n1604), 
	.CO(n1603), 
	.CI(n2260), 
	.B(n2200), 
	.A(n2230));
   FA_X1 U1203 (.S(n1606), 
	.CO(n1605), 
	.CI(n2170), 
	.B(n2410), 
	.A(n2140));
   FA_X1 U1204 (.S(n1608), 
	.CO(n1607), 
	.CI(n2440), 
	.B(n2470), 
	.A(n2110));
   FA_X1 U1205 (.S(n1610), 
	.CO(n1609), 
	.CI(n2050), 
	.B(n2501), 
	.A(n2080));
   FA_X1 U1206 (.S(n1612), 
	.CO(n1611), 
	.CI(n1614), 
	.B(n1616), 
	.A(n1641));
   FA_X1 U1207 (.S(n1614), 
	.CO(n1613), 
	.CI(n1643), 
	.B(n1620), 
	.A(n1618));
   FA_X1 U1208 (.S(n1616), 
	.CO(n1615), 
	.CI(n1645), 
	.B(n1622), 
	.A(n1647));
   FA_X1 U1209 (.S(n1618), 
	.CO(n1617), 
	.CI(n1624), 
	.B(n1649), 
	.A(n1626));
   FA_X1 U1210 (.S(n1620), 
	.CO(n1619), 
	.CI(n1651), 
	.B(n1653), 
	.A(n1628));
   FA_X1 U1211 (.S(n1622), 
	.CO(n1621), 
	.CI(n1636), 
	.B(n1634), 
	.A(n1632));
   FA_X1 U1212 (.S(n1624), 
	.CO(n1623), 
	.CI(n1630), 
	.B(n1659), 
	.A(n1655));
   FA_X1 U1213 (.S(n1626), 
	.CO(n1625), 
	.CI(n1661), 
	.B(n1657), 
	.A(n1663));
   FA_X1 U1214 (.S(n1628), 
	.CO(n1627), 
	.CI(n1638), 
	.B(n2351), 
	.A(n2381));
   FA_X1 U1215 (.S(n1630), 
	.CO(n1629), 
	.CI(n2231), 
	.B(n2411), 
	.A(n2201));
   FA_X1 U1216 (.S(n1632), 
	.CO(n1631), 
	.CI(n2171), 
	.B(n2321), 
	.A(n2441));
   FA_X1 U1217 (.S(n1634), 
	.CO(n1633), 
	.CI(n2141), 
	.B(n2261), 
	.A(n2471));
   FA_X1 U1218 (.S(n1636), 
	.CO(n1635), 
	.CI(n2111), 
	.B(n2291), 
	.A(n2502));
   HA_X1 U1219 (.S(n1638), 
	.CO(n1637), 
	.B(n2004), 
	.A(n2081));
   FA_X1 U1220 (.S(n1640), 
	.CO(n1639), 
	.CI(n1642), 
	.B(n1644), 
	.A(n1667));
   FA_X1 U1221 (.S(n1642), 
	.CO(n1641), 
	.CI(n1669), 
	.B(n1671), 
	.A(n1646));
   FA_X1 U1222 (.S(n1644), 
	.CO(n1643), 
	.CI(n1648), 
	.B(n1650), 
	.A(n1673));
   FA_X1 U1223 (.S(n1646), 
	.CO(n1645), 
	.CI(n1652), 
	.B(n1654), 
	.A(n1675));
   FA_X1 U1224 (.S(n1648), 
	.CO(n1647), 
	.CI(n1677), 
	.B(n1660), 
	.A(n1679));
   FA_X1 U1225 (.S(n1650), 
	.CO(n1649), 
	.CI(n1662), 
	.B(n1658), 
	.A(n1664));
   FA_X1 U1226 (.S(n1652), 
	.CO(n1651), 
	.CI(n1656), 
	.B(n1681), 
	.A(n1683));
   FA_X1 U1227 (.S(n1654), 
	.CO(n1653), 
	.CI(n1685), 
	.B(n1689), 
	.A(n1687));
   FA_X1 U1228 (.S(n1656), 
	.CO(n1655), 
	.CI(n2322), 
	.B(n2352), 
	.A(n2292));
   FA_X1 U1229 (.S(n1658), 
	.CO(n1657), 
	.CI(n2262), 
	.B(n2382), 
	.A(n2232));
   FA_X1 U1230 (.S(n1660), 
	.CO(n1659), 
	.CI(n2202), 
	.B(n2412), 
	.A(n2172));
   FA_X1 U1231 (.S(n1662), 
	.CO(n1661), 
	.CI(n2442), 
	.B(n2472), 
	.A(n2142));
   FA_X1 U1232 (.S(n1664), 
	.CO(n1663), 
	.CI(n2082), 
	.B(n2503), 
	.A(n2112));
   FA_X1 U1233 (.S(n1666), 
	.CO(n1665), 
	.CI(n1668), 
	.B(n1670), 
	.A(n1693));
   FA_X1 U1234 (.S(n1668), 
	.CO(n1667), 
	.CI(n1695), 
	.B(n1674), 
	.A(n1672));
   FA_X1 U1235 (.S(n1670), 
	.CO(n1669), 
	.CI(n1697), 
	.B(n1699), 
	.A(n1676));
   FA_X1 U1236 (.S(n1672), 
	.CO(n1671), 
	.CI(n1678), 
	.B(n1680), 
	.A(n1701));
   FA_X1 U1237 (.S(n1674), 
	.CO(n1673), 
	.CI(n1703), 
	.B(n1688), 
	.A(n1686));
   FA_X1 U1238 (.S(n1676), 
	.CO(n1675), 
	.CI(n1684), 
	.B(n1705), 
	.A(n1682));
   FA_X1 U1239 (.S(n1678), 
	.CO(n1677), 
	.CI(n1711), 
	.B(n1707), 
	.A(n1709));
   FA_X1 U1240 (.S(n1680), 
	.CO(n1679), 
	.CI(n1713), 
	.B(n2413), 
	.A(n1690));
   FA_X1 U1241 (.S(n1682), 
	.CO(n1681), 
	.CI(n2383), 
	.B(n2443), 
	.A(n2353));
   FA_X1 U1242 (.S(n1684), 
	.CO(n1683), 
	.CI(n2233), 
	.B(n2263), 
	.A(n2473));
   FA_X1 U1243 (.S(n1686), 
	.CO(n1685), 
	.CI(n2203), 
	.B(n2293), 
	.A(n2173));
   FA_X1 U1244 (.S(n1688), 
	.CO(n1687), 
	.CI(n2504), 
	.B(n2323), 
	.A(n2143));
   HA_X1 U1245 (.S(n1690), 
	.CO(n1689), 
	.B(n2005), 
	.A(n2113));
   FA_X1 U1246 (.S(n1692), 
	.CO(n1691), 
	.CI(n1694), 
	.B(n1696), 
	.A(n1717));
   FA_X1 U1247 (.S(n1694), 
	.CO(n1693), 
	.CI(n1698), 
	.B(n1721), 
	.A(n1719));
   FA_X1 U1248 (.S(n1696), 
	.CO(n1695), 
	.CI(n1700), 
	.B(n1704), 
	.A(n1702));
   FA_X1 U1249 (.S(n1698), 
	.CO(n1697), 
	.CI(n1723), 
	.B(n1727), 
	.A(n1725));
   FA_X1 U1250 (.S(n1700), 
	.CO(n1699), 
	.CI(n1706), 
	.B(n1714), 
	.A(n1712));
   FA_X1 U1251 (.S(n1702), 
	.CO(n1701), 
	.CI(n1710), 
	.B(n1735), 
	.A(n1708));
   FA_X1 U1252 (.S(n1704), 
	.CO(n1703), 
	.CI(n1733), 
	.B(n1731), 
	.A(n1729));
   FA_X1 U1253 (.S(n1706), 
	.CO(n1705), 
	.CI(n1737), 
	.B(n2384), 
	.A(n2354));
   FA_X1 U1254 (.S(n1708), 
	.CO(n1707), 
	.CI(n2324), 
	.B(n2414), 
	.A(n2294));
   FA_X1 U1255 (.S(n1710), 
	.CO(n1709), 
	.CI(n2264), 
	.B(n2444), 
	.A(n2234));
   FA_X1 U1256 (.S(n1712), 
	.CO(n1711), 
	.CI(n2204), 
	.B(n2474), 
	.A(n2174));
   FA_X1 U1257 (.S(n1714), 
	.CO(n1713), 
	.CI(n2114), 
	.B(n2505), 
	.A(n2144));
   FA_X1 U1258 (.S(n1716), 
	.CO(n1715), 
	.CI(n1718), 
	.B(n1720), 
	.A(n1741));
   FA_X1 U1259 (.S(n1718), 
	.CO(n1717), 
	.CI(n1743), 
	.B(n1745), 
	.A(n1722));
   FA_X1 U1260 (.S(n1720), 
	.CO(n1719), 
	.CI(n1724), 
	.B(n1747), 
	.A(n1726));
   FA_X1 U1261 (.S(n1722), 
	.CO(n1721), 
	.CI(n1728), 
	.B(n1751), 
	.A(n1749));
   FA_X1 U1262 (.S(n1724), 
	.CO(n1723), 
	.CI(n1734), 
	.B(n1732), 
	.A(n1736));
   FA_X1 U1263 (.S(n1726), 
	.CO(n1725), 
	.CI(n1730), 
	.B(n1755), 
	.A(n1753));
   FA_X1 U1264 (.S(n1728), 
	.CO(n1727), 
	.CI(n1757), 
	.B(n1738), 
	.A(n1759));
   FA_X1 U1265 (.S(n1730), 
	.CO(n1729), 
	.CI(n2355), 
	.B(n2385), 
	.A(n2265));
   FA_X1 U1266 (.S(n1732), 
	.CO(n1731), 
	.CI(n2235), 
	.B(n2415), 
	.A(n2205));
   FA_X1 U1267 (.S(n1734), 
	.CO(n1733), 
	.CI(n2445), 
	.B(n2295), 
	.A(n2475));
   FA_X1 U1268 (.S(n1736), 
	.CO(n1735), 
	.CI(n2175), 
	.B(n2325), 
	.A(n2506));
   HA_X1 U1269 (.S(n1738), 
	.CO(n1737), 
	.B(n2006), 
	.A(n2145));
   FA_X1 U1270 (.S(n1740), 
	.CO(n1739), 
	.CI(n1742), 
	.B(n1744), 
	.A(n1763));
   FA_X1 U1271 (.S(n1742), 
	.CO(n1741), 
	.CI(n1765), 
	.B(n1767), 
	.A(n1746));
   FA_X1 U1272 (.S(n1744), 
	.CO(n1743), 
	.CI(n1748), 
	.B(n1769), 
	.A(n1750));
   FA_X1 U1273 (.S(n1746), 
	.CO(n1745), 
	.CI(n1752), 
	.B(n1773), 
	.A(n1771));
   FA_X1 U1274 (.S(n1748), 
	.CO(n1747), 
	.CI(n1758), 
	.B(n1756), 
	.A(n1760));
   FA_X1 U1275 (.S(n1750), 
	.CO(n1749), 
	.CI(n1754), 
	.B(n1777), 
	.A(n1775));
   FA_X1 U1276 (.S(n1752), 
	.CO(n1751), 
	.CI(n1779), 
	.B(n2356), 
	.A(n1781));
   FA_X1 U1277 (.S(n1754), 
	.CO(n1753), 
	.CI(n2326), 
	.B(n2386), 
	.A(n2296));
   FA_X1 U1278 (.S(n1756), 
	.CO(n1755), 
	.CI(n2416), 
	.B(n2446), 
	.A(n2266));
   FA_X1 U1279 (.S(n1758), 
	.CO(n1757), 
	.CI(n2236), 
	.B(n2476), 
	.A(n2206));
   FA_X1 U1280 (.S(n1760), 
	.CO(n1759), 
	.CI(n2146), 
	.B(n2507), 
	.A(n2176));
   FA_X1 U1281 (.S(n1762), 
	.CO(n1761), 
	.CI(n1764), 
	.B(n1766), 
	.A(n1785));
   FA_X1 U1282 (.S(n1764), 
	.CO(n1763), 
	.CI(n1768), 
	.B(n1770), 
	.A(n1787));
   FA_X1 U1283 (.S(n1766), 
	.CO(n1765), 
	.CI(n1789), 
	.B(n1791), 
	.A(n1772));
   FA_X1 U1284 (.S(n1768), 
	.CO(n1767), 
	.CI(n1774), 
	.B(n1780), 
	.A(n1793));
   FA_X1 U1285 (.S(n1770), 
	.CO(n1769), 
	.CI(n1778), 
	.B(n1799), 
	.A(n1776));
   FA_X1 U1286 (.S(n1772), 
	.CO(n1771), 
	.CI(n1797), 
	.B(n1801), 
	.A(n1795));
   FA_X1 U1287 (.S(n1774), 
	.CO(n1773), 
	.CI(n1782), 
	.B(n2417), 
	.A(n2387));
   FA_X1 U1288 (.S(n1776), 
	.CO(n1775), 
	.CI(n2297), 
	.B(n2447), 
	.A(n2267));
   FA_X1 U1289 (.S(n1778), 
	.CO(n1777), 
	.CI(n2237), 
	.B(n2327), 
	.A(n2477));
   FA_X1 U1290 (.S(n1780), 
	.CO(n1779), 
	.CI(n2207), 
	.B(n2357), 
	.A(n2508));
   HA_X1 U1291 (.S(n1782), 
	.CO(n1781), 
	.B(n2007), 
	.A(n2177));
   FA_X1 U1292 (.S(n1784), 
	.CO(n1783), 
	.CI(n1786), 
	.B(n1788), 
	.A(n1805));
   FA_X1 U1293 (.S(n1786), 
	.CO(n1785), 
	.CI(n1807), 
	.B(n1792), 
	.A(n1790));
   FA_X1 U1294 (.S(n1788), 
	.CO(n1787), 
	.CI(n1809), 
	.B(n1811), 
	.A(n1794));
   FA_X1 U1295 (.S(n1790), 
	.CO(n1789), 
	.CI(n1813), 
	.B(n1800), 
	.A(n1802));
   FA_X1 U1296 (.S(n1792), 
	.CO(n1791), 
	.CI(n1798), 
	.B(n1815), 
	.A(n1796));
   FA_X1 U1297 (.S(n1794), 
	.CO(n1793), 
	.CI(n1817), 
	.B(n1821), 
	.A(n1819));
   FA_X1 U1298 (.S(n1796), 
	.CO(n1795), 
	.CI(n2388), 
	.B(n2418), 
	.A(n2358));
   FA_X1 U1299 (.S(n1798), 
	.CO(n1797), 
	.CI(n2328), 
	.B(n2448), 
	.A(n2298));
   FA_X1 U1300 (.S(n1800), 
	.CO(n1799), 
	.CI(n2268), 
	.B(n2478), 
	.A(n2238));
   FA_X1 U1301 (.S(n1802), 
	.CO(n1801), 
	.CI(n2178), 
	.B(n2509), 
	.A(n2208));
   FA_X1 U1302 (.S(n1804), 
	.CO(n1803), 
	.CI(n1806), 
	.B(n1808), 
	.A(n1825));
   FA_X1 U1303 (.S(n1806), 
	.CO(n1805), 
	.CI(n1827), 
	.B(n1812), 
	.A(n1810));
   FA_X1 U1304 (.S(n1808), 
	.CO(n1807), 
	.CI(n1829), 
	.B(n1831), 
	.A(n1814));
   FA_X1 U1305 (.S(n1810), 
	.CO(n1809), 
	.CI(n1818), 
	.B(n1816), 
	.A(n1820));
   FA_X1 U1306 (.S(n1812), 
	.CO(n1811), 
	.CI(n1833), 
	.B(n1837), 
	.A(n1835));
   FA_X1 U1307 (.S(n1814), 
	.CO(n1813), 
	.CI(n1839), 
	.B(n2389), 
	.A(n1822));
   FA_X1 U1308 (.S(n1816), 
	.CO(n1815), 
	.CI(n2299), 
	.B(n2419), 
	.A(n2269));
   FA_X1 U1309 (.S(n1818), 
	.CO(n1817), 
	.CI(n2449), 
	.B(n2329), 
	.A(n2239));
   FA_X1 U1310 (.S(n1820), 
	.CO(n1819), 
	.CI(n2479), 
	.B(n2359), 
	.A(n2510));
   HA_X1 U1311 (.S(n1822), 
	.CO(n1821), 
	.B(n2008), 
	.A(n2209));
   FA_X1 U1312 (.S(n1824), 
	.CO(n1823), 
	.CI(n1826), 
	.B(n1828), 
	.A(n1843));
   FA_X1 U1313 (.S(n1826), 
	.CO(n1825), 
	.CI(n1845), 
	.B(n1832), 
	.A(n1830));
   FA_X1 U1314 (.S(n1828), 
	.CO(n1827), 
	.CI(n1847), 
	.B(n1834), 
	.A(n1849));
   FA_X1 U1315 (.S(n1830), 
	.CO(n1829), 
	.CI(n1838), 
	.B(n1836), 
	.A(n1840));
   FA_X1 U1316 (.S(n1832), 
	.CO(n1831), 
	.CI(n1853), 
	.B(n1855), 
	.A(n1851));
   FA_X1 U1317 (.S(n1834), 
	.CO(n1833), 
	.CI(n1857), 
	.B(n2420), 
	.A(n2390));
   FA_X1 U1318 (.S(n1836), 
	.CO(n1835), 
	.CI(n2360), 
	.B(n2450), 
	.A(n2330));
   FA_X1 U1319 (.S(n1838), 
	.CO(n1837), 
	.CI(n2300), 
	.B(n2480), 
	.A(n2270));
   FA_X1 U1320 (.S(n1840), 
	.CO(n1839), 
	.CI(n2210), 
	.B(n2511), 
	.A(n2240));
   FA_X1 U1321 (.S(n1842), 
	.CO(n1841), 
	.CI(n1844), 
	.B(n1846), 
	.A(n1861));
   FA_X1 U1322 (.S(n1844), 
	.CO(n1843), 
	.CI(n1863), 
	.B(n1865), 
	.A(n1848));
   FA_X1 U1323 (.S(n1846), 
	.CO(n1845), 
	.CI(n1850), 
	.B(n1856), 
	.A(n1867));
   FA_X1 U1324 (.S(n1848), 
	.CO(n1847), 
	.CI(n1854), 
	.B(n1869), 
	.A(n1852));
   FA_X1 U1325 (.S(n1850), 
	.CO(n1849), 
	.CI(n1871), 
	.B(n1858), 
	.A(n1873));
   FA_X1 U1326 (.S(n1852), 
	.CO(n1851), 
	.CI(n2451), 
	.B(n2481), 
	.A(n2361));
   FA_X1 U1327 (.S(n1854), 
	.CO(n1853), 
	.CI(n2331), 
	.B(n2421), 
	.A(n2512));
   FA_X1 U1328 (.S(n1856), 
	.CO(n1855), 
	.CI(n2301), 
	.B(n2391), 
	.A(n2271));
   HA_X1 U1329 (.S(n1858), 
	.CO(n1857), 
	.B(n2009), 
	.A(n2241));
   FA_X1 U1330 (.S(n1860), 
	.CO(n1859), 
	.CI(n1862), 
	.B(n1864), 
	.A(n1877));
   FA_X1 U1331 (.S(n1862), 
	.CO(n1861), 
	.CI(n1879), 
	.B(n1868), 
	.A(n1866));
   FA_X1 U1332 (.S(n1864), 
	.CO(n1863), 
	.CI(n1881), 
	.B(n1874), 
	.A(n1883));
   FA_X1 U1333 (.S(n1866), 
	.CO(n1865), 
	.CI(n1872), 
	.B(n1885), 
	.A(n1870));
   FA_X1 U1334 (.S(n1868), 
	.CO(n1867), 
	.CI(n1887), 
	.B(n2422), 
	.A(n1889));
   FA_X1 U1335 (.S(n1870), 
	.CO(n1869), 
	.CI(n2392), 
	.B(n2452), 
	.A(n2362));
   FA_X1 U1336 (.S(n1872), 
	.CO(n1871), 
	.CI(n2332), 
	.B(n2482), 
	.A(n2302));
   FA_X1 U1337 (.S(n1874), 
	.CO(n1873), 
	.CI(n2242), 
	.B(n2513), 
	.A(n2272));
   FA_X1 U1338 (.S(n1876), 
	.CO(n1875), 
	.CI(n1878), 
	.B(n1893), 
	.A(n1880));
   FA_X1 U1339 (.S(n1878), 
	.CO(n1877), 
	.CI(n1882), 
	.B(n1884), 
	.A(n1895));
   FA_X1 U1340 (.S(n1880), 
	.CO(n1879), 
	.CI(n1897), 
	.B(n1886), 
	.A(n1888));
   FA_X1 U1341 (.S(n1882), 
	.CO(n1881), 
	.CI(n1901), 
	.B(n1903), 
	.A(n1899));
   FA_X1 U1342 (.S(n1884), 
	.CO(n1883), 
	.CI(n1890), 
	.B(n2483), 
	.A(n2453));
   FA_X1 U1343 (.S(n1886), 
	.CO(n1885), 
	.CI(n2363), 
	.B(n2423), 
	.A(n2333));
   FA_X1 U1344 (.S(n1888), 
	.CO(n1887), 
	.CI(n2514), 
	.B(n2393), 
	.A(n2303));
   HA_X1 U1345 (.S(n1890), 
	.CO(n1889), 
	.B(n2010), 
	.A(n2273));
   FA_X1 U1346 (.S(n1892), 
	.CO(n1891), 
	.CI(n1894), 
	.B(n1896), 
	.A(n1907));
   FA_X1 U1347 (.S(n1894), 
	.CO(n1893), 
	.CI(n1898), 
	.B(n1911), 
	.A(n1909));
   FA_X1 U1348 (.S(n1896), 
	.CO(n1895), 
	.CI(n1900), 
	.B(n1904), 
	.A(n1902));
   FA_X1 U1349 (.S(n1898), 
	.CO(n1897), 
	.CI(n1913), 
	.B(n1917), 
	.A(n1915));
   FA_X1 U1350 (.S(n1900), 
	.CO(n1899), 
	.CI(n2424), 
	.B(n2454), 
	.A(n2394));
   FA_X1 U1351 (.S(n1902), 
	.CO(n1901), 
	.CI(n2364), 
	.B(n2484), 
	.A(n2334));
   FA_X1 U1352 (.S(n1904), 
	.CO(n1903), 
	.CI(n2274), 
	.B(n2515), 
	.A(n2304));
   FA_X1 U1353 (.S(n1906), 
	.CO(n1905), 
	.CI(n1908), 
	.B(n1910), 
	.A(n1921));
   FA_X1 U1354 (.S(n1908), 
	.CO(n1907), 
	.CI(n1912), 
	.B(n1916), 
	.A(n1923));
   FA_X1 U1355 (.S(n1910), 
	.CO(n1909), 
	.CI(n1914), 
	.B(n1927), 
	.A(n1925));
   FA_X1 U1356 (.S(n1912), 
	.CO(n1911), 
	.CI(n1929), 
	.B(n2395), 
	.A(n1918));
   FA_X1 U1357 (.S(n1914), 
	.CO(n1913), 
	.CI(n2365), 
	.B(n2335), 
	.A(n2455));
   FA_X1 U1358 (.S(n1916), 
	.CO(n1915), 
	.CI(n2485), 
	.B(n2425), 
	.A(n2516));
   HA_X1 U1359 (.S(n1918), 
	.CO(n1917), 
	.B(n2011), 
	.A(n2305));
   FA_X1 U1360 (.S(n1920), 
	.CO(n1919), 
	.CI(n1922), 
	.B(n1924), 
	.A(n1933));
   FA_X1 U1361 (.S(n1922), 
	.CO(n1921), 
	.CI(n1935), 
	.B(n1930), 
	.A(n1926));
   FA_X1 U1362 (.S(n1924), 
	.CO(n1923), 
	.CI(n1928), 
	.B(n1939), 
	.A(n1937));
   FA_X1 U1363 (.S(n1926), 
	.CO(n1925), 
	.CI(n1941), 
	.B(n2456), 
	.A(n2426));
   FA_X1 U1364 (.S(n1928), 
	.CO(n1927), 
	.CI(n2396), 
	.B(n2486), 
	.A(n2366));
   FA_X1 U1365 (.S(n1930), 
	.CO(n1929), 
	.CI(n2306), 
	.B(n2517), 
	.A(n2336));
   FA_X1 U1366 (.S(n1932), 
	.CO(n1931), 
	.CI(n1934), 
	.B(n1936), 
	.A(n1945));
   FA_X1 U1367 (.S(n1934), 
	.CO(n1933), 
	.CI(n1947), 
	.B(n1938), 
	.A(n1940));
   FA_X1 U1368 (.S(n1936), 
	.CO(n1935), 
	.CI(n1949), 
	.B(n1942), 
	.A(n1951));
   FA_X1 U1369 (.S(n1938), 
	.CO(n1937), 
	.CI(n2397), 
	.B(n2457), 
	.A(n2367));
   FA_X1 U1370 (.S(n1940), 
	.CO(n1939), 
	.CI(n2487), 
	.B(n2427), 
	.A(n2518));
   HA_X1 U1371 (.S(n1942), 
	.CO(n1941), 
	.B(n2012), 
	.A(n2337));
   FA_X1 U1372 (.S(n1944), 
	.CO(n1943), 
	.CI(n1946), 
	.B(n1955), 
	.A(n1948));
   FA_X1 U1373 (.S(n1946), 
	.CO(n1945), 
	.CI(n1957), 
	.B(n1950), 
	.A(n1952));
   FA_X1 U1374 (.S(n1948), 
	.CO(n1947), 
	.CI(n1959), 
	.B(n2458), 
	.A(n1961));
   FA_X1 U1375 (.S(n1950), 
	.CO(n1949), 
	.CI(n2428), 
	.B(n2488), 
	.A(n2398));
   FA_X1 U1376 (.S(n1952), 
	.CO(n1951), 
	.CI(n2338), 
	.B(n2519), 
	.A(n2368));
   FA_X1 U1377 (.S(n1954), 
	.CO(n1953), 
	.CI(n1956), 
	.B(n1958), 
	.A(n1965));
   FA_X1 U1378 (.S(n1956), 
	.CO(n1955), 
	.CI(n1960), 
	.B(n1969), 
	.A(n1967));
   FA_X1 U1379 (.S(n1958), 
	.CO(n1957), 
	.CI(n1962), 
	.B(n2429), 
	.A(n2399));
   FA_X1 U1380 (.S(n1960), 
	.CO(n1959), 
	.CI(n2489), 
	.B(n2459), 
	.A(n2520));
   HA_X1 U1381 (.S(n1962), 
	.CO(n1961), 
	.B(n2013), 
	.A(n2369));
   FA_X1 U1382 (.S(n1964), 
	.CO(n1963), 
	.CI(n1966), 
	.B(n1970), 
	.A(n1973));
   FA_X1 U1383 (.S(n1966), 
	.CO(n1965), 
	.CI(n1968), 
	.B(n1977), 
	.A(n1975));
   FA_X1 U1384 (.S(n1968), 
	.CO(n1967), 
	.CI(n2460), 
	.B(n2490), 
	.A(n2430));
   FA_X1 U1385 (.S(n1970), 
	.CO(n1969), 
	.CI(n2370), 
	.B(n2521), 
	.A(n2400));
   FA_X1 U1386 (.S(n1972), 
	.CO(n1971), 
	.CI(n1974), 
	.B(n1981), 
	.A(n1976));
   FA_X1 U1387 (.S(n1974), 
	.CO(n1973), 
	.CI(n1983), 
	.B(n2522), 
	.A(n1978));
   FA_X1 U1388 (.S(n1976), 
	.CO(n1975), 
	.CI(n2491), 
	.B(n2461), 
	.A(n2431));
   HA_X1 U1389 (.S(n1978), 
	.CO(n1977), 
	.B(n2014), 
	.A(n2401));
   FA_X1 U1390 (.S(n1980), 
	.CO(n1979), 
	.CI(n1982), 
	.B(n1987), 
	.A(n1984));
   FA_X1 U1391 (.S(n1982), 
	.CO(n1981), 
	.CI(n1989), 
	.B(n2492), 
	.A(n2462));
   FA_X1 U1392 (.S(n1984), 
	.CO(n1983), 
	.CI(n2402), 
	.B(n2523), 
	.A(n2432));
   FA_X1 U1393 (.S(n1986), 
	.CO(n1985), 
	.CI(n1988), 
	.B(n1990), 
	.A(n1993));
   FA_X1 U1394 (.S(n1988), 
	.CO(n1987), 
	.CI(n2493), 
	.B(n2524), 
	.A(n2463));
   HA_X1 U1395 (.S(n1990), 
	.CO(n1989), 
	.B(n2015), 
	.A(n2433));
   FA_X1 U1396 (.S(n1992), 
	.CO(n1991), 
	.CI(n1994), 
	.B(n2494), 
	.A(n1997));
   FA_X1 U1397 (.S(n1994), 
	.CO(n1993), 
	.CI(n2434), 
	.B(n2525), 
	.A(n2464));
   FA_X1 U1398 (.S(n1996), 
	.CO(n1995), 
	.CI(n1998), 
	.B(n2526), 
	.A(n2495));
   HA_X1 U1399 (.S(n1998), 
	.CO(n1997), 
	.B(n2016), 
	.A(n2465));
   FA_X1 U1400 (.S(n2000), 
	.CO(n1999), 
	.CI(n2466), 
	.B(n2527), 
	.A(n2496));
   HA_X1 U1401 (.S(n2002), 
	.CO(n2001), 
	.B(n2497), 
	.A(n2528));
   OAI22_X1 U1402 (.ZN(n2003), 
	.B2(FE_OFN35_n3123), 
	.B1(n2563), 
	.A2(FE_PT1_n949), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1404 (.ZN(n2020), 
	.B2(FE_OFN35_n3123), 
	.B1(n2532), 
	.A2(n2533), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1405 (.ZN(n2021), 
	.B2(FE_OFN35_n3123), 
	.B1(n2533), 
	.A2(n2534), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1406 (.ZN(n2022), 
	.B2(FE_OFN35_n3123), 
	.B1(n2534), 
	.A2(n2535), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1407 (.ZN(n2023), 
	.B2(FE_OFN35_n3123), 
	.B1(n2535), 
	.A2(n2536), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1408 (.ZN(n2024), 
	.B2(FE_OFN35_n3123), 
	.B1(n2536), 
	.A2(n2537), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1409 (.ZN(n2025), 
	.B2(FE_OFN35_n3123), 
	.B1(n2537), 
	.A2(n2538), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1410 (.ZN(n2026), 
	.B2(FE_OFN35_n3123), 
	.B1(n2538), 
	.A2(n2539), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1411 (.ZN(n2027), 
	.B2(FE_OFN35_n3123), 
	.B1(n2539), 
	.A2(n2540), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1412 (.ZN(n2028), 
	.B2(FE_OFN35_n3123), 
	.B1(n2540), 
	.A2(n2541), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1413 (.ZN(n2029), 
	.B2(FE_OFN35_n3123), 
	.B1(n2541), 
	.A2(n2542), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1414 (.ZN(n2030), 
	.B2(FE_OFN35_n3123), 
	.B1(n2542), 
	.A2(n2543), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1415 (.ZN(n2031), 
	.B2(FE_OFN35_n3123), 
	.B1(n2543), 
	.A2(n2544), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1416 (.ZN(n2032), 
	.B2(FE_OFN35_n3123), 
	.B1(n2544), 
	.A2(n2545), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1417 (.ZN(n2033), 
	.B2(FE_OFN35_n3123), 
	.B1(n2545), 
	.A2(n2546), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1418 (.ZN(n2034), 
	.B2(FE_OFN35_n3123), 
	.B1(n2546), 
	.A2(n2547), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1419 (.ZN(n2035), 
	.B2(FE_OFN35_n3123), 
	.B1(n2547), 
	.A2(n2548), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1420 (.ZN(n2036), 
	.B2(FE_OFN35_n3123), 
	.B1(n2548), 
	.A2(n2549), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1421 (.ZN(n2037), 
	.B2(FE_OFN35_n3123), 
	.B1(n2549), 
	.A2(n2550), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1422 (.ZN(n2038), 
	.B2(FE_OFN35_n3123), 
	.B1(n2550), 
	.A2(n2551), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1423 (.ZN(n2039), 
	.B2(FE_OFN35_n3123), 
	.B1(n2551), 
	.A2(n2552), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1424 (.ZN(n2040), 
	.B2(FE_OFN35_n3123), 
	.B1(n2552), 
	.A2(n2553), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1425 (.ZN(n2041), 
	.B2(FE_OFN35_n3123), 
	.B1(n2553), 
	.A2(n2554), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1426 (.ZN(n2042), 
	.B2(FE_OFN35_n3123), 
	.B1(n2554), 
	.A2(n2555), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1427 (.ZN(n2043), 
	.B2(FE_OFN35_n3123), 
	.B1(n2555), 
	.A2(n2556), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1428 (.ZN(n2044), 
	.B2(FE_OFN35_n3123), 
	.B1(n2556), 
	.A2(n2557), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1429 (.ZN(n2045), 
	.B2(FE_OFN35_n3123), 
	.B1(n2557), 
	.A2(n2558), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1430 (.ZN(n2046), 
	.B2(FE_OFN35_n3123), 
	.B1(n2558), 
	.A2(n2559), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1431 (.ZN(n2047), 
	.B2(FE_OFN35_n3123), 
	.B1(n2559), 
	.A2(n2560), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1432 (.ZN(n2048), 
	.B2(FE_OFN35_n3123), 
	.B1(n2560), 
	.A2(n2561), 
	.A1(FE_OFN34_n3107));
   OAI22_X1 U1433 (.ZN(n2049), 
	.B2(FE_OFN35_n3123), 
	.B1(n2561), 
	.A2(n2562), 
	.A1(FE_OFN34_n3107));
   XNOR2_X1 U1434 (.ZN(n2531), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[31]));
   XNOR2_X1 U1435 (.ZN(n2532), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[30]));
   XNOR2_X1 U1436 (.ZN(n2533), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[29]));
   XNOR2_X1 U1437 (.ZN(n2534), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1438 (.ZN(n2535), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1439 (.ZN(n2536), 
	.B(a[31]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1440 (.ZN(n2537), 
	.B(a[31]), 
	.A(b[25]));
   XNOR2_X1 U1441 (.ZN(n2538), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1442 (.ZN(n2539), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1443 (.ZN(n2540), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1444 (.ZN(n2541), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1445 (.ZN(n2542), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1446 (.ZN(n2543), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[19]));
   XNOR2_X1 U1447 (.ZN(n2544), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1448 (.ZN(n2545), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[17]));
   XNOR2_X1 U1449 (.ZN(n2546), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[16]));
   XNOR2_X1 U1450 (.ZN(n2547), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[15]));
   XNOR2_X1 U1451 (.ZN(n2548), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[14]));
   XNOR2_X1 U1452 (.ZN(n2549), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1453 (.ZN(n2550), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1454 (.ZN(n2551), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1455 (.ZN(n2552), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1456 (.ZN(n2553), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(b[9]));
   XNOR2_X1 U1457 (.ZN(n2554), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1458 (.ZN(n2555), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1459 (.ZN(n2556), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1460 (.ZN(n2557), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1461 (.ZN(n2558), 
	.B(FE_OFN178_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1462 (.ZN(n2559), 
	.B(a[31]), 
	.A(b[3]));
   XNOR2_X1 U1463 (.ZN(n2560), 
	.B(a[31]), 
	.A(b[2]));
   XNOR2_X1 U1464 (.ZN(n2561), 
	.B(a[31]), 
	.A(b[1]));
   XNOR2_X1 U1465 (.ZN(n2562), 
	.B(a[31]), 
	.A(b[0]));
   OAI22_X1 U1466 (.ZN(n2004), 
	.B2(FE_OFN36_n3124), 
	.B1(n2596), 
	.A2(n3140), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1468 (.ZN(n2052), 
	.B2(FE_OFN36_n3124), 
	.B1(n2565), 
	.A2(n2566), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1469 (.ZN(n2053), 
	.B2(FE_OFN36_n3124), 
	.B1(n2566), 
	.A2(n2567), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1470 (.ZN(n2054), 
	.B2(FE_OFN36_n3124), 
	.B1(n2567), 
	.A2(n2568), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1471 (.ZN(n2055), 
	.B2(FE_OFN36_n3124), 
	.B1(n2568), 
	.A2(n2569), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1472 (.ZN(n2056), 
	.B2(FE_OFN36_n3124), 
	.B1(n2569), 
	.A2(n2570), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1473 (.ZN(n2057), 
	.B2(FE_OFN36_n3124), 
	.B1(n2570), 
	.A2(n2571), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1474 (.ZN(n2058), 
	.B2(FE_OFN36_n3124), 
	.B1(n2571), 
	.A2(n2572), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1475 (.ZN(n2059), 
	.B2(FE_OFN36_n3124), 
	.B1(n2572), 
	.A2(n2573), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1476 (.ZN(n2060), 
	.B2(FE_OFN36_n3124), 
	.B1(n2573), 
	.A2(n2574), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1477 (.ZN(n2061), 
	.B2(FE_OFN36_n3124), 
	.B1(n2574), 
	.A2(n2575), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1478 (.ZN(n2062), 
	.B2(FE_OFN36_n3124), 
	.B1(n2575), 
	.A2(n2576), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1479 (.ZN(n2063), 
	.B2(FE_OFN36_n3124), 
	.B1(n2576), 
	.A2(n2577), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1480 (.ZN(n2064), 
	.B2(FE_OFN36_n3124), 
	.B1(n2577), 
	.A2(n2578), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1481 (.ZN(n2065), 
	.B2(FE_OFN36_n3124), 
	.B1(n2578), 
	.A2(n2579), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1482 (.ZN(n2066), 
	.B2(FE_OFN36_n3124), 
	.B1(n2579), 
	.A2(n2580), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1483 (.ZN(n2067), 
	.B2(FE_OFN36_n3124), 
	.B1(n2580), 
	.A2(n2581), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1484 (.ZN(n2068), 
	.B2(FE_OFN36_n3124), 
	.B1(n2581), 
	.A2(n2582), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1485 (.ZN(n2069), 
	.B2(FE_OFN36_n3124), 
	.B1(n2582), 
	.A2(n2583), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1486 (.ZN(n2070), 
	.B2(FE_OFN36_n3124), 
	.B1(n2583), 
	.A2(n2584), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1487 (.ZN(n2071), 
	.B2(FE_OFN36_n3124), 
	.B1(n2584), 
	.A2(n2585), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1488 (.ZN(n2072), 
	.B2(FE_OFN36_n3124), 
	.B1(n2585), 
	.A2(n2586), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1489 (.ZN(n2073), 
	.B2(FE_OFN36_n3124), 
	.B1(n2586), 
	.A2(n2587), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1490 (.ZN(n2074), 
	.B2(FE_OFN36_n3124), 
	.B1(n2587), 
	.A2(n2588), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1491 (.ZN(n2075), 
	.B2(FE_OFN36_n3124), 
	.B1(n2588), 
	.A2(n2589), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1492 (.ZN(n2076), 
	.B2(FE_OFN36_n3124), 
	.B1(n2589), 
	.A2(n2590), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1493 (.ZN(n2077), 
	.B2(FE_OFN36_n3124), 
	.B1(n2590), 
	.A2(n2591), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1494 (.ZN(n2078), 
	.B2(FE_OFN36_n3124), 
	.B1(n2591), 
	.A2(n2592), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1495 (.ZN(n2079), 
	.B2(FE_OFN36_n3124), 
	.B1(n2592), 
	.A2(n2593), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1496 (.ZN(n2080), 
	.B2(FE_OFN36_n3124), 
	.B1(n2593), 
	.A2(n2594), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U1497 (.ZN(n2081), 
	.B2(FE_OFN36_n3124), 
	.B1(n2594), 
	.A2(n2595), 
	.A1(FE_OFN33_n3108));
   XNOR2_X1 U1498 (.ZN(n2564), 
	.B(a[29]), 
	.A(b[31]));
   XNOR2_X1 U1499 (.ZN(n2565), 
	.B(a[29]), 
	.A(b[30]));
   XNOR2_X1 U1500 (.ZN(n2566), 
	.B(a[29]), 
	.A(b[29]));
   XNOR2_X1 U1501 (.ZN(n2567), 
	.B(a[29]), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1502 (.ZN(n2568), 
	.B(a[29]), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1503 (.ZN(n2569), 
	.B(a[29]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1504 (.ZN(n2570), 
	.B(a[29]), 
	.A(b[25]));
   XNOR2_X1 U1505 (.ZN(n2571), 
	.B(a[29]), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1506 (.ZN(n2572), 
	.B(a[29]), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1507 (.ZN(n2573), 
	.B(a[29]), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1508 (.ZN(n2574), 
	.B(a[29]), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1509 (.ZN(n2575), 
	.B(a[29]), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1510 (.ZN(n2576), 
	.B(a[29]), 
	.A(b[19]));
   XNOR2_X1 U1511 (.ZN(n2577), 
	.B(a[29]), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1512 (.ZN(n2578), 
	.B(a[29]), 
	.A(b[17]));
   XNOR2_X1 U1513 (.ZN(n2579), 
	.B(a[29]), 
	.A(b[16]));
   XNOR2_X1 U1514 (.ZN(n2580), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(b[15]));
   XNOR2_X1 U1515 (.ZN(n2581), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(b[14]));
   XNOR2_X1 U1516 (.ZN(n2582), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1517 (.ZN(n2583), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1518 (.ZN(n2584), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1519 (.ZN(n2585), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1520 (.ZN(n2586), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(b[9]));
   XNOR2_X1 U1521 (.ZN(n2587), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1522 (.ZN(n2588), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1523 (.ZN(n2589), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1524 (.ZN(n2590), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1525 (.ZN(n2591), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1526 (.ZN(n2592), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1527 (.ZN(n2593), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(b[2]));
   XNOR2_X1 U1528 (.ZN(n2594), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(b[1]));
   XNOR2_X1 U1529 (.ZN(n2595), 
	.B(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1530 (.ZN(n2005), 
	.B2(FE_OFN38_n3125), 
	.B1(n2629), 
	.A2(n3141), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1532 (.ZN(n2084), 
	.B2(FE_OFN38_n3125), 
	.B1(n2598), 
	.A2(n2599), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1533 (.ZN(n2085), 
	.B2(FE_OFN38_n3125), 
	.B1(n2599), 
	.A2(n2600), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1534 (.ZN(n2086), 
	.B2(FE_OFN38_n3125), 
	.B1(n2600), 
	.A2(n2601), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1535 (.ZN(n2087), 
	.B2(FE_OFN38_n3125), 
	.B1(n2601), 
	.A2(n2602), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1536 (.ZN(n2088), 
	.B2(FE_OFN38_n3125), 
	.B1(n2602), 
	.A2(n2603), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1537 (.ZN(n2089), 
	.B2(FE_OFN38_n3125), 
	.B1(n2603), 
	.A2(n2604), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1538 (.ZN(n2090), 
	.B2(FE_OFN38_n3125), 
	.B1(n2604), 
	.A2(n2605), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1539 (.ZN(n2091), 
	.B2(FE_OFN38_n3125), 
	.B1(n2605), 
	.A2(n2606), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1540 (.ZN(n2092), 
	.B2(FE_OFN38_n3125), 
	.B1(n2606), 
	.A2(n2607), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1541 (.ZN(n2093), 
	.B2(FE_OFN38_n3125), 
	.B1(n2607), 
	.A2(n2608), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1542 (.ZN(n2094), 
	.B2(FE_OFN38_n3125), 
	.B1(n2608), 
	.A2(n2609), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1543 (.ZN(n2095), 
	.B2(FE_OFN38_n3125), 
	.B1(n2609), 
	.A2(n2610), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1544 (.ZN(n2096), 
	.B2(FE_OFN38_n3125), 
	.B1(n2610), 
	.A2(n2611), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1545 (.ZN(n2097), 
	.B2(FE_OFN38_n3125), 
	.B1(n2611), 
	.A2(n2612), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1546 (.ZN(n2098), 
	.B2(FE_OFN38_n3125), 
	.B1(n2612), 
	.A2(n2613), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1547 (.ZN(n2099), 
	.B2(FE_OFN38_n3125), 
	.B1(n2613), 
	.A2(n2614), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1548 (.ZN(n2100), 
	.B2(FE_OFN38_n3125), 
	.B1(n2614), 
	.A2(n2615), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1549 (.ZN(n2101), 
	.B2(FE_OFN38_n3125), 
	.B1(n2615), 
	.A2(n2616), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1550 (.ZN(n2102), 
	.B2(FE_OFN38_n3125), 
	.B1(n2616), 
	.A2(n2617), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1551 (.ZN(n2103), 
	.B2(FE_OFN38_n3125), 
	.B1(n2617), 
	.A2(n2618), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1552 (.ZN(n2104), 
	.B2(FE_OFN38_n3125), 
	.B1(n2618), 
	.A2(n2619), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1553 (.ZN(n2105), 
	.B2(FE_OFN38_n3125), 
	.B1(n2619), 
	.A2(n2620), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1554 (.ZN(n2106), 
	.B2(FE_OFN38_n3125), 
	.B1(n2620), 
	.A2(n2621), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1555 (.ZN(n2107), 
	.B2(FE_OFN38_n3125), 
	.B1(n2621), 
	.A2(n2622), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1556 (.ZN(n2108), 
	.B2(FE_OFN38_n3125), 
	.B1(n2622), 
	.A2(n2623), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1557 (.ZN(n2109), 
	.B2(FE_OFN38_n3125), 
	.B1(n2623), 
	.A2(n2624), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1558 (.ZN(n2110), 
	.B2(FE_OFN38_n3125), 
	.B1(n2624), 
	.A2(n2625), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1559 (.ZN(n2111), 
	.B2(FE_OFN38_n3125), 
	.B1(n2625), 
	.A2(n2626), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1560 (.ZN(n2112), 
	.B2(FE_OFN38_n3125), 
	.B1(n2626), 
	.A2(n2627), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U1561 (.ZN(n2113), 
	.B2(FE_OFN38_n3125), 
	.B1(n2627), 
	.A2(n2628), 
	.A1(FE_OFN37_n3109));
   XNOR2_X1 U1562 (.ZN(n2597), 
	.B(a[27]), 
	.A(b[31]));
   XNOR2_X1 U1563 (.ZN(n2598), 
	.B(a[27]), 
	.A(b[30]));
   XNOR2_X1 U1564 (.ZN(n2599), 
	.B(a[27]), 
	.A(b[29]));
   XNOR2_X1 U1565 (.ZN(n2600), 
	.B(a[27]), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1566 (.ZN(n2601), 
	.B(a[27]), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1567 (.ZN(n2602), 
	.B(a[27]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1568 (.ZN(n2603), 
	.B(a[27]), 
	.A(b[25]));
   XNOR2_X1 U1569 (.ZN(n2604), 
	.B(a[27]), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1570 (.ZN(n2605), 
	.B(a[27]), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1571 (.ZN(n2606), 
	.B(a[27]), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1572 (.ZN(n2607), 
	.B(a[27]), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1573 (.ZN(n2608), 
	.B(a[27]), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1574 (.ZN(n2609), 
	.B(a[27]), 
	.A(b[19]));
   XNOR2_X1 U1575 (.ZN(n2610), 
	.B(a[27]), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1576 (.ZN(n2611), 
	.B(a[27]), 
	.A(b[17]));
   XNOR2_X1 U1577 (.ZN(n2612), 
	.B(a[27]), 
	.A(b[16]));
   XNOR2_X1 U1578 (.ZN(n2613), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(b[15]));
   XNOR2_X1 U1579 (.ZN(n2614), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(b[14]));
   XNOR2_X1 U1580 (.ZN(n2615), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1581 (.ZN(n2616), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1582 (.ZN(n2617), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1583 (.ZN(n2618), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1584 (.ZN(n2619), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(b[9]));
   XNOR2_X1 U1585 (.ZN(n2620), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1586 (.ZN(n2621), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1587 (.ZN(n2622), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1588 (.ZN(n2623), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1589 (.ZN(n2624), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1590 (.ZN(n2625), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1591 (.ZN(n2626), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(b[2]));
   XNOR2_X1 U1592 (.ZN(n2627), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(b[1]));
   XNOR2_X1 U1593 (.ZN(n2628), 
	.B(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1594 (.ZN(n2006), 
	.B2(FE_OFN40_n3126), 
	.B1(n2662), 
	.A2(n3142), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1596 (.ZN(n2116), 
	.B2(FE_OFN40_n3126), 
	.B1(n2631), 
	.A2(n2632), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1597 (.ZN(n2117), 
	.B2(FE_OFN40_n3126), 
	.B1(n2632), 
	.A2(n2633), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1598 (.ZN(n2118), 
	.B2(FE_OFN40_n3126), 
	.B1(n2633), 
	.A2(n2634), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1599 (.ZN(n2119), 
	.B2(FE_OFN40_n3126), 
	.B1(n2634), 
	.A2(n2635), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1600 (.ZN(n2120), 
	.B2(FE_OFN40_n3126), 
	.B1(n2635), 
	.A2(n2636), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1601 (.ZN(n2121), 
	.B2(FE_OFN40_n3126), 
	.B1(n2636), 
	.A2(n2637), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1602 (.ZN(n2122), 
	.B2(FE_OFN40_n3126), 
	.B1(n2637), 
	.A2(n2638), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1603 (.ZN(n2123), 
	.B2(FE_OFN40_n3126), 
	.B1(n2638), 
	.A2(n2639), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1604 (.ZN(n2124), 
	.B2(FE_OFN40_n3126), 
	.B1(n2639), 
	.A2(n2640), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1605 (.ZN(n2125), 
	.B2(FE_OFN40_n3126), 
	.B1(n2640), 
	.A2(n2641), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1606 (.ZN(n2126), 
	.B2(FE_OFN40_n3126), 
	.B1(n2641), 
	.A2(n2642), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1607 (.ZN(n2127), 
	.B2(FE_OFN40_n3126), 
	.B1(n2642), 
	.A2(n2643), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1608 (.ZN(n2128), 
	.B2(FE_OFN40_n3126), 
	.B1(n2643), 
	.A2(n2644), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1609 (.ZN(n2129), 
	.B2(FE_OFN40_n3126), 
	.B1(n2644), 
	.A2(n2645), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1610 (.ZN(n2130), 
	.B2(FE_OFN40_n3126), 
	.B1(n2645), 
	.A2(n2646), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1611 (.ZN(n2131), 
	.B2(FE_OFN40_n3126), 
	.B1(n2646), 
	.A2(n2647), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1612 (.ZN(n2132), 
	.B2(FE_OFN40_n3126), 
	.B1(n2647), 
	.A2(n2648), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1613 (.ZN(n2133), 
	.B2(FE_OFN40_n3126), 
	.B1(n2648), 
	.A2(n2649), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1614 (.ZN(n2134), 
	.B2(FE_OFN40_n3126), 
	.B1(n2649), 
	.A2(n2650), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1615 (.ZN(n2135), 
	.B2(FE_OFN40_n3126), 
	.B1(n2650), 
	.A2(n2651), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1616 (.ZN(n2136), 
	.B2(FE_OFN40_n3126), 
	.B1(n2651), 
	.A2(n2652), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1617 (.ZN(n2137), 
	.B2(FE_OFN40_n3126), 
	.B1(n2652), 
	.A2(n2653), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1618 (.ZN(n2138), 
	.B2(FE_OFN40_n3126), 
	.B1(n2653), 
	.A2(n2654), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1619 (.ZN(n2139), 
	.B2(FE_OFN40_n3126), 
	.B1(n2654), 
	.A2(n2655), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1620 (.ZN(n2140), 
	.B2(FE_OFN40_n3126), 
	.B1(n2655), 
	.A2(n2656), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1621 (.ZN(n2141), 
	.B2(FE_OFN40_n3126), 
	.B1(n2656), 
	.A2(n2657), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1622 (.ZN(n2142), 
	.B2(FE_OFN40_n3126), 
	.B1(n2657), 
	.A2(n2658), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1623 (.ZN(n2143), 
	.B2(FE_OFN40_n3126), 
	.B1(n2658), 
	.A2(n2659), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1624 (.ZN(n2144), 
	.B2(FE_OFN40_n3126), 
	.B1(n2659), 
	.A2(n2660), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U1625 (.ZN(n2145), 
	.B2(FE_OFN40_n3126), 
	.B1(n2660), 
	.A2(n2661), 
	.A1(FE_OFN39_n3110));
   XNOR2_X1 U1626 (.ZN(n2630), 
	.B(a[25]), 
	.A(b[31]));
   XNOR2_X1 U1627 (.ZN(n2631), 
	.B(a[25]), 
	.A(b[30]));
   XNOR2_X1 U1628 (.ZN(n2632), 
	.B(a[25]), 
	.A(b[29]));
   XNOR2_X1 U1629 (.ZN(n2633), 
	.B(a[25]), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1630 (.ZN(n2634), 
	.B(a[25]), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1631 (.ZN(n2635), 
	.B(a[25]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1632 (.ZN(n2636), 
	.B(a[25]), 
	.A(b[25]));
   XNOR2_X1 U1633 (.ZN(n2637), 
	.B(a[25]), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1634 (.ZN(n2638), 
	.B(a[25]), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1635 (.ZN(n2639), 
	.B(a[25]), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1636 (.ZN(n2640), 
	.B(a[25]), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1637 (.ZN(n2641), 
	.B(a[25]), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1638 (.ZN(n2642), 
	.B(a[25]), 
	.A(b[19]));
   XNOR2_X1 U1639 (.ZN(n2643), 
	.B(a[25]), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1640 (.ZN(n2644), 
	.B(a[25]), 
	.A(b[17]));
   XNOR2_X1 U1641 (.ZN(n2645), 
	.B(a[25]), 
	.A(b[16]));
   XNOR2_X1 U1642 (.ZN(n2646), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(b[15]));
   XNOR2_X1 U1643 (.ZN(n2647), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(b[14]));
   XNOR2_X1 U1644 (.ZN(n2648), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1645 (.ZN(n2649), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1646 (.ZN(n2650), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1647 (.ZN(n2651), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1648 (.ZN(n2652), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(b[9]));
   XNOR2_X1 U1649 (.ZN(n2653), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1650 (.ZN(n2654), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1651 (.ZN(n2655), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1652 (.ZN(n2656), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1653 (.ZN(n2657), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1654 (.ZN(n2658), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1655 (.ZN(n2659), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(b[2]));
   XNOR2_X1 U1656 (.ZN(n2660), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(b[1]));
   XNOR2_X1 U1657 (.ZN(n2661), 
	.B(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1658 (.ZN(n2007), 
	.B2(FE_OFN42_n3127), 
	.B1(n2695), 
	.A2(FE_PT1_n808), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1660 (.ZN(n2148), 
	.B2(FE_OFN42_n3127), 
	.B1(n2664), 
	.A2(n2665), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1661 (.ZN(n2149), 
	.B2(FE_OFN42_n3127), 
	.B1(n2665), 
	.A2(n2666), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1662 (.ZN(n2150), 
	.B2(FE_OFN42_n3127), 
	.B1(n2666), 
	.A2(n2667), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1663 (.ZN(n2151), 
	.B2(FE_OFN42_n3127), 
	.B1(n2667), 
	.A2(n2668), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1664 (.ZN(n2152), 
	.B2(FE_OFN42_n3127), 
	.B1(n2668), 
	.A2(n2669), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1665 (.ZN(n2153), 
	.B2(FE_OFN42_n3127), 
	.B1(n2669), 
	.A2(n2670), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1666 (.ZN(n2154), 
	.B2(FE_OFN42_n3127), 
	.B1(n2670), 
	.A2(n2671), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1667 (.ZN(n2155), 
	.B2(FE_OFN42_n3127), 
	.B1(n2671), 
	.A2(n2672), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1668 (.ZN(n2156), 
	.B2(FE_OFN42_n3127), 
	.B1(n2672), 
	.A2(n2673), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1669 (.ZN(n2157), 
	.B2(FE_OFN42_n3127), 
	.B1(n2673), 
	.A2(n2674), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1670 (.ZN(n2158), 
	.B2(FE_OFN42_n3127), 
	.B1(n2674), 
	.A2(n2675), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1671 (.ZN(n2159), 
	.B2(FE_OFN42_n3127), 
	.B1(n2675), 
	.A2(n2676), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1672 (.ZN(n2160), 
	.B2(FE_OFN42_n3127), 
	.B1(n2676), 
	.A2(n2677), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1673 (.ZN(n2161), 
	.B2(FE_OFN42_n3127), 
	.B1(n2677), 
	.A2(n2678), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1674 (.ZN(n2162), 
	.B2(FE_OFN42_n3127), 
	.B1(n2678), 
	.A2(n2679), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1675 (.ZN(n2163), 
	.B2(FE_OFN42_n3127), 
	.B1(n2679), 
	.A2(n2680), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1676 (.ZN(n2164), 
	.B2(FE_OFN42_n3127), 
	.B1(n2680), 
	.A2(n2681), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1677 (.ZN(n2165), 
	.B2(FE_OFN42_n3127), 
	.B1(n2681), 
	.A2(n2682), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1678 (.ZN(n2166), 
	.B2(FE_OFN42_n3127), 
	.B1(n2682), 
	.A2(n2683), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1679 (.ZN(n2167), 
	.B2(FE_OFN42_n3127), 
	.B1(n2683), 
	.A2(n2684), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1680 (.ZN(n2168), 
	.B2(FE_OFN42_n3127), 
	.B1(n2684), 
	.A2(n2685), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1681 (.ZN(n2169), 
	.B2(FE_OFN42_n3127), 
	.B1(n2685), 
	.A2(n2686), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1682 (.ZN(n2170), 
	.B2(FE_OFN42_n3127), 
	.B1(n2686), 
	.A2(n2687), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1683 (.ZN(n2171), 
	.B2(FE_OFN42_n3127), 
	.B1(n2687), 
	.A2(n2688), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1684 (.ZN(n2172), 
	.B2(FE_OFN42_n3127), 
	.B1(n2688), 
	.A2(n2689), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1685 (.ZN(n2173), 
	.B2(FE_OFN42_n3127), 
	.B1(n2689), 
	.A2(n2690), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1686 (.ZN(n2174), 
	.B2(FE_OFN42_n3127), 
	.B1(n2690), 
	.A2(n2691), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1687 (.ZN(n2175), 
	.B2(FE_OFN42_n3127), 
	.B1(n2691), 
	.A2(n2692), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1688 (.ZN(n2176), 
	.B2(FE_OFN42_n3127), 
	.B1(n2692), 
	.A2(n2693), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U1689 (.ZN(n2177), 
	.B2(FE_OFN42_n3127), 
	.B1(n2693), 
	.A2(n2694), 
	.A1(FE_OFN41_n3111));
   XNOR2_X1 U1690 (.ZN(n2663), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U1691 (.ZN(n2664), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U1692 (.ZN(n2665), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[29]));
   XNOR2_X1 U1693 (.ZN(n2666), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1694 (.ZN(n2667), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1695 (.ZN(n2668), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1696 (.ZN(n2669), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[25]));
   XNOR2_X1 U1697 (.ZN(n2670), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1698 (.ZN(n2671), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1699 (.ZN(n2672), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1700 (.ZN(n2673), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1701 (.ZN(n2674), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1702 (.ZN(n2675), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[19]));
   XNOR2_X1 U1703 (.ZN(n2676), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1704 (.ZN(n2677), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[17]));
   XNOR2_X1 U1705 (.ZN(n2678), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[16]));
   XNOR2_X1 U1706 (.ZN(n2679), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[15]));
   XNOR2_X1 U1707 (.ZN(n2680), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[14]));
   XNOR2_X1 U1708 (.ZN(n2681), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1709 (.ZN(n2682), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1710 (.ZN(n2683), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1711 (.ZN(n2684), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1712 (.ZN(n2685), 
	.B(FE_OFN174_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(b[9]));
   XNOR2_X1 U1713 (.ZN(n2686), 
	.B(a[23]), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1714 (.ZN(n2687), 
	.B(a[23]), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1715 (.ZN(n2688), 
	.B(a[23]), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1716 (.ZN(n2689), 
	.B(a[23]), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1717 (.ZN(n2690), 
	.B(a[23]), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1718 (.ZN(n2691), 
	.B(a[23]), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1719 (.ZN(n2692), 
	.B(a[23]), 
	.A(b[2]));
   XNOR2_X1 U1720 (.ZN(n2693), 
	.B(a[23]), 
	.A(b[1]));
   XNOR2_X1 U1721 (.ZN(n2694), 
	.B(a[23]), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1722 (.ZN(n2008), 
	.B2(FE_OFN44_n3128), 
	.B1(n2728), 
	.A2(n338), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1724 (.ZN(n2180), 
	.B2(FE_OFN44_n3128), 
	.B1(n2697), 
	.A2(n2698), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1725 (.ZN(n2181), 
	.B2(FE_OFN44_n3128), 
	.B1(n2698), 
	.A2(n2699), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1726 (.ZN(n2182), 
	.B2(FE_OFN44_n3128), 
	.B1(n2699), 
	.A2(n2700), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1727 (.ZN(n2183), 
	.B2(FE_OFN44_n3128), 
	.B1(n2700), 
	.A2(n2701), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1728 (.ZN(n2184), 
	.B2(FE_OFN44_n3128), 
	.B1(n2701), 
	.A2(n2702), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1729 (.ZN(n2185), 
	.B2(FE_OFN44_n3128), 
	.B1(n2702), 
	.A2(n2703), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1730 (.ZN(n2186), 
	.B2(FE_OFN44_n3128), 
	.B1(n2703), 
	.A2(n2704), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1731 (.ZN(n2187), 
	.B2(FE_OFN44_n3128), 
	.B1(n2704), 
	.A2(n2705), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1732 (.ZN(n2188), 
	.B2(FE_OFN44_n3128), 
	.B1(n2705), 
	.A2(n2706), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1733 (.ZN(n2189), 
	.B2(FE_OFN44_n3128), 
	.B1(n2706), 
	.A2(n2707), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1734 (.ZN(n2190), 
	.B2(FE_OFN44_n3128), 
	.B1(n2707), 
	.A2(n2708), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1735 (.ZN(n2191), 
	.B2(FE_OFN44_n3128), 
	.B1(n2708), 
	.A2(n2709), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1736 (.ZN(n2192), 
	.B2(FE_OFN44_n3128), 
	.B1(n2709), 
	.A2(n2710), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1737 (.ZN(n2193), 
	.B2(FE_OFN44_n3128), 
	.B1(n2710), 
	.A2(n2711), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1738 (.ZN(n2194), 
	.B2(FE_OFN44_n3128), 
	.B1(n2711), 
	.A2(n2712), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1739 (.ZN(n2195), 
	.B2(FE_OFN44_n3128), 
	.B1(n2712), 
	.A2(n2713), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1740 (.ZN(n2196), 
	.B2(FE_OFN44_n3128), 
	.B1(n2713), 
	.A2(n2714), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1741 (.ZN(n2197), 
	.B2(FE_OFN44_n3128), 
	.B1(n2714), 
	.A2(n2715), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1742 (.ZN(n2198), 
	.B2(FE_OFN44_n3128), 
	.B1(n2715), 
	.A2(n2716), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1743 (.ZN(n2199), 
	.B2(FE_OFN44_n3128), 
	.B1(n2716), 
	.A2(n2717), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1744 (.ZN(n2200), 
	.B2(FE_OFN44_n3128), 
	.B1(n2717), 
	.A2(n2718), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1745 (.ZN(n2201), 
	.B2(FE_OFN44_n3128), 
	.B1(n2718), 
	.A2(n2719), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1746 (.ZN(n2202), 
	.B2(FE_OFN44_n3128), 
	.B1(n2719), 
	.A2(n2720), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1747 (.ZN(n2203), 
	.B2(FE_OFN44_n3128), 
	.B1(n2720), 
	.A2(n2721), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1748 (.ZN(n2204), 
	.B2(FE_OFN44_n3128), 
	.B1(n2721), 
	.A2(n2722), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1749 (.ZN(n2205), 
	.B2(FE_OFN44_n3128), 
	.B1(n2722), 
	.A2(n2723), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1750 (.ZN(n2206), 
	.B2(FE_OFN44_n3128), 
	.B1(n2723), 
	.A2(n2724), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1751 (.ZN(n2207), 
	.B2(FE_OFN44_n3128), 
	.B1(n2724), 
	.A2(n2725), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1752 (.ZN(n2208), 
	.B2(FE_OFN44_n3128), 
	.B1(n2725), 
	.A2(n2726), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U1753 (.ZN(n2209), 
	.B2(FE_OFN44_n3128), 
	.B1(n2726), 
	.A2(n2727), 
	.A1(FE_OFN43_n3112));
   XNOR2_X1 U1754 (.ZN(n2696), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[31]));
   XNOR2_X1 U1755 (.ZN(n2697), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U1756 (.ZN(n2698), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[29]));
   XNOR2_X1 U1757 (.ZN(n2699), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1758 (.ZN(n2700), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1759 (.ZN(n2701), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1760 (.ZN(n2702), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[25]));
   XNOR2_X1 U1761 (.ZN(n2703), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1762 (.ZN(n2704), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1763 (.ZN(n2705), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1764 (.ZN(n2706), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1765 (.ZN(n2707), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1766 (.ZN(n2708), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[19]));
   XNOR2_X1 U1767 (.ZN(n2709), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1768 (.ZN(n2710), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[17]));
   XNOR2_X1 U1769 (.ZN(n2711), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[16]));
   XNOR2_X1 U1770 (.ZN(n2712), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[15]));
   XNOR2_X1 U1771 (.ZN(n2713), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[14]));
   XNOR2_X1 U1772 (.ZN(n2714), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1773 (.ZN(n2715), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1774 (.ZN(n2716), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1775 (.ZN(n2717), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1776 (.ZN(n2718), 
	.B(FE_OFN127_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(b[9]));
   XNOR2_X1 U1777 (.ZN(n2719), 
	.B(a[21]), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1778 (.ZN(n2720), 
	.B(a[21]), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1779 (.ZN(n2721), 
	.B(a[21]), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1780 (.ZN(n2722), 
	.B(a[21]), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1781 (.ZN(n2723), 
	.B(a[21]), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1782 (.ZN(n2724), 
	.B(a[21]), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1783 (.ZN(n2725), 
	.B(a[21]), 
	.A(b[2]));
   XNOR2_X1 U1784 (.ZN(n2726), 
	.B(a[21]), 
	.A(b[1]));
   XNOR2_X1 U1785 (.ZN(n2727), 
	.B(a[21]), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1786 (.ZN(n2009), 
	.B2(FE_OFN46_n3129), 
	.B1(n2761), 
	.A2(n3145), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1788 (.ZN(n2212), 
	.B2(FE_OFN46_n3129), 
	.B1(n2730), 
	.A2(n2731), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1789 (.ZN(n2213), 
	.B2(FE_OFN46_n3129), 
	.B1(n2731), 
	.A2(n2732), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1790 (.ZN(n2214), 
	.B2(FE_OFN46_n3129), 
	.B1(n2732), 
	.A2(n2733), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1791 (.ZN(n2215), 
	.B2(FE_OFN46_n3129), 
	.B1(n2733), 
	.A2(n2734), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1792 (.ZN(n2216), 
	.B2(FE_OFN46_n3129), 
	.B1(n2734), 
	.A2(n2735), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1793 (.ZN(n2217), 
	.B2(FE_OFN46_n3129), 
	.B1(n2735), 
	.A2(n2736), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1794 (.ZN(n2218), 
	.B2(FE_OFN46_n3129), 
	.B1(n2736), 
	.A2(n2737), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1795 (.ZN(n2219), 
	.B2(FE_OFN46_n3129), 
	.B1(n2737), 
	.A2(n2738), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1796 (.ZN(n2220), 
	.B2(FE_OFN46_n3129), 
	.B1(n2738), 
	.A2(n2739), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1797 (.ZN(n2221), 
	.B2(FE_OFN46_n3129), 
	.B1(n2739), 
	.A2(n2740), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1798 (.ZN(n2222), 
	.B2(FE_OFN46_n3129), 
	.B1(n2740), 
	.A2(n2741), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1799 (.ZN(n2223), 
	.B2(FE_OFN46_n3129), 
	.B1(n2741), 
	.A2(n2742), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1800 (.ZN(n2224), 
	.B2(FE_OFN46_n3129), 
	.B1(n2742), 
	.A2(n2743), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1801 (.ZN(n2225), 
	.B2(FE_OFN46_n3129), 
	.B1(n2743), 
	.A2(n2744), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1802 (.ZN(n2226), 
	.B2(FE_OFN46_n3129), 
	.B1(n2744), 
	.A2(n2745), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1803 (.ZN(n2227), 
	.B2(FE_OFN46_n3129), 
	.B1(n2745), 
	.A2(n2746), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1804 (.ZN(n2228), 
	.B2(FE_OFN46_n3129), 
	.B1(n2746), 
	.A2(n2747), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1805 (.ZN(n2229), 
	.B2(FE_OFN46_n3129), 
	.B1(n2747), 
	.A2(n2748), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1806 (.ZN(n2230), 
	.B2(FE_OFN46_n3129), 
	.B1(n2748), 
	.A2(n2749), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1807 (.ZN(n2231), 
	.B2(FE_OFN46_n3129), 
	.B1(n2749), 
	.A2(n2750), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1808 (.ZN(n2232), 
	.B2(FE_OFN46_n3129), 
	.B1(n2750), 
	.A2(n2751), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1809 (.ZN(n2233), 
	.B2(FE_OFN46_n3129), 
	.B1(n2751), 
	.A2(n2752), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1810 (.ZN(n2234), 
	.B2(FE_OFN46_n3129), 
	.B1(n2752), 
	.A2(n2753), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1811 (.ZN(n2235), 
	.B2(FE_OFN46_n3129), 
	.B1(n2753), 
	.A2(n2754), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1812 (.ZN(n2236), 
	.B2(FE_OFN46_n3129), 
	.B1(n2754), 
	.A2(n2755), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1813 (.ZN(n2237), 
	.B2(FE_OFN46_n3129), 
	.B1(n2755), 
	.A2(n2756), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1814 (.ZN(n2238), 
	.B2(FE_OFN46_n3129), 
	.B1(n2756), 
	.A2(n2757), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1815 (.ZN(n2239), 
	.B2(FE_OFN46_n3129), 
	.B1(n2757), 
	.A2(n2758), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1816 (.ZN(n2240), 
	.B2(FE_OFN46_n3129), 
	.B1(n2758), 
	.A2(n2759), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U1817 (.ZN(n2241), 
	.B2(FE_OFN46_n3129), 
	.B1(n2759), 
	.A2(n2760), 
	.A1(FE_OFN45_n3113));
   XNOR2_X1 U1818 (.ZN(n2729), 
	.B(a[19]), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U1819 (.ZN(n2730), 
	.B(a[19]), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U1820 (.ZN(n2731), 
	.B(a[19]), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U1821 (.ZN(n2732), 
	.B(a[19]), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1822 (.ZN(n2733), 
	.B(a[19]), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1823 (.ZN(n2734), 
	.B(a[19]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1824 (.ZN(n2735), 
	.B(a[19]), 
	.A(b[25]));
   XNOR2_X1 U1825 (.ZN(n2736), 
	.B(a[19]), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1826 (.ZN(n2737), 
	.B(a[19]), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1827 (.ZN(n2738), 
	.B(a[19]), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1828 (.ZN(n2739), 
	.B(a[19]), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1829 (.ZN(n2740), 
	.B(a[19]), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1830 (.ZN(n2741), 
	.B(a[19]), 
	.A(b[19]));
   XNOR2_X1 U1831 (.ZN(n2742), 
	.B(a[19]), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1832 (.ZN(n2743), 
	.B(a[19]), 
	.A(b[17]));
   XNOR2_X1 U1833 (.ZN(n2744), 
	.B(a[19]), 
	.A(b[16]));
   XNOR2_X1 U1834 (.ZN(n2745), 
	.B(a[19]), 
	.A(b[15]));
   XNOR2_X1 U1835 (.ZN(n2746), 
	.B(a[19]), 
	.A(b[14]));
   XNOR2_X1 U1836 (.ZN(n2747), 
	.B(a[19]), 
	.A(b[13]));
   XNOR2_X1 U1837 (.ZN(n2748), 
	.B(a[19]), 
	.A(b[12]));
   XNOR2_X1 U1838 (.ZN(n2749), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1839 (.ZN(n2750), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1840 (.ZN(n2751), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U1841 (.ZN(n2752), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1842 (.ZN(n2753), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1843 (.ZN(n2754), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1844 (.ZN(n2755), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1845 (.ZN(n2756), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1846 (.ZN(n2757), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1847 (.ZN(n2758), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(b[2]));
   XNOR2_X1 U1848 (.ZN(n2759), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(b[1]));
   XNOR2_X1 U1849 (.ZN(n2760), 
	.B(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1850 (.ZN(n2010), 
	.B2(FE_OFN48_n3130), 
	.B1(n2794), 
	.A2(n3146), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1852 (.ZN(n2244), 
	.B2(FE_OFN48_n3130), 
	.B1(n2763), 
	.A2(n2764), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1853 (.ZN(n2245), 
	.B2(FE_OFN48_n3130), 
	.B1(n2764), 
	.A2(n2765), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1854 (.ZN(n2246), 
	.B2(FE_OFN48_n3130), 
	.B1(n2765), 
	.A2(n2766), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1855 (.ZN(n2247), 
	.B2(FE_OFN48_n3130), 
	.B1(n2766), 
	.A2(n2767), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1856 (.ZN(n2248), 
	.B2(FE_OFN48_n3130), 
	.B1(n2767), 
	.A2(n2768), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1857 (.ZN(n2249), 
	.B2(FE_OFN48_n3130), 
	.B1(n2768), 
	.A2(n2769), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1858 (.ZN(n2250), 
	.B2(FE_OFN48_n3130), 
	.B1(n2769), 
	.A2(n2770), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1859 (.ZN(n2251), 
	.B2(FE_OFN48_n3130), 
	.B1(n2770), 
	.A2(n2771), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1860 (.ZN(n2252), 
	.B2(FE_OFN48_n3130), 
	.B1(n2771), 
	.A2(n2772), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1861 (.ZN(n2253), 
	.B2(FE_OFN48_n3130), 
	.B1(n2772), 
	.A2(n2773), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1862 (.ZN(n2254), 
	.B2(FE_OFN48_n3130), 
	.B1(n2773), 
	.A2(n2774), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1863 (.ZN(n2255), 
	.B2(FE_OFN48_n3130), 
	.B1(n2774), 
	.A2(n2775), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1864 (.ZN(n2256), 
	.B2(FE_OFN48_n3130), 
	.B1(n2775), 
	.A2(n2776), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1865 (.ZN(n2257), 
	.B2(FE_OFN48_n3130), 
	.B1(n2776), 
	.A2(n2777), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1866 (.ZN(n2258), 
	.B2(FE_OFN48_n3130), 
	.B1(n2777), 
	.A2(n2778), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1867 (.ZN(n2259), 
	.B2(FE_OFN48_n3130), 
	.B1(n2778), 
	.A2(n2779), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1868 (.ZN(n2260), 
	.B2(FE_OFN48_n3130), 
	.B1(n2779), 
	.A2(n2780), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1869 (.ZN(n2261), 
	.B2(FE_OFN48_n3130), 
	.B1(n2780), 
	.A2(n2781), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1870 (.ZN(n2262), 
	.B2(FE_OFN48_n3130), 
	.B1(n2781), 
	.A2(n2782), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1871 (.ZN(n2263), 
	.B2(FE_OFN48_n3130), 
	.B1(n2782), 
	.A2(n2783), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1872 (.ZN(n2264), 
	.B2(FE_OFN48_n3130), 
	.B1(n2783), 
	.A2(n2784), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1873 (.ZN(n2265), 
	.B2(FE_OFN48_n3130), 
	.B1(n2784), 
	.A2(n2785), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1874 (.ZN(n2266), 
	.B2(FE_OFN48_n3130), 
	.B1(n2785), 
	.A2(n2786), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1875 (.ZN(n2267), 
	.B2(FE_OFN48_n3130), 
	.B1(n2786), 
	.A2(n2787), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1876 (.ZN(n2268), 
	.B2(FE_OFN48_n3130), 
	.B1(n2787), 
	.A2(n2788), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1877 (.ZN(n2269), 
	.B2(FE_OFN48_n3130), 
	.B1(n2788), 
	.A2(n2789), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1878 (.ZN(n2270), 
	.B2(FE_OFN48_n3130), 
	.B1(n2789), 
	.A2(n2790), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1879 (.ZN(n2271), 
	.B2(FE_OFN48_n3130), 
	.B1(n2790), 
	.A2(n2791), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1880 (.ZN(n2272), 
	.B2(FE_OFN48_n3130), 
	.B1(n2791), 
	.A2(n2792), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U1881 (.ZN(n2273), 
	.B2(FE_OFN48_n3130), 
	.B1(n2792), 
	.A2(n2793), 
	.A1(FE_OFN47_n3114));
   XNOR2_X1 U1882 (.ZN(n2762), 
	.B(a[17]), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U1883 (.ZN(n2763), 
	.B(a[17]), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U1884 (.ZN(n2764), 
	.B(a[17]), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U1885 (.ZN(n2765), 
	.B(a[17]), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1886 (.ZN(n2766), 
	.B(a[17]), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1887 (.ZN(n2767), 
	.B(a[17]), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1888 (.ZN(n2768), 
	.B(a[17]), 
	.A(b[25]));
   XNOR2_X1 U1889 (.ZN(n2769), 
	.B(a[17]), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1890 (.ZN(n2770), 
	.B(a[17]), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1891 (.ZN(n2771), 
	.B(a[17]), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1892 (.ZN(n2772), 
	.B(a[17]), 
	.A(b[21]));
   XNOR2_X1 U1893 (.ZN(n2773), 
	.B(a[17]), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1894 (.ZN(n2774), 
	.B(a[17]), 
	.A(b[19]));
   XNOR2_X1 U1895 (.ZN(n2775), 
	.B(a[17]), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1896 (.ZN(n2776), 
	.B(a[17]), 
	.A(b[17]));
   XNOR2_X1 U1897 (.ZN(n2777), 
	.B(a[17]), 
	.A(b[16]));
   XNOR2_X1 U1898 (.ZN(n2778), 
	.B(a[17]), 
	.A(b[15]));
   XNOR2_X1 U1899 (.ZN(n2779), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(b[14]));
   XNOR2_X1 U1900 (.ZN(n2780), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(b[13]));
   XNOR2_X1 U1901 (.ZN(n2781), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1902 (.ZN(n2782), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN145_UUT_Mpath_the_mult_x_operand2_11_));
   XNOR2_X1 U1903 (.ZN(n2783), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN108_UUT_Mpath_the_mult_x_operand2_10_));
   XNOR2_X1 U1904 (.ZN(n2784), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U1905 (.ZN(n2785), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1906 (.ZN(n2786), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1907 (.ZN(n2787), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1908 (.ZN(n2788), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1909 (.ZN(n2789), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1910 (.ZN(n2790), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1911 (.ZN(n2791), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(b[2]));
   XNOR2_X1 U1912 (.ZN(n2792), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(b[1]));
   XNOR2_X1 U1913 (.ZN(n2793), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(FE_OFN106_UUT_Mpath_the_mult_x_operand2_0_));
   OAI22_X1 U1914 (.ZN(n2011), 
	.B2(n3131), 
	.B1(n2827), 
	.A2(FE_PT1_n477), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1916 (.ZN(n2276), 
	.B2(FE_OFN52_n3131), 
	.B1(n2796), 
	.A2(n2797), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1917 (.ZN(n2277), 
	.B2(FE_OFN52_n3131), 
	.B1(n2797), 
	.A2(n2798), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1918 (.ZN(n2278), 
	.B2(FE_OFN52_n3131), 
	.B1(n2798), 
	.A2(n2799), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1919 (.ZN(n2279), 
	.B2(FE_OFN52_n3131), 
	.B1(n2799), 
	.A2(n2800), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1920 (.ZN(n2280), 
	.B2(FE_OFN52_n3131), 
	.B1(n2800), 
	.A2(n2801), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1921 (.ZN(n2281), 
	.B2(FE_OFN52_n3131), 
	.B1(n2801), 
	.A2(n2802), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1922 (.ZN(n2282), 
	.B2(FE_OFN52_n3131), 
	.B1(n2802), 
	.A2(n2803), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1923 (.ZN(n2283), 
	.B2(FE_OFN52_n3131), 
	.B1(n2803), 
	.A2(n2804), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1924 (.ZN(n2284), 
	.B2(FE_OFN52_n3131), 
	.B1(n2804), 
	.A2(n2805), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1925 (.ZN(n2285), 
	.B2(FE_OFN52_n3131), 
	.B1(n2805), 
	.A2(n2806), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1926 (.ZN(n2286), 
	.B2(FE_OFN52_n3131), 
	.B1(n2806), 
	.A2(n2807), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1927 (.ZN(n2287), 
	.B2(FE_OFN52_n3131), 
	.B1(n2807), 
	.A2(n2808), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1928 (.ZN(n2288), 
	.B2(FE_OFN52_n3131), 
	.B1(n2808), 
	.A2(n2809), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1929 (.ZN(n2289), 
	.B2(FE_OFN52_n3131), 
	.B1(n2809), 
	.A2(n2810), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1930 (.ZN(n2290), 
	.B2(FE_OFN52_n3131), 
	.B1(n2810), 
	.A2(n2811), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1931 (.ZN(n2291), 
	.B2(FE_OFN52_n3131), 
	.B1(n2811), 
	.A2(n2812), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1932 (.ZN(n2292), 
	.B2(FE_OFN52_n3131), 
	.B1(n2812), 
	.A2(n2813), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1933 (.ZN(n2293), 
	.B2(FE_OFN52_n3131), 
	.B1(n2813), 
	.A2(n2814), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1934 (.ZN(n2294), 
	.B2(FE_OFN52_n3131), 
	.B1(n2814), 
	.A2(n2815), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1935 (.ZN(n2295), 
	.B2(FE_OFN52_n3131), 
	.B1(n2815), 
	.A2(n2816), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1936 (.ZN(n2296), 
	.B2(FE_OFN52_n3131), 
	.B1(n2816), 
	.A2(n2817), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1937 (.ZN(n2297), 
	.B2(FE_OFN52_n3131), 
	.B1(n2817), 
	.A2(n2818), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1938 (.ZN(n2298), 
	.B2(FE_OFN52_n3131), 
	.B1(n2818), 
	.A2(n2819), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1939 (.ZN(n2299), 
	.B2(FE_OFN52_n3131), 
	.B1(n2819), 
	.A2(n2820), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1940 (.ZN(n2300), 
	.B2(FE_OFN52_n3131), 
	.B1(n2820), 
	.A2(n2821), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1941 (.ZN(n2301), 
	.B2(FE_OFN52_n3131), 
	.B1(n2821), 
	.A2(n2822), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1942 (.ZN(n2302), 
	.B2(FE_OFN52_n3131), 
	.B1(n2822), 
	.A2(n2823), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1943 (.ZN(n2303), 
	.B2(FE_OFN52_n3131), 
	.B1(n2823), 
	.A2(n2824), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1944 (.ZN(n2304), 
	.B2(FE_OFN52_n3131), 
	.B1(n2824), 
	.A2(n2825), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U1945 (.ZN(n2305), 
	.B2(FE_OFN52_n3131), 
	.B1(n2825), 
	.A2(n2826), 
	.A1(FE_OFN51_n3115));
   XNOR2_X1 U1946 (.ZN(n2795), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U1947 (.ZN(n2796), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U1948 (.ZN(n2797), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U1949 (.ZN(n2798), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN115_UUT_Mpath_the_mult_x_operand2_28_));
   XNOR2_X1 U1950 (.ZN(n2799), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN116_UUT_Mpath_the_mult_x_operand2_27_));
   XNOR2_X1 U1951 (.ZN(n2800), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN119_UUT_Mpath_the_mult_x_operand2_26_));
   XNOR2_X1 U1952 (.ZN(n2801), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[25]));
   XNOR2_X1 U1953 (.ZN(n2802), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN123_UUT_Mpath_the_mult_x_operand2_24_));
   XNOR2_X1 U1954 (.ZN(n2803), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN110_UUT_Mpath_the_mult_x_operand2_23_));
   XNOR2_X1 U1955 (.ZN(n2804), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN124_UUT_Mpath_the_mult_x_operand2_22_));
   XNOR2_X1 U1956 (.ZN(n2805), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U1957 (.ZN(n2806), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN128_UUT_Mpath_the_mult_x_operand2_20_));
   XNOR2_X1 U1958 (.ZN(n2807), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[19]));
   XNOR2_X1 U1959 (.ZN(n2808), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN132_UUT_Mpath_the_mult_x_operand2_18_));
   XNOR2_X1 U1960 (.ZN(n2809), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[17]));
   XNOR2_X1 U1961 (.ZN(n2810), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[16]));
   XNOR2_X1 U1962 (.ZN(n2811), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[15]));
   XNOR2_X1 U1963 (.ZN(n2812), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[14]));
   XNOR2_X1 U1964 (.ZN(n2813), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U1965 (.ZN(n2814), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN144_UUT_Mpath_the_mult_x_operand2_12_));
   XNOR2_X1 U1966 (.ZN(n2815), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[11]));
   XNOR2_X1 U1967 (.ZN(n2816), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(b[10]));
   XNOR2_X1 U1968 (.ZN(n2817), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U1969 (.ZN(n2818), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN109_UUT_Mpath_the_mult_x_operand2_8_));
   XNOR2_X1 U1970 (.ZN(n2819), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN151_UUT_Mpath_the_mult_x_operand2_7_));
   XNOR2_X1 U1971 (.ZN(n2820), 
	.B(FE_OFN139_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(FE_OFN154_UUT_Mpath_the_mult_x_operand2_6_));
   XNOR2_X1 U1972 (.ZN(n2821), 
	.B(a[15]), 
	.A(FE_OFN155_UUT_Mpath_the_mult_x_operand2_5_));
   XNOR2_X1 U1973 (.ZN(n2822), 
	.B(a[15]), 
	.A(FE_OFN158_UUT_Mpath_the_mult_x_operand2_4_));
   XNOR2_X1 U1974 (.ZN(n2823), 
	.B(a[15]), 
	.A(FE_OFN161_UUT_Mpath_the_mult_x_operand2_3_));
   XNOR2_X1 U1975 (.ZN(n2824), 
	.B(a[15]), 
	.A(b[2]));
   XNOR2_X1 U1976 (.ZN(n2825), 
	.B(a[15]), 
	.A(b[1]));
   XNOR2_X1 U1977 (.ZN(n2826), 
	.B(a[15]), 
	.A(b[0]));
   OAI22_X1 U1978 (.ZN(n2012), 
	.B2(FE_OFN58_n3132), 
	.B1(n2860), 
	.A2(n531), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1980 (.ZN(n2308), 
	.B2(FE_OFN58_n3132), 
	.B1(n2829), 
	.A2(n2830), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1981 (.ZN(n2309), 
	.B2(FE_OFN58_n3132), 
	.B1(n2830), 
	.A2(n2831), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1982 (.ZN(n2310), 
	.B2(FE_OFN58_n3132), 
	.B1(n2831), 
	.A2(n2832), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1983 (.ZN(n2311), 
	.B2(FE_OFN58_n3132), 
	.B1(n2832), 
	.A2(n2833), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1984 (.ZN(n2312), 
	.B2(FE_OFN58_n3132), 
	.B1(n2833), 
	.A2(n2834), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1985 (.ZN(n2313), 
	.B2(FE_OFN58_n3132), 
	.B1(n2834), 
	.A2(n2835), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1986 (.ZN(n2314), 
	.B2(FE_OFN58_n3132), 
	.B1(n2835), 
	.A2(n2836), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1987 (.ZN(n2315), 
	.B2(FE_OFN58_n3132), 
	.B1(n2836), 
	.A2(n2837), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1988 (.ZN(n2316), 
	.B2(FE_OFN58_n3132), 
	.B1(n2837), 
	.A2(n2838), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1989 (.ZN(n2317), 
	.B2(FE_OFN58_n3132), 
	.B1(n2838), 
	.A2(n2839), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1990 (.ZN(n2318), 
	.B2(FE_OFN58_n3132), 
	.B1(n2839), 
	.A2(n2840), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1991 (.ZN(n2319), 
	.B2(FE_OFN58_n3132), 
	.B1(n2840), 
	.A2(n2841), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1992 (.ZN(n2320), 
	.B2(FE_OFN58_n3132), 
	.B1(n2841), 
	.A2(n2842), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1993 (.ZN(n2321), 
	.B2(FE_OFN58_n3132), 
	.B1(n2842), 
	.A2(n2843), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1994 (.ZN(n2322), 
	.B2(FE_OFN58_n3132), 
	.B1(n2843), 
	.A2(n2844), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1995 (.ZN(n2323), 
	.B2(FE_OFN58_n3132), 
	.B1(n2844), 
	.A2(n2845), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1996 (.ZN(n2324), 
	.B2(FE_OFN58_n3132), 
	.B1(n2845), 
	.A2(n2846), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1997 (.ZN(n2325), 
	.B2(FE_OFN58_n3132), 
	.B1(n2846), 
	.A2(n2847), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1998 (.ZN(n2326), 
	.B2(FE_OFN58_n3132), 
	.B1(n2847), 
	.A2(n2848), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U1999 (.ZN(n2327), 
	.B2(FE_OFN58_n3132), 
	.B1(n2848), 
	.A2(n2849), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2000 (.ZN(n2328), 
	.B2(FE_OFN58_n3132), 
	.B1(n2849), 
	.A2(n2850), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2001 (.ZN(n2329), 
	.B2(FE_OFN58_n3132), 
	.B1(n2850), 
	.A2(n2851), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2002 (.ZN(n2330), 
	.B2(FE_OFN58_n3132), 
	.B1(n2851), 
	.A2(n2852), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2003 (.ZN(n2331), 
	.B2(FE_OFN58_n3132), 
	.B1(n2852), 
	.A2(n2853), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2004 (.ZN(n2332), 
	.B2(FE_OFN58_n3132), 
	.B1(n2853), 
	.A2(n2854), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2005 (.ZN(n2333), 
	.B2(FE_OFN58_n3132), 
	.B1(n2854), 
	.A2(n2855), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2006 (.ZN(n2334), 
	.B2(FE_OFN58_n3132), 
	.B1(n2855), 
	.A2(n2856), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2007 (.ZN(n2335), 
	.B2(FE_OFN58_n3132), 
	.B1(n2856), 
	.A2(n2857), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2008 (.ZN(n2336), 
	.B2(FE_OFN58_n3132), 
	.B1(n2857), 
	.A2(n2858), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2009 (.ZN(n2337), 
	.B2(FE_OFN58_n3132), 
	.B1(n2858), 
	.A2(n2859), 
	.A1(FE_OFN55_n3116));
   XNOR2_X1 U2010 (.ZN(n2828), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U2011 (.ZN(n2829), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U2012 (.ZN(n2830), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2013 (.ZN(n2831), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[28]));
   XNOR2_X1 U2014 (.ZN(n2832), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[27]));
   XNOR2_X1 U2015 (.ZN(n2833), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[26]));
   XNOR2_X1 U2016 (.ZN(n2834), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[25]));
   XNOR2_X1 U2017 (.ZN(n2835), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[24]));
   XNOR2_X1 U2018 (.ZN(n2836), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[23]));
   XNOR2_X1 U2019 (.ZN(n2837), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[22]));
   XNOR2_X1 U2020 (.ZN(n2838), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN125_UUT_Mpath_the_mult_x_operand2_21_));
   XNOR2_X1 U2021 (.ZN(n2839), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[20]));
   XNOR2_X1 U2022 (.ZN(n2840), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[19]));
   XNOR2_X1 U2023 (.ZN(n2841), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[18]));
   XNOR2_X1 U2024 (.ZN(n2842), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[17]));
   XNOR2_X1 U2025 (.ZN(n2843), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[16]));
   XNOR2_X1 U2026 (.ZN(n2844), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[15]));
   XNOR2_X1 U2027 (.ZN(n2845), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[14]));
   XNOR2_X1 U2028 (.ZN(n2846), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN141_UUT_Mpath_the_mult_x_operand2_13_));
   XNOR2_X1 U2029 (.ZN(n2847), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[12]));
   XNOR2_X1 U2030 (.ZN(n2848), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[11]));
   XNOR2_X1 U2031 (.ZN(n2849), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[10]));
   XNOR2_X1 U2032 (.ZN(n2850), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U2033 (.ZN(n2851), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[8]));
   XNOR2_X1 U2034 (.ZN(n2852), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[7]));
   XNOR2_X1 U2035 (.ZN(n2853), 
	.B(FE_OFN143_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(b[6]));
   XNOR2_X1 U2036 (.ZN(n2854), 
	.B(a[13]), 
	.A(b[5]));
   XNOR2_X1 U2037 (.ZN(n2855), 
	.B(a[13]), 
	.A(b[4]));
   XNOR2_X1 U2038 (.ZN(n2856), 
	.B(a[13]), 
	.A(b[3]));
   XNOR2_X1 U2039 (.ZN(n2857), 
	.B(a[13]), 
	.A(b[2]));
   XNOR2_X1 U2040 (.ZN(n2858), 
	.B(a[13]), 
	.A(b[1]));
   XNOR2_X1 U2041 (.ZN(n2859), 
	.B(a[13]), 
	.A(b[0]));
   OAI22_X1 U2042 (.ZN(n2013), 
	.B2(FE_OFN64_n3133), 
	.B1(n2893), 
	.A2(FE_PT1_n582), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2044 (.ZN(n2340), 
	.B2(FE_OFN64_n3133), 
	.B1(n2862), 
	.A2(n2863), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2045 (.ZN(n2341), 
	.B2(FE_OFN64_n3133), 
	.B1(n2863), 
	.A2(n2864), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2046 (.ZN(n2342), 
	.B2(FE_OFN64_n3133), 
	.B1(n2864), 
	.A2(n2865), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2047 (.ZN(n2343), 
	.B2(FE_OFN64_n3133), 
	.B1(n2865), 
	.A2(n2866), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2048 (.ZN(n2344), 
	.B2(FE_OFN64_n3133), 
	.B1(n2866), 
	.A2(n2867), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2049 (.ZN(n2345), 
	.B2(FE_OFN64_n3133), 
	.B1(n2867), 
	.A2(n2868), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2050 (.ZN(n2346), 
	.B2(FE_OFN64_n3133), 
	.B1(n2868), 
	.A2(n2869), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2051 (.ZN(n2347), 
	.B2(FE_OFN64_n3133), 
	.B1(n2869), 
	.A2(n2870), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2052 (.ZN(n2348), 
	.B2(FE_OFN64_n3133), 
	.B1(n2870), 
	.A2(n2871), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2053 (.ZN(n2349), 
	.B2(FE_OFN64_n3133), 
	.B1(n2871), 
	.A2(n2872), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2054 (.ZN(n2350), 
	.B2(FE_OFN64_n3133), 
	.B1(n2872), 
	.A2(n2873), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2055 (.ZN(n2351), 
	.B2(FE_OFN64_n3133), 
	.B1(n2873), 
	.A2(n2874), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2056 (.ZN(n2352), 
	.B2(FE_OFN64_n3133), 
	.B1(n2874), 
	.A2(n2875), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2057 (.ZN(n2353), 
	.B2(FE_OFN64_n3133), 
	.B1(n2875), 
	.A2(n2876), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2058 (.ZN(n2354), 
	.B2(FE_OFN64_n3133), 
	.B1(n2876), 
	.A2(n2877), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2059 (.ZN(n2355), 
	.B2(FE_OFN64_n3133), 
	.B1(n2877), 
	.A2(n2878), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2060 (.ZN(n2356), 
	.B2(FE_OFN64_n3133), 
	.B1(n2878), 
	.A2(n2879), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2061 (.ZN(n2357), 
	.B2(FE_OFN64_n3133), 
	.B1(n2879), 
	.A2(n2880), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2062 (.ZN(n2358), 
	.B2(FE_OFN64_n3133), 
	.B1(n2880), 
	.A2(n2881), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2063 (.ZN(n2359), 
	.B2(FE_OFN64_n3133), 
	.B1(n2881), 
	.A2(n2882), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2064 (.ZN(n2360), 
	.B2(FE_OFN64_n3133), 
	.B1(n2882), 
	.A2(n2883), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2065 (.ZN(n2361), 
	.B2(FE_OFN64_n3133), 
	.B1(n2883), 
	.A2(n2884), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2066 (.ZN(n2362), 
	.B2(FE_OFN64_n3133), 
	.B1(n2884), 
	.A2(n2885), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2067 (.ZN(n2363), 
	.B2(FE_OFN64_n3133), 
	.B1(n2885), 
	.A2(n2886), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2068 (.ZN(n2364), 
	.B2(FE_OFN64_n3133), 
	.B1(n2886), 
	.A2(n2887), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2069 (.ZN(n2365), 
	.B2(FE_OFN64_n3133), 
	.B1(n2887), 
	.A2(n2888), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2070 (.ZN(n2366), 
	.B2(FE_OFN64_n3133), 
	.B1(n2888), 
	.A2(n2889), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2071 (.ZN(n2367), 
	.B2(FE_OFN64_n3133), 
	.B1(n2889), 
	.A2(n2890), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2072 (.ZN(n2368), 
	.B2(FE_OFN64_n3133), 
	.B1(n2890), 
	.A2(n2891), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2073 (.ZN(n2369), 
	.B2(FE_OFN64_n3133), 
	.B1(n2891), 
	.A2(n2892), 
	.A1(FE_OFN61_n3117));
   XNOR2_X1 U2074 (.ZN(n2861), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U2075 (.ZN(n2862), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U2076 (.ZN(n2863), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2077 (.ZN(n2864), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[28]));
   XNOR2_X1 U2078 (.ZN(n2865), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[27]));
   XNOR2_X1 U2079 (.ZN(n2866), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[26]));
   XNOR2_X1 U2080 (.ZN(n2867), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[25]));
   XNOR2_X1 U2081 (.ZN(n2868), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[24]));
   XNOR2_X1 U2082 (.ZN(n2869), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[23]));
   XNOR2_X1 U2083 (.ZN(n2870), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[22]));
   XNOR2_X1 U2084 (.ZN(n2871), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[21]));
   XNOR2_X1 U2085 (.ZN(n2872), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[20]));
   XNOR2_X1 U2086 (.ZN(n2873), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[19]));
   XNOR2_X1 U2087 (.ZN(n2874), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[18]));
   XNOR2_X1 U2088 (.ZN(n2875), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[17]));
   XNOR2_X1 U2089 (.ZN(n2876), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[16]));
   XNOR2_X1 U2090 (.ZN(n2877), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[15]));
   XNOR2_X1 U2091 (.ZN(n2878), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[14]));
   XNOR2_X1 U2092 (.ZN(n2879), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[13]));
   XNOR2_X1 U2093 (.ZN(n2880), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[12]));
   XNOR2_X1 U2094 (.ZN(n2881), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[11]));
   XNOR2_X1 U2095 (.ZN(n2882), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[10]));
   XNOR2_X1 U2096 (.ZN(n2883), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U2097 (.ZN(n2884), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[8]));
   XNOR2_X1 U2098 (.ZN(n2885), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[7]));
   XNOR2_X1 U2099 (.ZN(n2886), 
	.B(FE_OFN147_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(b[6]));
   XNOR2_X1 U2100 (.ZN(n2887), 
	.B(a[11]), 
	.A(b[5]));
   XNOR2_X1 U2101 (.ZN(n2888), 
	.B(a[11]), 
	.A(b[4]));
   XNOR2_X1 U2102 (.ZN(n2889), 
	.B(a[11]), 
	.A(b[3]));
   XNOR2_X1 U2103 (.ZN(n2890), 
	.B(a[11]), 
	.A(b[2]));
   XNOR2_X1 U2104 (.ZN(n2891), 
	.B(a[11]), 
	.A(b[1]));
   XNOR2_X1 U2105 (.ZN(n2892), 
	.B(a[11]), 
	.A(b[0]));
   OAI22_X1 U2106 (.ZN(n2014), 
	.B2(FE_OFN66_n3134), 
	.B1(n2926), 
	.A2(FE_PT1_n617), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2108 (.ZN(n2372), 
	.B2(FE_OFN66_n3134), 
	.B1(n2895), 
	.A2(n2896), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2109 (.ZN(n2373), 
	.B2(FE_OFN66_n3134), 
	.B1(n2896), 
	.A2(n2897), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2110 (.ZN(n2374), 
	.B2(FE_OFN66_n3134), 
	.B1(n2897), 
	.A2(n2898), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2111 (.ZN(n2375), 
	.B2(FE_OFN66_n3134), 
	.B1(n2898), 
	.A2(n2899), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2112 (.ZN(n2376), 
	.B2(FE_OFN66_n3134), 
	.B1(n2899), 
	.A2(n2900), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2113 (.ZN(n2377), 
	.B2(FE_OFN66_n3134), 
	.B1(n2900), 
	.A2(n2901), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2114 (.ZN(n2378), 
	.B2(FE_OFN66_n3134), 
	.B1(n2901), 
	.A2(n2902), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2115 (.ZN(n2379), 
	.B2(FE_OFN66_n3134), 
	.B1(n2902), 
	.A2(n2903), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2116 (.ZN(n2380), 
	.B2(FE_OFN66_n3134), 
	.B1(n2903), 
	.A2(n2904), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2117 (.ZN(n2381), 
	.B2(FE_OFN66_n3134), 
	.B1(n2904), 
	.A2(n2905), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2118 (.ZN(n2382), 
	.B2(FE_OFN66_n3134), 
	.B1(n2905), 
	.A2(n2906), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2119 (.ZN(n2383), 
	.B2(FE_OFN66_n3134), 
	.B1(n2906), 
	.A2(n2907), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2120 (.ZN(n2384), 
	.B2(FE_OFN66_n3134), 
	.B1(n2907), 
	.A2(n2908), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2121 (.ZN(n2385), 
	.B2(FE_OFN66_n3134), 
	.B1(n2908), 
	.A2(n2909), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2122 (.ZN(n2386), 
	.B2(FE_OFN66_n3134), 
	.B1(n2909), 
	.A2(n2910), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2123 (.ZN(n2387), 
	.B2(FE_OFN66_n3134), 
	.B1(n2910), 
	.A2(n2911), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2124 (.ZN(n2388), 
	.B2(FE_OFN66_n3134), 
	.B1(n2911), 
	.A2(n2912), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2125 (.ZN(n2389), 
	.B2(FE_OFN66_n3134), 
	.B1(n2912), 
	.A2(n2913), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2126 (.ZN(n2390), 
	.B2(FE_OFN66_n3134), 
	.B1(n2913), 
	.A2(n2914), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2127 (.ZN(n2391), 
	.B2(FE_OFN66_n3134), 
	.B1(n2914), 
	.A2(n2915), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2128 (.ZN(n2392), 
	.B2(FE_OFN66_n3134), 
	.B1(n2915), 
	.A2(n2916), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2129 (.ZN(n2393), 
	.B2(FE_OFN66_n3134), 
	.B1(n2916), 
	.A2(n2917), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2130 (.ZN(n2394), 
	.B2(FE_OFN66_n3134), 
	.B1(n2917), 
	.A2(n2918), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2131 (.ZN(n2395), 
	.B2(FE_OFN66_n3134), 
	.B1(n2918), 
	.A2(n2919), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2132 (.ZN(n2396), 
	.B2(FE_OFN66_n3134), 
	.B1(n2919), 
	.A2(n2920), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2133 (.ZN(n2397), 
	.B2(FE_OFN66_n3134), 
	.B1(n2920), 
	.A2(n2921), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2134 (.ZN(n2398), 
	.B2(FE_OFN66_n3134), 
	.B1(n2921), 
	.A2(n2922), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2135 (.ZN(n2399), 
	.B2(FE_OFN66_n3134), 
	.B1(n2922), 
	.A2(n2923), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2136 (.ZN(n2400), 
	.B2(FE_OFN66_n3134), 
	.B1(n2923), 
	.A2(n2924), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2137 (.ZN(n2401), 
	.B2(FE_OFN66_n3134), 
	.B1(n2924), 
	.A2(n2925), 
	.A1(FE_OFN65_n3118));
   XNOR2_X1 U2138 (.ZN(n2894), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U2139 (.ZN(n2895), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U2140 (.ZN(n2896), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2141 (.ZN(n2897), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[28]));
   XNOR2_X1 U2142 (.ZN(n2898), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[27]));
   XNOR2_X1 U2143 (.ZN(n2899), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[26]));
   XNOR2_X1 U2144 (.ZN(n2900), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[25]));
   XNOR2_X1 U2145 (.ZN(n2901), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[24]));
   XNOR2_X1 U2146 (.ZN(n2902), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[23]));
   XNOR2_X1 U2147 (.ZN(n2903), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[22]));
   XNOR2_X1 U2148 (.ZN(n2904), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[21]));
   XNOR2_X1 U2149 (.ZN(n2905), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[20]));
   XNOR2_X1 U2150 (.ZN(n2906), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[19]));
   XNOR2_X1 U2151 (.ZN(n2907), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[18]));
   XNOR2_X1 U2152 (.ZN(n2908), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[17]));
   XNOR2_X1 U2153 (.ZN(n2909), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[16]));
   XNOR2_X1 U2154 (.ZN(n2910), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[15]));
   XNOR2_X1 U2155 (.ZN(n2911), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[14]));
   XNOR2_X1 U2156 (.ZN(n2912), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[13]));
   XNOR2_X1 U2157 (.ZN(n2913), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[12]));
   XNOR2_X1 U2158 (.ZN(n2914), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[11]));
   XNOR2_X1 U2159 (.ZN(n2915), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[10]));
   XNOR2_X1 U2160 (.ZN(n2916), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U2161 (.ZN(n2917), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[8]));
   XNOR2_X1 U2162 (.ZN(n2918), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[7]));
   XNOR2_X1 U2163 (.ZN(n2919), 
	.B(FE_OFN150_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(b[6]));
   XNOR2_X1 U2164 (.ZN(n2920), 
	.B(a[9]), 
	.A(b[5]));
   XNOR2_X1 U2165 (.ZN(n2921), 
	.B(a[9]), 
	.A(b[4]));
   XNOR2_X1 U2166 (.ZN(n2922), 
	.B(a[9]), 
	.A(b[3]));
   XNOR2_X1 U2167 (.ZN(n2923), 
	.B(a[9]), 
	.A(b[2]));
   XNOR2_X1 U2168 (.ZN(n2924), 
	.B(a[9]), 
	.A(b[1]));
   XNOR2_X1 U2169 (.ZN(n2925), 
	.B(a[9]), 
	.A(b[0]));
   OAI22_X1 U2170 (.ZN(n2015), 
	.B2(FE_OFN70_n3135), 
	.B1(n2959), 
	.A2(FE_PT1_n654), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2172 (.ZN(n2404), 
	.B2(FE_OFN70_n3135), 
	.B1(n2928), 
	.A2(n2929), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2173 (.ZN(n2405), 
	.B2(FE_OFN70_n3135), 
	.B1(n2929), 
	.A2(n2930), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2174 (.ZN(n2406), 
	.B2(FE_OFN70_n3135), 
	.B1(n2930), 
	.A2(n2931), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2175 (.ZN(n2407), 
	.B2(FE_OFN70_n3135), 
	.B1(n2931), 
	.A2(n2932), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2176 (.ZN(n2408), 
	.B2(FE_OFN70_n3135), 
	.B1(n2932), 
	.A2(n2933), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2177 (.ZN(n2409), 
	.B2(FE_OFN70_n3135), 
	.B1(n2933), 
	.A2(n2934), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2178 (.ZN(n2410), 
	.B2(FE_OFN70_n3135), 
	.B1(n2934), 
	.A2(n2935), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2179 (.ZN(n2411), 
	.B2(FE_OFN70_n3135), 
	.B1(n2935), 
	.A2(n2936), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2180 (.ZN(n2412), 
	.B2(FE_OFN70_n3135), 
	.B1(n2936), 
	.A2(n2937), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2181 (.ZN(n2413), 
	.B2(FE_OFN70_n3135), 
	.B1(n2937), 
	.A2(n2938), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2182 (.ZN(n2414), 
	.B2(FE_OFN70_n3135), 
	.B1(n2938), 
	.A2(n2939), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2183 (.ZN(n2415), 
	.B2(FE_OFN70_n3135), 
	.B1(n2939), 
	.A2(n2940), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2184 (.ZN(n2416), 
	.B2(FE_OFN70_n3135), 
	.B1(n2940), 
	.A2(n2941), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2185 (.ZN(n2417), 
	.B2(FE_OFN70_n3135), 
	.B1(n2941), 
	.A2(n2942), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2186 (.ZN(n2418), 
	.B2(FE_OFN70_n3135), 
	.B1(n2942), 
	.A2(n2943), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2187 (.ZN(n2419), 
	.B2(FE_OFN70_n3135), 
	.B1(n2943), 
	.A2(n2944), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2188 (.ZN(n2420), 
	.B2(FE_OFN70_n3135), 
	.B1(n2944), 
	.A2(n2945), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2189 (.ZN(n2421), 
	.B2(FE_OFN70_n3135), 
	.B1(n2945), 
	.A2(n2946), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2190 (.ZN(n2422), 
	.B2(FE_OFN70_n3135), 
	.B1(n2946), 
	.A2(n2947), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2191 (.ZN(n2423), 
	.B2(FE_OFN70_n3135), 
	.B1(n2947), 
	.A2(n2948), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2192 (.ZN(n2424), 
	.B2(FE_OFN70_n3135), 
	.B1(n2948), 
	.A2(n2949), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2193 (.ZN(n2425), 
	.B2(FE_OFN70_n3135), 
	.B1(n2949), 
	.A2(n2950), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2194 (.ZN(n2426), 
	.B2(FE_OFN70_n3135), 
	.B1(n2950), 
	.A2(n2951), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2195 (.ZN(n2427), 
	.B2(FE_OFN70_n3135), 
	.B1(n2951), 
	.A2(n2952), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2196 (.ZN(n2428), 
	.B2(FE_OFN70_n3135), 
	.B1(n2952), 
	.A2(n2953), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2197 (.ZN(n2429), 
	.B2(FE_OFN70_n3135), 
	.B1(n2953), 
	.A2(n2954), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2198 (.ZN(n2430), 
	.B2(FE_OFN70_n3135), 
	.B1(n2954), 
	.A2(n2955), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2199 (.ZN(n2431), 
	.B2(FE_OFN70_n3135), 
	.B1(n2955), 
	.A2(n2956), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2200 (.ZN(n2432), 
	.B2(FE_OFN70_n3135), 
	.B1(n2956), 
	.A2(n2957), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2201 (.ZN(n2433), 
	.B2(FE_OFN70_n3135), 
	.B1(n2957), 
	.A2(n2958), 
	.A1(FE_OFN67_n3119));
   XNOR2_X1 U2202 (.ZN(n2927), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U2203 (.ZN(n2928), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U2204 (.ZN(n2929), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2205 (.ZN(n2930), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[28]));
   XNOR2_X1 U2206 (.ZN(n2931), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[27]));
   XNOR2_X1 U2207 (.ZN(n2932), 
	.B(a[7]), 
	.A(b[26]));
   XNOR2_X1 U2208 (.ZN(n2933), 
	.B(a[7]), 
	.A(b[25]));
   XNOR2_X1 U2209 (.ZN(n2934), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[24]));
   XNOR2_X1 U2210 (.ZN(n2935), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[23]));
   XNOR2_X1 U2211 (.ZN(n2936), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[22]));
   XNOR2_X1 U2212 (.ZN(n2937), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[21]));
   XNOR2_X1 U2213 (.ZN(n2938), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[20]));
   XNOR2_X1 U2214 (.ZN(n2939), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[19]));
   XNOR2_X1 U2215 (.ZN(n2940), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[18]));
   XNOR2_X1 U2216 (.ZN(n2941), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[17]));
   XNOR2_X1 U2217 (.ZN(n2942), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[16]));
   XNOR2_X1 U2218 (.ZN(n2943), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[15]));
   XNOR2_X1 U2219 (.ZN(n2944), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[14]));
   XNOR2_X1 U2220 (.ZN(n2945), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[13]));
   XNOR2_X1 U2221 (.ZN(n2946), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[12]));
   XNOR2_X1 U2222 (.ZN(n2947), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[11]));
   XNOR2_X1 U2223 (.ZN(n2948), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[10]));
   XNOR2_X1 U2224 (.ZN(n2949), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U2225 (.ZN(n2950), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[8]));
   XNOR2_X1 U2226 (.ZN(n2951), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[7]));
   XNOR2_X1 U2227 (.ZN(n2952), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[6]));
   XNOR2_X1 U2228 (.ZN(n2953), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[5]));
   XNOR2_X1 U2229 (.ZN(n2954), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(b[4]));
   XNOR2_X1 U2230 (.ZN(n2955), 
	.B(a[7]), 
	.A(b[3]));
   XNOR2_X1 U2231 (.ZN(n2956), 
	.B(a[7]), 
	.A(b[2]));
   XNOR2_X1 U2232 (.ZN(n2957), 
	.B(a[7]), 
	.A(b[1]));
   XNOR2_X1 U2233 (.ZN(n2958), 
	.B(a[7]), 
	.A(b[0]));
   OAI22_X1 U2234 (.ZN(n2016), 
	.B2(FE_OFN75_n3136), 
	.B1(n2992), 
	.A2(FE_PT1_n705), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2236 (.ZN(n2436), 
	.B2(FE_OFN75_n3136), 
	.B1(n2961), 
	.A2(n2962), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2237 (.ZN(n2437), 
	.B2(FE_OFN75_n3136), 
	.B1(n2962), 
	.A2(n2963), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2238 (.ZN(n2438), 
	.B2(FE_OFN75_n3136), 
	.B1(n2963), 
	.A2(n2964), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2239 (.ZN(n2439), 
	.B2(FE_OFN75_n3136), 
	.B1(n2964), 
	.A2(n2965), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2240 (.ZN(n2440), 
	.B2(FE_OFN75_n3136), 
	.B1(n2965), 
	.A2(n2966), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2241 (.ZN(n2441), 
	.B2(FE_OFN75_n3136), 
	.B1(n2966), 
	.A2(n2967), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2242 (.ZN(n2442), 
	.B2(FE_OFN75_n3136), 
	.B1(n2967), 
	.A2(n2968), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2243 (.ZN(n2443), 
	.B2(FE_OFN75_n3136), 
	.B1(n2968), 
	.A2(n2969), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2244 (.ZN(n2444), 
	.B2(FE_OFN75_n3136), 
	.B1(n2969), 
	.A2(n2970), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2245 (.ZN(n2445), 
	.B2(FE_OFN75_n3136), 
	.B1(n2970), 
	.A2(n2971), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2246 (.ZN(n2446), 
	.B2(FE_OFN75_n3136), 
	.B1(n2971), 
	.A2(n2972), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2247 (.ZN(n2447), 
	.B2(FE_OFN75_n3136), 
	.B1(n2972), 
	.A2(n2973), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2248 (.ZN(n2448), 
	.B2(FE_OFN75_n3136), 
	.B1(n2973), 
	.A2(n2974), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2249 (.ZN(n2449), 
	.B2(FE_OFN75_n3136), 
	.B1(n2974), 
	.A2(n2975), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2250 (.ZN(n2450), 
	.B2(FE_OFN75_n3136), 
	.B1(n2975), 
	.A2(n2976), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2251 (.ZN(n2451), 
	.B2(FE_OFN75_n3136), 
	.B1(n2976), 
	.A2(n2977), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2252 (.ZN(n2452), 
	.B2(FE_OFN75_n3136), 
	.B1(n2977), 
	.A2(n2978), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2253 (.ZN(n2453), 
	.B2(FE_OFN75_n3136), 
	.B1(n2978), 
	.A2(n2979), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2254 (.ZN(n2454), 
	.B2(FE_OFN75_n3136), 
	.B1(n2979), 
	.A2(n2980), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2255 (.ZN(n2455), 
	.B2(FE_OFN75_n3136), 
	.B1(n2980), 
	.A2(n2981), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2256 (.ZN(n2456), 
	.B2(FE_OFN75_n3136), 
	.B1(n2981), 
	.A2(n2982), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2257 (.ZN(n2457), 
	.B2(FE_OFN75_n3136), 
	.B1(n2982), 
	.A2(n2983), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2258 (.ZN(n2458), 
	.B2(FE_OFN75_n3136), 
	.B1(n2983), 
	.A2(n2984), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2259 (.ZN(n2459), 
	.B2(FE_OFN75_n3136), 
	.B1(n2984), 
	.A2(n2985), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2260 (.ZN(n2460), 
	.B2(FE_OFN75_n3136), 
	.B1(n2985), 
	.A2(n2986), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2261 (.ZN(n2461), 
	.B2(FE_OFN75_n3136), 
	.B1(n2986), 
	.A2(n2987), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2262 (.ZN(n2462), 
	.B2(FE_OFN75_n3136), 
	.B1(n2987), 
	.A2(n2988), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2263 (.ZN(n2463), 
	.B2(FE_OFN75_n3136), 
	.B1(n2988), 
	.A2(n2989), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2264 (.ZN(n2464), 
	.B2(FE_OFN75_n3136), 
	.B1(n2989), 
	.A2(n2990), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2265 (.ZN(n2465), 
	.B2(FE_OFN75_n3136), 
	.B1(n2990), 
	.A2(n2991), 
	.A1(FE_OFN72_n3120));
   XNOR2_X1 U2266 (.ZN(n2960), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(FE_OFN107_UUT_Mpath_the_mult_x_operand2_31_));
   XNOR2_X1 U2267 (.ZN(n2961), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(FE_OFN111_UUT_Mpath_the_mult_x_operand2_30_));
   XNOR2_X1 U2268 (.ZN(n2962), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2269 (.ZN(n2963), 
	.B(a[5]), 
	.A(b[28]));
   XNOR2_X1 U2270 (.ZN(n2964), 
	.B(a[5]), 
	.A(b[27]));
   XNOR2_X1 U2271 (.ZN(n2965), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[26]));
   XNOR2_X1 U2272 (.ZN(n2966), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[25]));
   XNOR2_X1 U2273 (.ZN(n2967), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[24]));
   XNOR2_X1 U2274 (.ZN(n2968), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[23]));
   XNOR2_X1 U2275 (.ZN(n2969), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[22]));
   XNOR2_X1 U2276 (.ZN(n2970), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[21]));
   XNOR2_X1 U2277 (.ZN(n2971), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[20]));
   XNOR2_X1 U2278 (.ZN(n2972), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[19]));
   XNOR2_X1 U2279 (.ZN(n2973), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[18]));
   XNOR2_X1 U2280 (.ZN(n2974), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[17]));
   XNOR2_X1 U2281 (.ZN(n2975), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[16]));
   XNOR2_X1 U2282 (.ZN(n2976), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[15]));
   XNOR2_X1 U2283 (.ZN(n2977), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[14]));
   XNOR2_X1 U2284 (.ZN(n2978), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[13]));
   XNOR2_X1 U2285 (.ZN(n2979), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[12]));
   XNOR2_X1 U2286 (.ZN(n2980), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[11]));
   XNOR2_X1 U2287 (.ZN(n2981), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[10]));
   XNOR2_X1 U2288 (.ZN(n2982), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(FE_OFN148_UUT_Mpath_the_mult_x_operand2_9_));
   XNOR2_X1 U2289 (.ZN(n2983), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[8]));
   XNOR2_X1 U2290 (.ZN(n2984), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[7]));
   XNOR2_X1 U2291 (.ZN(n2985), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[6]));
   XNOR2_X1 U2292 (.ZN(n2986), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(b[5]));
   XNOR2_X1 U2293 (.ZN(n2987), 
	.B(a[5]), 
	.A(b[4]));
   XNOR2_X1 U2294 (.ZN(n2988), 
	.B(a[5]), 
	.A(b[3]));
   XNOR2_X1 U2295 (.ZN(n2989), 
	.B(a[5]), 
	.A(b[2]));
   XNOR2_X1 U2296 (.ZN(n2990), 
	.B(a[5]), 
	.A(b[1]));
   XNOR2_X1 U2297 (.ZN(n2991), 
	.B(a[5]), 
	.A(b[0]));
   OAI22_X1 U2298 (.ZN(n2017), 
	.B2(FE_OFN81_n3137), 
	.B1(n3025), 
	.A2(n3153), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2300 (.ZN(n2468), 
	.B2(FE_OFN81_n3137), 
	.B1(n2994), 
	.A2(n2995), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2301 (.ZN(n2469), 
	.B2(FE_OFN81_n3137), 
	.B1(n2995), 
	.A2(n2996), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2302 (.ZN(n2470), 
	.B2(FE_OFN81_n3137), 
	.B1(n2996), 
	.A2(n2997), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2303 (.ZN(n2471), 
	.B2(FE_OFN81_n3137), 
	.B1(n2997), 
	.A2(n2998), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2304 (.ZN(n2472), 
	.B2(FE_OFN81_n3137), 
	.B1(n2998), 
	.A2(n2999), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2305 (.ZN(n2473), 
	.B2(FE_OFN81_n3137), 
	.B1(n2999), 
	.A2(n3000), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2306 (.ZN(n2474), 
	.B2(FE_OFN81_n3137), 
	.B1(n3000), 
	.A2(n3001), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2307 (.ZN(n2475), 
	.B2(FE_OFN81_n3137), 
	.B1(n3001), 
	.A2(n3002), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2308 (.ZN(n2476), 
	.B2(FE_OFN81_n3137), 
	.B1(n3002), 
	.A2(n3003), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2309 (.ZN(n2477), 
	.B2(FE_OFN81_n3137), 
	.B1(n3003), 
	.A2(n3004), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2310 (.ZN(n2478), 
	.B2(FE_OFN81_n3137), 
	.B1(n3004), 
	.A2(n3005), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2311 (.ZN(n2479), 
	.B2(FE_OFN81_n3137), 
	.B1(n3005), 
	.A2(n3006), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2312 (.ZN(n2480), 
	.B2(FE_OFN81_n3137), 
	.B1(n3006), 
	.A2(n3007), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2313 (.ZN(n2481), 
	.B2(FE_OFN81_n3137), 
	.B1(n3007), 
	.A2(n3008), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2314 (.ZN(n2482), 
	.B2(FE_OFN81_n3137), 
	.B1(n3008), 
	.A2(n3009), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2315 (.ZN(n2483), 
	.B2(FE_OFN81_n3137), 
	.B1(n3009), 
	.A2(n3010), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2316 (.ZN(n2484), 
	.B2(FE_OFN81_n3137), 
	.B1(n3010), 
	.A2(n3011), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2317 (.ZN(n2485), 
	.B2(FE_OFN81_n3137), 
	.B1(n3011), 
	.A2(n3012), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2318 (.ZN(n2486), 
	.B2(FE_OFN81_n3137), 
	.B1(n3012), 
	.A2(n3013), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2319 (.ZN(n2487), 
	.B2(FE_OFN81_n3137), 
	.B1(n3013), 
	.A2(n3014), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2320 (.ZN(n2488), 
	.B2(FE_OFN81_n3137), 
	.B1(n3014), 
	.A2(n3015), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2321 (.ZN(n2489), 
	.B2(FE_OFN81_n3137), 
	.B1(n3015), 
	.A2(n3016), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2322 (.ZN(n2490), 
	.B2(FE_OFN81_n3137), 
	.B1(n3016), 
	.A2(n3017), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2323 (.ZN(n2491), 
	.B2(FE_OFN81_n3137), 
	.B1(n3017), 
	.A2(n3018), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2324 (.ZN(n2492), 
	.B2(FE_OFN81_n3137), 
	.B1(n3018), 
	.A2(n3019), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2325 (.ZN(n2493), 
	.B2(FE_OFN81_n3137), 
	.B1(n3019), 
	.A2(n3020), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2326 (.ZN(n2494), 
	.B2(FE_OFN81_n3137), 
	.B1(n3020), 
	.A2(n3021), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2327 (.ZN(n2495), 
	.B2(FE_OFN81_n3137), 
	.B1(n3021), 
	.A2(n3022), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2328 (.ZN(n2496), 
	.B2(FE_OFN81_n3137), 
	.B1(n3022), 
	.A2(n3023), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2329 (.ZN(n2497), 
	.B2(FE_OFN81_n3137), 
	.B1(n3023), 
	.A2(n3024), 
	.A1(FE_OFN78_n3121));
   XNOR2_X1 U2330 (.ZN(n2993), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[31]));
   XNOR2_X1 U2331 (.ZN(n2994), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[30]));
   XNOR2_X1 U2332 (.ZN(n2995), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[29]));
   XNOR2_X1 U2333 (.ZN(n2996), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[28]));
   XNOR2_X1 U2334 (.ZN(n2997), 
	.B(a[3]), 
	.A(b[27]));
   XNOR2_X1 U2335 (.ZN(n2998), 
	.B(a[3]), 
	.A(b[26]));
   XNOR2_X1 U2336 (.ZN(n2999), 
	.B(a[3]), 
	.A(b[25]));
   XNOR2_X1 U2337 (.ZN(n3000), 
	.B(a[3]), 
	.A(b[24]));
   XNOR2_X1 U2338 (.ZN(n3001), 
	.B(a[3]), 
	.A(b[23]));
   XNOR2_X1 U2339 (.ZN(n3002), 
	.B(a[3]), 
	.A(b[22]));
   XNOR2_X1 U2340 (.ZN(n3003), 
	.B(a[3]), 
	.A(b[21]));
   XNOR2_X1 U2341 (.ZN(n3004), 
	.B(a[3]), 
	.A(b[20]));
   XNOR2_X1 U2342 (.ZN(n3005), 
	.B(a[3]), 
	.A(b[19]));
   XNOR2_X1 U2343 (.ZN(n3006), 
	.B(a[3]), 
	.A(b[18]));
   XNOR2_X1 U2344 (.ZN(n3007), 
	.B(a[3]), 
	.A(b[17]));
   XNOR2_X1 U2345 (.ZN(n3008), 
	.B(a[3]), 
	.A(b[16]));
   XNOR2_X1 U2346 (.ZN(n3009), 
	.B(a[3]), 
	.A(b[15]));
   XNOR2_X1 U2347 (.ZN(n3010), 
	.B(a[3]), 
	.A(b[14]));
   XNOR2_X1 U2348 (.ZN(n3011), 
	.B(a[3]), 
	.A(b[13]));
   XNOR2_X1 U2349 (.ZN(n3012), 
	.B(a[3]), 
	.A(b[12]));
   XNOR2_X1 U2350 (.ZN(n3013), 
	.B(a[3]), 
	.A(b[11]));
   XNOR2_X1 U2351 (.ZN(n3014), 
	.B(a[3]), 
	.A(b[10]));
   XNOR2_X1 U2352 (.ZN(n3015), 
	.B(a[3]), 
	.A(b[9]));
   XNOR2_X1 U2353 (.ZN(n3016), 
	.B(a[3]), 
	.A(b[8]));
   XNOR2_X1 U2354 (.ZN(n3017), 
	.B(a[3]), 
	.A(b[7]));
   XNOR2_X1 U2355 (.ZN(n3018), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[6]));
   XNOR2_X1 U2356 (.ZN(n3019), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[5]));
   XNOR2_X1 U2357 (.ZN(n3020), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[4]));
   XNOR2_X1 U2358 (.ZN(n3021), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[3]));
   XNOR2_X1 U2359 (.ZN(n3022), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[2]));
   XNOR2_X1 U2360 (.ZN(n3023), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[1]));
   XNOR2_X1 U2361 (.ZN(n3024), 
	.B(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(b[0]));
   OAI22_X1 U2362 (.ZN(n2018), 
	.B2(n3138), 
	.B1(n3058), 
	.A2(FE_PT1_n796), 
	.A1(n3122));
   OAI22_X1 U2363 (.ZN(n2500), 
	.B2(n3138), 
	.B1(n3026), 
	.A2(n3027), 
	.A1(n3122));
   OAI22_X1 U2364 (.ZN(n2501), 
	.B2(n3138), 
	.B1(n3027), 
	.A2(n3028), 
	.A1(n3122));
   OAI22_X1 U2365 (.ZN(n2502), 
	.B2(n3138), 
	.B1(n3028), 
	.A2(n3029), 
	.A1(n3122));
   OAI22_X1 U2366 (.ZN(n2503), 
	.B2(n3138), 
	.B1(n3029), 
	.A2(n3030), 
	.A1(n3122));
   OAI22_X1 U2367 (.ZN(n2504), 
	.B2(n3138), 
	.B1(n3030), 
	.A2(n3031), 
	.A1(n3122));
   OAI22_X1 U2368 (.ZN(n2505), 
	.B2(n3138), 
	.B1(n3031), 
	.A2(n3032), 
	.A1(n3122));
   OAI22_X1 U2369 (.ZN(n2506), 
	.B2(n3138), 
	.B1(n3032), 
	.A2(n3033), 
	.A1(n3122));
   OAI22_X1 U2370 (.ZN(n2507), 
	.B2(n3138), 
	.B1(n3033), 
	.A2(n3034), 
	.A1(n3122));
   OAI22_X1 U2371 (.ZN(n2508), 
	.B2(n3138), 
	.B1(n3034), 
	.A2(n3035), 
	.A1(n3122));
   OAI22_X1 U2372 (.ZN(n2509), 
	.B2(n3138), 
	.B1(n3035), 
	.A2(n3036), 
	.A1(n3122));
   OAI22_X1 U2373 (.ZN(n2510), 
	.B2(n3138), 
	.B1(n3036), 
	.A2(n3037), 
	.A1(n3122));
   OAI22_X1 U2374 (.ZN(n2511), 
	.B2(n3138), 
	.B1(n3037), 
	.A2(n3038), 
	.A1(n3122));
   OAI22_X1 U2375 (.ZN(n2512), 
	.B2(n3138), 
	.B1(n3038), 
	.A2(n3039), 
	.A1(n3122));
   OAI22_X1 U2376 (.ZN(n2513), 
	.B2(n3138), 
	.B1(n3039), 
	.A2(n3040), 
	.A1(n3122));
   OAI22_X1 U2377 (.ZN(n2514), 
	.B2(n3138), 
	.B1(n3040), 
	.A2(n3041), 
	.A1(n3122));
   OAI22_X1 U2378 (.ZN(n2515), 
	.B2(n3138), 
	.B1(n3041), 
	.A2(n3042), 
	.A1(n3122));
   OAI22_X1 U2379 (.ZN(n2516), 
	.B2(n3138), 
	.B1(n3042), 
	.A2(n3043), 
	.A1(n3122));
   OAI22_X1 U2380 (.ZN(n2517), 
	.B2(n3138), 
	.B1(n3043), 
	.A2(n3044), 
	.A1(n3122));
   OAI22_X1 U2381 (.ZN(n2518), 
	.B2(n3138), 
	.B1(n3044), 
	.A2(n3045), 
	.A1(n3122));
   OAI22_X1 U2382 (.ZN(n2519), 
	.B2(n3138), 
	.B1(n3045), 
	.A2(n3046), 
	.A1(n3122));
   OAI22_X1 U2383 (.ZN(n2520), 
	.B2(n3138), 
	.B1(n3046), 
	.A2(n3047), 
	.A1(n3122));
   OAI22_X1 U2384 (.ZN(n2521), 
	.B2(n3138), 
	.B1(n3047), 
	.A2(n3048), 
	.A1(n3122));
   OAI22_X1 U2385 (.ZN(n2522), 
	.B2(n3138), 
	.B1(n3048), 
	.A2(n3049), 
	.A1(n3122));
   OAI22_X1 U2386 (.ZN(n2523), 
	.B2(n3138), 
	.B1(n3049), 
	.A2(n3050), 
	.A1(n3122));
   OAI22_X1 U2387 (.ZN(n2524), 
	.B2(n3138), 
	.B1(n3050), 
	.A2(n3051), 
	.A1(n3122));
   OAI22_X1 U2388 (.ZN(n2525), 
	.B2(n3138), 
	.B1(n3051), 
	.A2(n3052), 
	.A1(n3122));
   OAI22_X1 U2389 (.ZN(n2526), 
	.B2(n3138), 
	.B1(n3052), 
	.A2(n3053), 
	.A1(n3122));
   OAI22_X1 U2390 (.ZN(n2527), 
	.B2(n3138), 
	.B1(n3053), 
	.A2(n3054), 
	.A1(n3122));
   OAI22_X1 U2391 (.ZN(n2528), 
	.B2(n3138), 
	.B1(n3054), 
	.A2(n3055), 
	.A1(n3122));
   OAI22_X1 U2392 (.ZN(n2529), 
	.B2(n3138), 
	.B1(n3055), 
	.A2(n3056), 
	.A1(n3122));
   OAI22_X1 U2393 (.ZN(n2530), 
	.B2(n3138), 
	.B1(n3056), 
	.A2(n3057), 
	.A1(n3122));
   XNOR2_X1 U2394 (.ZN(n3026), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[31]));
   XNOR2_X1 U2395 (.ZN(n3027), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[30]));
   XNOR2_X1 U2396 (.ZN(n3028), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(FE_OFN112_UUT_Mpath_the_mult_x_operand2_29_));
   XNOR2_X1 U2397 (.ZN(n3029), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[28]));
   XNOR2_X1 U2398 (.ZN(n3030), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[27]));
   XNOR2_X1 U2399 (.ZN(n3031), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[26]));
   XNOR2_X1 U2400 (.ZN(n3032), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[25]));
   XNOR2_X1 U2401 (.ZN(n3033), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[24]));
   XNOR2_X1 U2402 (.ZN(n3034), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[23]));
   XNOR2_X1 U2403 (.ZN(n3035), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[22]));
   XNOR2_X1 U2404 (.ZN(n3036), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[21]));
   XNOR2_X1 U2405 (.ZN(n3037), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[20]));
   XNOR2_X1 U2406 (.ZN(n3038), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[19]));
   XNOR2_X1 U2407 (.ZN(n3039), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[18]));
   XNOR2_X1 U2408 (.ZN(n3040), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[17]));
   XNOR2_X1 U2409 (.ZN(n3041), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[16]));
   XNOR2_X1 U2410 (.ZN(n3042), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[15]));
   XNOR2_X1 U2411 (.ZN(n3043), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[14]));
   XNOR2_X1 U2412 (.ZN(n3044), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[13]));
   XNOR2_X1 U2413 (.ZN(n3045), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[12]));
   XNOR2_X1 U2414 (.ZN(n3046), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[11]));
   XNOR2_X1 U2415 (.ZN(n3047), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[10]));
   XNOR2_X1 U2416 (.ZN(n3048), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[9]));
   XNOR2_X1 U2417 (.ZN(n3049), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[8]));
   XNOR2_X1 U2418 (.ZN(n3050), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[7]));
   XNOR2_X1 U2419 (.ZN(n3051), 
	.B(FE_OFN172_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(b[6]));
   XNOR2_X1 U2420 (.ZN(n3052), 
	.B(a[1]), 
	.A(b[5]));
   XNOR2_X1 U2421 (.ZN(n3053), 
	.B(a[1]), 
	.A(b[4]));
   XNOR2_X1 U2422 (.ZN(n3054), 
	.B(a[1]), 
	.A(b[3]));
   XNOR2_X1 U2423 (.ZN(n3055), 
	.B(a[1]), 
	.A(b[2]));
   XNOR2_X1 U2424 (.ZN(n3056), 
	.B(a[1]), 
	.A(b[1]));
   XNOR2_X1 U2425 (.ZN(n3057), 
	.B(a[1]), 
	.A(b[0]));
   INV_X1 U2458 (.ZN(n3140), 
	.A(FE_OFN114_UUT_Mpath_the_mult_x_operand1_29_));
   INV_X1 U2460 (.ZN(n3141), 
	.A(FE_OFN118_UUT_Mpath_the_mult_x_operand1_27_));
   INV_X1 U2462 (.ZN(n3142), 
	.A(FE_OFN122_UUT_Mpath_the_mult_x_operand1_25_));
   INV_X1 U2468 (.ZN(n3145), 
	.A(FE_OFN131_UUT_Mpath_the_mult_x_operand1_19_));
   INV_X1 U2470 (.ZN(n3146), 
	.A(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_));
   INV_X1 U2484 (.ZN(n3153), 
	.A(FE_OFN166_UUT_Mpath_the_mult_x_operand1_3_));
   XOR2_X1 U2489 (.Z(n3091), 
	.B(a[31]), 
	.A(a[30]));
   XOR2_X1 U2492 (.Z(n3092), 
	.B(a[29]), 
	.A(a[28]));
   XOR2_X1 U2495 (.Z(n3093), 
	.B(a[27]), 
	.A(a[26]));
   XOR2_X1 U2498 (.Z(n3094), 
	.B(a[25]), 
	.A(a[24]));
   XOR2_X1 U2501 (.Z(n3095), 
	.B(a[23]), 
	.A(a[22]));
   XOR2_X1 U2504 (.Z(n3096), 
	.B(a[21]), 
	.A(a[20]));
   XOR2_X1 U2507 (.Z(n3097), 
	.B(a[19]), 
	.A(a[18]));
   XOR2_X1 U2510 (.Z(n3098), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(a[16]));
   XOR2_X1 U2513 (.Z(n3099), 
	.B(a[15]), 
	.A(a[14]));
   XOR2_X1 U2516 (.Z(n3100), 
	.B(a[13]), 
	.A(a[12]));
   XOR2_X1 U2519 (.Z(n3101), 
	.B(a[11]), 
	.A(a[10]));
   XOR2_X1 U2522 (.Z(n3102), 
	.B(a[9]), 
	.A(a[8]));
   XOR2_X1 U2525 (.Z(n3103), 
	.B(a[7]), 
	.A(a[6]));
   XOR2_X1 U2528 (.Z(n3104), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(a[4]));
   XOR2_X1 U2531 (.Z(n3105), 
	.B(a[3]), 
	.A(a[2]));
   NAND2_X2 U2533 (.ZN(n3122), 
	.A2(n3138), 
	.A1(n3106));
   XOR2_X1 U2534 (.Z(n3106), 
	.B(a[1]), 
	.A(a[0]));
   INV_X2 U2535 (.ZN(n3138), 
	.A(a[0]));
   OAI22_X1 U2538 (.ZN(n1103), 
	.B2(FE_OFN40_n3126), 
	.B1(n2630), 
	.A2(n2631), 
	.A1(FE_OFN39_n3110));
   OAI22_X1 U2540 (.ZN(n1233), 
	.B2(FE_OFN52_n3131), 
	.B1(n2795), 
	.A2(n2796), 
	.A1(FE_OFN51_n3115));
   OAI22_X1 U2542 (.ZN(n1271), 
	.B2(FE_OFN58_n3132), 
	.B1(n2828), 
	.A2(n2829), 
	.A1(FE_OFN55_n3116));
   OAI22_X1 U2544 (.ZN(n1409), 
	.B2(FE_OFN70_n3135), 
	.B1(n2927), 
	.A2(n2928), 
	.A1(FE_OFN67_n3119));
   OAI22_X1 U2546 (.ZN(n1313), 
	.B2(FE_OFN64_n3133), 
	.B1(n2861), 
	.A2(n2862), 
	.A1(FE_OFN61_n3117));
   OAI22_X1 U2548 (.ZN(n1079), 
	.B2(FE_OFN36_n3124), 
	.B1(n2564), 
	.A2(n2565), 
	.A1(FE_OFN33_n3108));
   OAI22_X1 U2550 (.ZN(n1089), 
	.B2(FE_OFN38_n3125), 
	.B1(n2597), 
	.A2(n2598), 
	.A1(FE_OFN37_n3109));
   OAI22_X1 U2552 (.ZN(n1121), 
	.B2(FE_OFN42_n3127), 
	.B1(n2663), 
	.A2(n2664), 
	.A1(FE_OFN41_n3111));
   OAI22_X1 U2554 (.ZN(n1463), 
	.B2(FE_OFN75_n3136), 
	.B1(n2960), 
	.A2(n2961), 
	.A1(FE_OFN72_n3120));
   OAI22_X1 U2556 (.ZN(n1169), 
	.B2(FE_OFN46_n3129), 
	.B1(n2729), 
	.A2(n2730), 
	.A1(FE_OFN45_n3113));
   OAI22_X1 U2558 (.ZN(n1199), 
	.B2(FE_OFN48_n3130), 
	.B1(n2762), 
	.A2(n2763), 
	.A1(FE_OFN47_n3114));
   OAI22_X1 U2560 (.ZN(n1521), 
	.B2(FE_OFN81_n3137), 
	.B1(n2993), 
	.A2(n2994), 
	.A1(FE_OFN78_n3121));
   OAI22_X1 U2562 (.ZN(n1143), 
	.B2(FE_OFN44_n3128), 
	.B1(n2696), 
	.A2(n2697), 
	.A1(FE_OFN43_n3112));
   OAI22_X1 U2564 (.ZN(n1359), 
	.B2(FE_OFN66_n3134), 
	.B1(n2894), 
	.A2(n2895), 
	.A1(FE_OFN65_n3118));
   OAI22_X1 U2566 (.ZN(n1073), 
	.B2(FE_OFN35_n3123), 
	.B1(n2531), 
	.A2(n2532), 
	.A1(FE_OFN34_n3107));
   NAND2_X1 U2571 (.ZN(n3113), 
	.A2(FE_OFN46_n3129), 
	.A1(n3097));
   XNOR2_X1 U2572 (.ZN(n3129), 
	.B(FE_OFN135_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(a[18]));
   NAND2_X1 U2576 (.ZN(n3117), 
	.A2(n3133), 
	.A1(n3101));
   XNOR2_X1 U2577 (.ZN(n3133), 
	.B(a[9]), 
	.A(a[10]));
   NAND2_X1 U2581 (.ZN(n3112), 
	.A2(FE_OFN44_n3128), 
	.A1(n3096));
   XNOR2_X1 U2582 (.ZN(n3128), 
	.B(a[19]), 
	.A(a[20]));
   NAND2_X1 U2586 (.ZN(n3116), 
	.A2(n3132), 
	.A1(n3100));
   XNOR2_X1 U2587 (.ZN(n3132), 
	.B(a[11]), 
	.A(a[12]));
   NAND2_X1 U2591 (.ZN(n3115), 
	.A2(n3131), 
	.A1(n3099));
   XNOR2_X1 U2592 (.ZN(n3131), 
	.B(a[13]), 
	.A(a[14]));
   NAND2_X1 U2596 (.ZN(n3114), 
	.A2(FE_OFN48_n3130), 
	.A1(n3098));
   XNOR2_X1 U2597 (.ZN(n3130), 
	.B(a[15]), 
	.A(a[16]));
   NAND2_X1 U2601 (.ZN(n3111), 
	.A2(FE_OFN42_n3127), 
	.A1(n3095));
   XNOR2_X1 U2602 (.ZN(n3127), 
	.B(a[21]), 
	.A(a[22]));
   NAND2_X1 U2606 (.ZN(n3109), 
	.A2(n3125), 
	.A1(n3093));
   XNOR2_X1 U2607 (.ZN(n3125), 
	.B(a[25]), 
	.A(a[26]));
   NAND2_X1 U2611 (.ZN(n3110), 
	.A2(n3126), 
	.A1(n3094));
   XNOR2_X1 U2612 (.ZN(n3126), 
	.B(a[23]), 
	.A(a[24]));
   NAND2_X1 U2616 (.ZN(n3108), 
	.A2(n3124), 
	.A1(n3092));
   XNOR2_X1 U2617 (.ZN(n3124), 
	.B(a[27]), 
	.A(a[28]));
   NAND2_X1 U2621 (.ZN(n3121), 
	.A2(FE_OFN81_n3137), 
	.A1(n3105));
   XNOR2_X1 U2622 (.ZN(n3137), 
	.B(a[1]), 
	.A(a[2]));
   NAND2_X1 U2626 (.ZN(n3120), 
	.A2(FE_OFN75_n3136), 
	.A1(n3104));
   XNOR2_X1 U2627 (.ZN(n3136), 
	.B(a[3]), 
	.A(a[4]));
   NAND2_X1 U2631 (.ZN(n3119), 
	.A2(FE_OFN70_n3135), 
	.A1(n3103));
   XNOR2_X1 U2632 (.ZN(n3135), 
	.B(FE_OFN157_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(a[6]));
   NAND2_X1 U2636 (.ZN(n3118), 
	.A2(n3134), 
	.A1(n3102));
   XNOR2_X1 U2637 (.ZN(n3134), 
	.B(FE_OFN153_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(a[8]));
   NAND2_X1 U2641 (.ZN(n3107), 
	.A2(n3123), 
	.A1(n3091));
   XNOR2_X1 U2642 (.ZN(n3123), 
	.B(a[29]), 
	.A(a[30]));
endmodule

module up_island_DW01_add_3 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	FE_PT1__UUT_Mpath_the_alu_N182_, 
	FE_PT1__UUT_Mpath_the_alu_N183_, 
	FE_PT1__UUT_Mpath_the_alu_N169_, 
	FE_PT1__UUT_Mpath_the_alu_N170_, 
	FE_PT1__UUT_Mpath_the_alu_N164_, 
	FE_PT1__UUT_Mpath_the_alu_N165_, 
	FE_PT1__UUT_Mpath_the_alu_N162_, 
	FE_PT1__UUT_Mpath_the_alu_N171_, 
	FE_PT1__UUT_Mpath_the_alu_N184_, 
	FE_PT1__UUT_Mpath_the_alu_N163_, 
	FE_PT1__UUT_Mpath_the_alu_N172_, 
	FE_PT1__UUT_Mpath_the_alu_N166_, 
	FE_PT1__UUT_Mpath_the_alu_N173_, 
	FE_PT1__UUT_Mpath_the_alu_N167_, 
	FE_PT1__UUT_Mpath_the_alu_N174_, 
	FE_PT1__UUT_Mpath_the_alu_N168_, 
	FE_PT1__UUT_Mpath_the_alu_N175_, 
	FE_PT1__UUT_Mpath_the_alu_N159_, 
	FE_PT1__UUT_Mpath_the_alu_N176_, 
	FE_PT1__UUT_Mpath_the_alu_N177_, 
	FE_PT1__UUT_Mpath_the_alu_N178_, 
	FE_OFN181_UUT_Mpath_out_regB_0_);
   input [31:0] A;
   input [31:0] B;
   input CI;
   output [31:0] SUM;
   output CO;
   input FE_PT1__UUT_Mpath_the_alu_N182_;
   input FE_PT1__UUT_Mpath_the_alu_N183_;
   input FE_PT1__UUT_Mpath_the_alu_N169_;
   input FE_PT1__UUT_Mpath_the_alu_N170_;
   input FE_PT1__UUT_Mpath_the_alu_N164_;
   input FE_PT1__UUT_Mpath_the_alu_N165_;
   input FE_PT1__UUT_Mpath_the_alu_N162_;
   input FE_PT1__UUT_Mpath_the_alu_N171_;
   input FE_PT1__UUT_Mpath_the_alu_N184_;
   input FE_PT1__UUT_Mpath_the_alu_N163_;
   input FE_PT1__UUT_Mpath_the_alu_N172_;
   input FE_PT1__UUT_Mpath_the_alu_N166_;
   input FE_PT1__UUT_Mpath_the_alu_N173_;
   input FE_PT1__UUT_Mpath_the_alu_N167_;
   input FE_PT1__UUT_Mpath_the_alu_N174_;
   input FE_PT1__UUT_Mpath_the_alu_N168_;
   input FE_PT1__UUT_Mpath_the_alu_N175_;
   input FE_PT1__UUT_Mpath_the_alu_N159_;
   input FE_PT1__UUT_Mpath_the_alu_N176_;
   input FE_PT1__UUT_Mpath_the_alu_N177_;
   input FE_PT1__UUT_Mpath_the_alu_N178_;
   input FE_OFN181_UUT_Mpath_out_regB_0_;

   // Internal wires
   wire \carry[31] ;
   wire \carry[29] ;
   wire \carry[28] ;
   wire \carry[26] ;
   wire \carry[21] ;
   wire \carry[16] ;
   wire \carry[15] ;
   wire \carry[14] ;
   wire \carry[13] ;
   wire \carry[12] ;
   wire \carry[11] ;
   wire \carry[10] ;
   wire \carry[9] ;
   wire \carry[8] ;
   wire \carry[7] ;
   wire \carry[1] ;
   wire n3;
   wire n5;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n18;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n37;
   wire n38;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n54;
   wire n55;
   wire n56;
   wire n58;
   wire n60;
   wire n62;
   wire n63;
   wire n64;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n73;
   wire n74;
   wire n75;
   wire n77;
   wire n79;
   wire n80;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n91;
   wire n92;
   wire n93;
   wire n95;
   wire n96;
   wire n98;
   wire n99;
   wire n101;
   wire n102;
   wire n103;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n115;
   wire n116;
   wire n117;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n124;
   wire n125;
   wire n126;
   wire n130;
   wire n133;
   wire n134;
   wire n135;
   wire n137;
   wire n138;
   wire n139;
   wire n141;
   wire n142;
   wire n143;
   wire n145;
   wire n146;
   wire n147;
   wire n150;
   wire n151;
   wire n152;
   wire n154;
   wire n155;
   wire n156;
   wire n158;
   wire n159;
   wire n161;
   wire n162;
   wire n163;

   FA_X1 U1_10 (.S(SUM[10]), 
	.CO(\carry[11] ), 
	.CI(\carry[10] ), 
	.B(B[10]), 
	.A(A[10]));
   FA_X1 U1_9 (.S(SUM[9]), 
	.CO(\carry[10] ), 
	.CI(\carry[9] ), 
	.B(B[9]), 
	.A(A[9]));
   FA_X1 U1_8 (.S(SUM[8]), 
	.CO(\carry[9] ), 
	.CI(\carry[8] ), 
	.B(B[8]), 
	.A(A[8]));
   NAND2_X1 U1 (.ZN(n49), 
	.A2(B[12]), 
	.A1(A[12]));
   NAND2_X1 U2 (.ZN(n158), 
	.A2(B[6]), 
	.A1(A[6]));
   INV_X1 U3 (.ZN(n38), 
	.A(n44));
   INV_X1 U4 (.ZN(n50), 
	.A(FE_PT1__UUT_Mpath_the_alu_N163_));
   INV_X1 U5 (.ZN(n99), 
	.A(n108));
   INV_X1 U6 (.ZN(n51), 
	.A(FE_PT1__UUT_Mpath_the_alu_N162_));
   NAND3_X2 U7 (.ZN(\carry[16] ), 
	.A3(n92), 
	.A2(n93), 
	.A1(n91));
   NAND3_X1 U8 (.ZN(\carry[12] ), 
	.A3(n41), 
	.A2(n42), 
	.A1(n40));
   NAND3_X1 U9 (.ZN(\carry[29] ), 
	.A3(n112), 
	.A2(n113), 
	.A1(n111));
   NAND3_X1 U10 (.ZN(\carry[13] ), 
	.A3(n48), 
	.A2(n49), 
	.A1(n47));
   NAND3_X1 U12 (.ZN(\carry[14] ), 
	.A3(n55), 
	.A2(n56), 
	.A1(n54));
   XNOR2_X1 U14 (.ZN(SUM[29]), 
	.B(n3), 
	.A(\carry[29] ));
   XNOR2_X1 U15 (.ZN(n3), 
	.B(B[29]), 
	.A(A[29]));
   NAND3_X1 U17 (.ZN(n5), 
	.A3(n22), 
	.A2(n23), 
	.A1(n21));
   NAND2_X1 U20 (.ZN(n7), 
	.A2(A[6]), 
	.A1(n66));
   NAND3_X1 U21 (.ZN(n8), 
	.A3(n7), 
	.A2(n158), 
	.A1(n159));
   NAND3_X1 U22 (.ZN(\carry[15] ), 
	.A3(n74), 
	.A2(n75), 
	.A1(n73));
   NAND3_X1 U23 (.ZN(\carry[7] ), 
	.A3(n158), 
	.A2(n159), 
	.A1(n7));
   NAND2_X1 U24 (.ZN(n9), 
	.A2(B[5]), 
	.A1(n10));
   NAND3_X1 U25 (.ZN(n10), 
	.A3(n86), 
	.A2(n88), 
	.A1(n87));
   AND3_X1 U26 (.ZN(n11), 
	.A3(n146), 
	.A2(n147), 
	.A1(n145));
   NAND3_X1 U28 (.ZN(n12), 
	.A3(n28), 
	.A2(n29), 
	.A1(n27));
   NAND3_X1 U29 (.ZN(n13), 
	.A3(n142), 
	.A2(n143), 
	.A1(n141));
   NAND2_X1 U30 (.ZN(n14), 
	.A2(A[29]), 
	.A1(\carry[29] ));
   NAND3_X1 U35 (.ZN(n18), 
	.A3(n69), 
	.A2(n70), 
	.A1(n68));
   AND2_X1 U36 (.ZN(\carry[1] ), 
	.A2(FE_OFN181_UUT_Mpath_out_regB_0_), 
	.A1(A[0]));
   XOR2_X1 U38 (.Z(n20), 
	.B(A[1]), 
	.A(B[1]));
   XOR2_X1 U39 (.Z(SUM[1]), 
	.B(n20), 
	.A(\carry[1] ));
   NAND2_X1 U40 (.ZN(n21), 
	.A2(B[1]), 
	.A1(\carry[1] ));
   NAND2_X1 U41 (.ZN(n22), 
	.A2(A[1]), 
	.A1(\carry[1] ));
   NAND2_X1 U42 (.ZN(n23), 
	.A2(A[1]), 
	.A1(B[1]));
   NAND2_X1 U44 (.ZN(n24), 
	.A2(A[5]), 
	.A1(n10));
   XOR2_X1 U46 (.Z(n26), 
	.B(A[2]), 
	.A(B[2]));
   XOR2_X1 U47 (.Z(SUM[2]), 
	.B(n26), 
	.A(n5));
   NAND2_X1 U48 (.ZN(n27), 
	.A2(B[2]), 
	.A1(n5));
   NAND2_X1 U49 (.ZN(n28), 
	.A2(A[2]), 
	.A1(n5));
   NAND2_X1 U50 (.ZN(n29), 
	.A2(A[2]), 
	.A1(B[2]));
   NAND3_X1 U52 (.ZN(n30), 
	.A3(n60), 
	.A2(n58), 
	.A1(n14));
   NAND2_X1 U54 (.ZN(n125), 
	.A2(B[26]), 
	.A1(\carry[26] ));
   INV_X1 U61 (.ZN(n37), 
	.A(n11));
   XNOR2_X1 U62 (.ZN(SUM[28]), 
	.B(n38), 
	.A(n43));
   XOR2_X1 U64 (.Z(SUM[11]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N178_), 
	.A(\carry[11] ));
   NAND2_X1 U65 (.ZN(n40), 
	.A2(A[11]), 
	.A1(\carry[11] ));
   NAND2_X1 U66 (.ZN(n41), 
	.A2(B[11]), 
	.A1(\carry[11] ));
   NAND2_X1 U67 (.ZN(n42), 
	.A2(B[11]), 
	.A1(A[11]));
   AND3_X1 U68 (.ZN(n43), 
	.A3(n138), 
	.A2(n139), 
	.A1(n137));
   XNOR2_X1 U69 (.ZN(n44), 
	.B(B[28]), 
	.A(A[28]));
   NAND2_X1 U70 (.ZN(n45), 
	.A2(A[26]), 
	.A1(n37));
   XOR2_X1 U72 (.Z(SUM[12]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N177_), 
	.A(\carry[12] ));
   NAND2_X1 U73 (.ZN(n47), 
	.A2(A[12]), 
	.A1(\carry[12] ));
   NAND2_X1 U74 (.ZN(n48), 
	.A2(B[12]), 
	.A1(\carry[12] ));
   XNOR2_X1 U75 (.ZN(SUM[26]), 
	.B(n50), 
	.A(n37));
   XNOR2_X1 U76 (.ZN(SUM[27]), 
	.B(n51), 
	.A(n96));
   XOR2_X1 U79 (.Z(SUM[13]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N176_), 
	.A(\carry[13] ));
   NAND2_X1 U80 (.ZN(n54), 
	.A2(A[13]), 
	.A1(\carry[13] ));
   NAND2_X1 U81 (.ZN(n55), 
	.A2(B[13]), 
	.A1(\carry[13] ));
   NAND2_X1 U82 (.ZN(n56), 
	.A2(B[13]), 
	.A1(A[13]));
   NAND2_X1 U84 (.ZN(n58), 
	.A2(B[29]), 
	.A1(A[29]));
   NAND2_X1 U85 (.ZN(n60), 
	.A2(\carry[29] ), 
	.A1(B[29]));
   XOR2_X1 U87 (.Z(SUM[30]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N159_), 
	.A(n30));
   NAND2_X1 U88 (.ZN(n62), 
	.A2(B[30]), 
	.A1(A[30]));
   NAND2_X1 U89 (.ZN(n63), 
	.A2(A[30]), 
	.A1(n30));
   NAND2_X1 U90 (.ZN(n64), 
	.A2(B[30]), 
	.A1(n30));
   NAND3_X1 U91 (.ZN(\carry[31] ), 
	.A3(n62), 
	.A2(n64), 
	.A1(n63));
   NAND3_X1 U93 (.ZN(n66), 
	.A3(n9), 
	.A2(n130), 
	.A1(n24));
   XOR2_X1 U94 (.Z(n67), 
	.B(B[3]), 
	.A(A[3]));
   XOR2_X1 U95 (.Z(SUM[3]), 
	.B(n67), 
	.A(n12));
   NAND2_X1 U96 (.ZN(n68), 
	.A2(A[3]), 
	.A1(n12));
   NAND2_X1 U97 (.ZN(n69), 
	.A2(B[3]), 
	.A1(n12));
   NAND2_X1 U98 (.ZN(n70), 
	.A2(B[3]), 
	.A1(A[3]));
   XOR2_X1 U102 (.Z(SUM[14]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N175_), 
	.A(\carry[14] ));
   NAND2_X1 U103 (.ZN(n73), 
	.A2(A[14]), 
	.A1(\carry[14] ));
   NAND2_X1 U104 (.ZN(n74), 
	.A2(B[14]), 
	.A1(\carry[14] ));
   NAND2_X1 U105 (.ZN(n75), 
	.A2(B[14]), 
	.A1(A[14]));
   NAND3_X1 U107 (.ZN(n77), 
	.A3(n83), 
	.A2(n84), 
	.A1(n82));
   NAND3_X1 U109 (.ZN(n79), 
	.A3(n116), 
	.A2(n117), 
	.A1(n115));
   NAND3_X1 U110 (.ZN(n80), 
	.A3(n120), 
	.A2(n121), 
	.A1(n119));
   XOR2_X1 U112 (.Z(SUM[21]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N168_), 
	.A(\carry[21] ));
   NAND2_X1 U113 (.ZN(n82), 
	.A2(A[21]), 
	.A1(\carry[21] ));
   NAND2_X1 U114 (.ZN(n83), 
	.A2(B[21]), 
	.A1(\carry[21] ));
   NAND2_X1 U115 (.ZN(n84), 
	.A2(B[21]), 
	.A1(A[21]));
   XOR2_X1 U117 (.Z(n85), 
	.B(A[4]), 
	.A(B[4]));
   XOR2_X1 U118 (.Z(SUM[4]), 
	.B(n85), 
	.A(n18));
   NAND2_X1 U119 (.ZN(n86), 
	.A2(B[4]), 
	.A1(n18));
   NAND2_X1 U120 (.ZN(n87), 
	.A2(A[4]), 
	.A1(n18));
   NAND2_X1 U121 (.ZN(n88), 
	.A2(A[4]), 
	.A1(B[4]));
   NAND3_X1 U122 (.ZN(n89), 
	.A3(n106), 
	.A2(n107), 
	.A1(n105));
   XOR2_X1 U124 (.Z(SUM[15]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N174_), 
	.A(\carry[15] ));
   NAND2_X1 U125 (.ZN(n91), 
	.A2(A[15]), 
	.A1(\carry[15] ));
   NAND2_X1 U126 (.ZN(n92), 
	.A2(B[15]), 
	.A1(\carry[15] ));
   NAND2_X1 U127 (.ZN(n93), 
	.A2(B[15]), 
	.A1(A[15]));
   NAND2_X1 U129 (.ZN(n124), 
	.A2(A[26]), 
	.A1(\carry[26] ));
   NAND3_X1 U130 (.ZN(n96), 
	.A3(n125), 
	.A2(n126), 
	.A1(n45));
   NAND3_X1 U131 (.ZN(n95), 
	.A3(n124), 
	.A2(n126), 
	.A1(n125));
   NAND3_X1 U133 (.ZN(n98), 
	.A3(n102), 
	.A2(n103), 
	.A1(n101));
   XNOR2_X1 U134 (.ZN(SUM[31]), 
	.B(n99), 
	.A(\carry[31] ));
   XOR2_X1 U136 (.Z(SUM[22]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N167_), 
	.A(n77));
   NAND2_X1 U137 (.ZN(n101), 
	.A2(A[22]), 
	.A1(n77));
   NAND2_X1 U138 (.ZN(n102), 
	.A2(B[22]), 
	.A1(n77));
   NAND2_X1 U139 (.ZN(n103), 
	.A2(B[22]), 
	.A1(A[22]));
   XOR2_X1 U142 (.Z(SUM[16]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N173_), 
	.A(\carry[16] ));
   NAND2_X1 U143 (.ZN(n105), 
	.A2(A[16]), 
	.A1(\carry[16] ));
   NAND2_X1 U144 (.ZN(n106), 
	.A2(B[16]), 
	.A1(\carry[16] ));
   NAND2_X1 U145 (.ZN(n107), 
	.A2(B[16]), 
	.A1(A[16]));
   XOR2_X1 U147 (.Z(n108), 
	.B(B[31]), 
	.A(A[31]));
   NAND3_X1 U149 (.ZN(n110), 
	.A3(n134), 
	.A2(n135), 
	.A1(n133));
   NAND3_X1 U150 (.ZN(\carry[26] ), 
	.A3(n146), 
	.A2(n147), 
	.A1(n145));
   NAND2_X1 U151 (.ZN(n111), 
	.A2(A[28]), 
	.A1(\carry[28] ));
   NAND2_X1 U152 (.ZN(n112), 
	.A2(B[28]), 
	.A1(\carry[28] ));
   NAND2_X1 U153 (.ZN(n113), 
	.A2(B[28]), 
	.A1(A[28]));
   XOR2_X1 U155 (.Z(SUM[23]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N166_), 
	.A(n98));
   NAND2_X1 U156 (.ZN(n115), 
	.A2(A[23]), 
	.A1(n98));
   NAND2_X1 U157 (.ZN(n116), 
	.A2(B[23]), 
	.A1(n98));
   NAND2_X1 U158 (.ZN(n117), 
	.A2(B[23]), 
	.A1(A[23]));
   XOR2_X1 U160 (.Z(SUM[17]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N172_), 
	.A(n89));
   NAND2_X1 U161 (.ZN(n119), 
	.A2(A[17]), 
	.A1(n89));
   NAND2_X1 U162 (.ZN(n120), 
	.A2(B[17]), 
	.A1(n89));
   NAND2_X1 U163 (.ZN(n121), 
	.A2(B[17]), 
	.A1(A[17]));
   NAND3_X1 U165 (.ZN(n122), 
	.A3(n151), 
	.A2(n152), 
	.A1(n150));
   NAND2_X1 U167 (.ZN(n126), 
	.A2(B[26]), 
	.A1(A[26]));
   XOR2_X1 U169 (.Z(SUM[5]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N184_), 
	.A(n10));
   NAND2_X1 U172 (.ZN(n130), 
	.A2(B[5]), 
	.A1(A[5]));
   XOR2_X1 U175 (.Z(SUM[18]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N171_), 
	.A(n80));
   NAND2_X1 U176 (.ZN(n133), 
	.A2(A[18]), 
	.A1(n80));
   NAND2_X1 U177 (.ZN(n134), 
	.A2(B[18]), 
	.A1(n80));
   NAND2_X1 U178 (.ZN(n135), 
	.A2(B[18]), 
	.A1(A[18]));
   NAND2_X1 U181 (.ZN(n137), 
	.A2(A[27]), 
	.A1(n95));
   NAND2_X1 U182 (.ZN(n138), 
	.A2(B[27]), 
	.A1(n95));
   NAND2_X1 U183 (.ZN(n139), 
	.A2(B[27]), 
	.A1(A[27]));
   NAND3_X1 U184 (.ZN(\carry[28] ), 
	.A3(n139), 
	.A2(n138), 
	.A1(n137));
   XOR2_X1 U186 (.Z(SUM[24]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N165_), 
	.A(n79));
   NAND2_X1 U187 (.ZN(n141), 
	.A2(A[24]), 
	.A1(n79));
   NAND2_X1 U188 (.ZN(n142), 
	.A2(B[24]), 
	.A1(n79));
   NAND2_X1 U189 (.ZN(n143), 
	.A2(B[24]), 
	.A1(A[24]));
   XOR2_X1 U191 (.Z(SUM[25]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N164_), 
	.A(n13));
   NAND2_X1 U192 (.ZN(n145), 
	.A2(A[25]), 
	.A1(n13));
   NAND2_X1 U193 (.ZN(n146), 
	.A2(B[25]), 
	.A1(n13));
   NAND2_X1 U194 (.ZN(n147), 
	.A2(B[25]), 
	.A1(A[25]));
   XOR2_X1 U197 (.Z(SUM[19]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N170_), 
	.A(n110));
   NAND2_X1 U198 (.ZN(n150), 
	.A2(A[19]), 
	.A1(n110));
   NAND2_X1 U199 (.ZN(n151), 
	.A2(B[19]), 
	.A1(n110));
   NAND2_X1 U200 (.ZN(n152), 
	.A2(B[19]), 
	.A1(A[19]));
   XOR2_X1 U203 (.Z(SUM[20]), 
	.B(FE_PT1__UUT_Mpath_the_alu_N169_), 
	.A(n122));
   NAND2_X1 U204 (.ZN(n154), 
	.A2(A[20]), 
	.A1(n122));
   NAND2_X1 U205 (.ZN(n155), 
	.A2(B[20]), 
	.A1(n122));
   NAND2_X1 U206 (.ZN(n156), 
	.A2(B[20]), 
	.A1(A[20]));
   NAND3_X1 U207 (.ZN(\carry[21] ), 
	.A3(n155), 
	.A2(n156), 
	.A1(n154));
   XOR2_X1 U209 (.Z(SUM[6]), 
	.B(n66), 
	.A(FE_PT1__UUT_Mpath_the_alu_N183_));
   NAND2_X1 U210 (.ZN(n159), 
	.A2(n66), 
	.A1(B[6]));
   XOR2_X1 U212 (.Z(SUM[7]), 
	.B(n8), 
	.A(FE_PT1__UUT_Mpath_the_alu_N182_));
   NAND2_X1 U213 (.ZN(n161), 
	.A2(B[7]), 
	.A1(A[7]));
   NAND2_X1 U214 (.ZN(n162), 
	.A2(\carry[7] ), 
	.A1(A[7]));
   NAND2_X1 U215 (.ZN(n163), 
	.A2(B[7]), 
	.A1(n8));
   NAND3_X1 U216 (.ZN(\carry[8] ), 
	.A3(n161), 
	.A2(n163), 
	.A1(n162));
   XOR2_X1 U217 (.Z(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module up_island_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [31:0] A;
   input [31:0] B;
   input CI;
   output [31:0] DIFF;
   output CO;

   // Internal wires
   wire \carry[31] ;
   wire \carry[30] ;
   wire \carry[29] ;
   wire \carry[28] ;
   wire \carry[27] ;
   wire \carry[24] ;
   wire \carry[23] ;
   wire \carry[22] ;
   wire \carry[21] ;
   wire \carry[20] ;
   wire \carry[19] ;
   wire \carry[18] ;
   wire \carry[17] ;
   wire \carry[16] ;
   wire \carry[15] ;
   wire \carry[13] ;
   wire \carry[11] ;
   wire \carry[10] ;
   wire \carry[9] ;
   wire \carry[8] ;
   wire \carry[6] ;
   wire \carry[5] ;
   wire \carry[2] ;
   wire \carry[1] ;
   wire \B_not[31] ;
   wire \B_not[30] ;
   wire \B_not[29] ;
   wire \B_not[28] ;
   wire \B_not[27] ;
   wire \B_not[26] ;
   wire \B_not[25] ;
   wire \B_not[24] ;
   wire \B_not[23] ;
   wire \B_not[22] ;
   wire \B_not[21] ;
   wire \B_not[20] ;
   wire \B_not[19] ;
   wire \B_not[18] ;
   wire \B_not[17] ;
   wire \B_not[16] ;
   wire \B_not[15] ;
   wire \B_not[14] ;
   wire \B_not[13] ;
   wire \B_not[12] ;
   wire \B_not[11] ;
   wire \B_not[10] ;
   wire \B_not[9] ;
   wire \B_not[8] ;
   wire \B_not[7] ;
   wire \B_not[6] ;
   wire \B_not[5] ;
   wire n1;
   wire n2;
   wire n7;
   wire n8;
   wire n9;
   wire n12;
   wire n14;
   wire n16;
   wire n21;
   wire n23;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n40;
   wire n44;
   wire n45;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n53;
   wire n54;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n64;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n87;
   wire n88;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;

   FA_X1 U2_18 (.S(DIFF[18]), 
	.CO(\carry[19] ), 
	.CI(\carry[18] ), 
	.B(\B_not[18] ), 
	.A(A[18]));
   FA_X1 U2_15 (.S(DIFF[15]), 
	.CO(\carry[16] ), 
	.CI(\carry[15] ), 
	.B(\B_not[15] ), 
	.A(A[15]));
   NAND2_X1 U1 (.ZN(n109), 
	.A2(A[9]), 
	.A1(\B_not[9] ));
   NAND2_X1 U2 (.ZN(n113), 
	.A2(A[10]), 
	.A1(\B_not[10] ));
   NAND2_X1 U3 (.ZN(n34), 
	.A2(\B_not[22] ), 
	.A1(A[22]));
   NAND2_X1 U4 (.ZN(n169), 
	.A2(A[23]), 
	.A1(\B_not[23] ));
   NAND2_X1 U5 (.ZN(n160), 
	.A2(A[8]), 
	.A1(\B_not[8] ));
   NAND2_X1 U6 (.ZN(n80), 
	.A2(A[16]), 
	.A1(\B_not[16] ));
   NAND2_X1 U7 (.ZN(n173), 
	.A2(A[17]), 
	.A1(\B_not[17] ));
   NAND2_X1 U8 (.ZN(n164), 
	.A2(A[7]), 
	.A1(\B_not[7] ));
   NAND2_X1 U9 (.ZN(n156), 
	.A2(A[14]), 
	.A1(\B_not[14] ));
   NAND2_X1 U10 (.ZN(n148), 
	.A2(A[13]), 
	.A1(\B_not[13] ));
   NAND2_X1 U11 (.ZN(n105), 
	.A2(A[11]), 
	.A1(\B_not[11] ));
   NAND2_X1 U12 (.ZN(n140), 
	.A2(A[12]), 
	.A1(\B_not[12] ));
   NAND2_X1 U13 (.ZN(n123), 
	.A2(\B_not[24] ), 
	.A1(A[24]));
   NAND2_X1 U14 (.ZN(n144), 
	.A2(A[6]), 
	.A1(\B_not[6] ));
   INV_X1 U15 (.ZN(n72), 
	.A(n118));
   NAND2_X1 U17 (.ZN(n1), 
	.A2(\B_not[12] ), 
	.A1(n64));
   NAND2_X1 U18 (.ZN(n125), 
	.A2(\B_not[24] ), 
	.A1(n71));
   NAND2_X1 U19 (.ZN(n2), 
	.A2(A[24]), 
	.A1(\carry[24] ));
   NAND3_X1 U24 (.ZN(\carry[8] ), 
	.A3(n162), 
	.A2(n164), 
	.A1(n163));
   NAND2_X1 U25 (.ZN(n147), 
	.A2(A[13]), 
	.A1(\carry[13] ));
   NAND3_X1 U26 (.ZN(\carry[6] ), 
	.A3(n100), 
	.A2(n102), 
	.A1(n101));
   NAND2_X1 U28 (.ZN(n7), 
	.A2(A[11]), 
	.A1(\carry[11] ));
   NAND2_X1 U29 (.ZN(n8), 
	.A2(\B_not[11] ), 
	.A1(n29));
   NAND2_X1 U30 (.ZN(n146), 
	.A2(\B_not[13] ), 
	.A1(n87));
   NAND3_X1 U31 (.ZN(\carry[10] ), 
	.A3(n107), 
	.A2(n109), 
	.A1(n108));
   NAND3_X1 U32 (.ZN(n9), 
	.A3(n158), 
	.A2(n160), 
	.A1(n159));
   NAND2_X1 U35 (.ZN(n12), 
	.A2(A[3]), 
	.A1(n21));
   NAND3_X1 U37 (.ZN(n14), 
	.A3(n146), 
	.A2(n148), 
	.A1(n147));
   NAND3_X1 U39 (.ZN(n16), 
	.A3(n69), 
	.A2(n68), 
	.A1(n67));
   NAND3_X1 U44 (.ZN(\carry[23] ), 
	.A3(n33), 
	.A2(n34), 
	.A1(n32));
   NAND3_X1 U45 (.ZN(\carry[9] ), 
	.A3(n160), 
	.A2(n158), 
	.A1(n159));
   NAND3_X1 U46 (.ZN(n21), 
	.A3(n133), 
	.A2(n131), 
	.A1(n132));
   NAND2_X1 U49 (.ZN(n23), 
	.A2(\B_not[25] ), 
	.A1(n90));
   NAND3_X1 U52 (.ZN(n26), 
	.A3(n94), 
	.A2(n93), 
	.A1(n92));
   NAND3_X1 U53 (.ZN(n27), 
	.A3(n98), 
	.A2(n97), 
	.A1(n96));
   NAND3_X1 U54 (.ZN(\carry[22] ), 
	.A3(n93), 
	.A2(n94), 
	.A1(n92));
   NAND3_X1 U55 (.ZN(\carry[5] ), 
	.A3(n59), 
	.A2(n60), 
	.A1(n58));
   NAND3_X1 U56 (.ZN(n28), 
	.A3(n115), 
	.A2(n117), 
	.A1(n12));
   NAND3_X1 U57 (.ZN(n29), 
	.A3(n111), 
	.A2(n113), 
	.A1(n112));
   XOR2_X1 U59 (.Z(n31), 
	.B(\B_not[22] ), 
	.A(A[22]));
   XOR2_X1 U60 (.Z(DIFF[22]), 
	.B(n31), 
	.A(n26));
   NAND2_X1 U61 (.ZN(n32), 
	.A2(A[22]), 
	.A1(n26));
   NAND2_X1 U62 (.ZN(n33), 
	.A2(\B_not[22] ), 
	.A1(\carry[22] ));
   NAND3_X1 U63 (.ZN(n35), 
	.A3(n49), 
	.A2(n50), 
	.A1(n48));
   INV_X1 U64 (.ZN(\B_not[22] ), 
	.A(B[22]));
   AND3_X1 U65 (.ZN(n40), 
	.A3(n152), 
	.A2(n151), 
	.A1(n150));
   NAND3_X1 U67 (.ZN(\carry[11] ), 
	.A3(n113), 
	.A2(n111), 
	.A1(n112));
   NAND2_X1 U68 (.ZN(n111), 
	.A2(\B_not[10] ), 
	.A1(\carry[10] ));
   XNOR2_X1 U69 (.ZN(DIFF[31]), 
	.B(n45), 
	.A(\carry[31] ));
   XNOR2_X1 U73 (.ZN(DIFF[30]), 
	.B(n134), 
	.A(n40));
   XNOR2_X1 U78 (.ZN(DIFF[28]), 
	.B(n81), 
	.A(n44));
   AND3_X1 U79 (.ZN(n44), 
	.A3(n121), 
	.A2(n120), 
	.A1(n119));
   XNOR2_X1 U80 (.ZN(n45), 
	.B(\B_not[31] ), 
	.A(A[31]));
   XOR2_X1 U81 (.Z(n47), 
	.B(\B_not[19] ), 
	.A(A[19]));
   XOR2_X1 U82 (.Z(DIFF[19]), 
	.B(n47), 
	.A(\carry[19] ));
   NAND2_X1 U83 (.ZN(n48), 
	.A2(A[19]), 
	.A1(\carry[19] ));
   NAND2_X1 U84 (.ZN(n49), 
	.A2(\B_not[19] ), 
	.A1(\carry[19] ));
   NAND2_X1 U85 (.ZN(n50), 
	.A2(\B_not[19] ), 
	.A1(A[19]));
   NAND3_X1 U86 (.ZN(\carry[20] ), 
	.A3(n50), 
	.A2(n49), 
	.A1(n48));
   NAND3_X1 U89 (.ZN(n53), 
	.A3(n23), 
	.A2(n127), 
	.A1(n128));
   NAND3_X1 U90 (.ZN(n54), 
	.A3(n78), 
	.A2(n80), 
	.A1(n79));
   NAND3_X1 U92 (.ZN(n56), 
	.A3(n142), 
	.A2(n144), 
	.A1(n143));
   XOR2_X1 U93 (.Z(n57), 
	.B(n174), 
	.A(A[4]));
   XOR2_X1 U94 (.Z(DIFF[4]), 
	.B(n57), 
	.A(n28));
   NAND2_X1 U95 (.ZN(n58), 
	.A2(A[4]), 
	.A1(n28));
   NAND2_X1 U96 (.ZN(n59), 
	.A2(n174), 
	.A1(n28));
   NAND2_X1 U97 (.ZN(n60), 
	.A2(n174), 
	.A1(A[4]));
   NAND3_X1 U98 (.ZN(n61), 
	.A3(n83), 
	.A2(n84), 
	.A1(n82));
   NAND3_X1 U99 (.ZN(\carry[17] ), 
	.A3(n79), 
	.A2(n80), 
	.A1(n78));
   NAND3_X1 U102 (.ZN(n64), 
	.A3(n7), 
	.A2(n105), 
	.A1(n8));
   XOR2_X1 U104 (.Z(n66), 
	.B(\B_not[26] ), 
	.A(A[26]));
   XOR2_X1 U105 (.Z(DIFF[26]), 
	.B(n66), 
	.A(n53));
   NAND2_X1 U106 (.ZN(n67), 
	.A2(A[26]), 
	.A1(n53));
   NAND2_X1 U107 (.ZN(n68), 
	.A2(\B_not[26] ), 
	.A1(n53));
   NAND2_X1 U108 (.ZN(n69), 
	.A2(\B_not[26] ), 
	.A1(A[26]));
   NAND3_X1 U109 (.ZN(\carry[27] ), 
	.A3(n68), 
	.A2(n69), 
	.A1(n67));
   NAND3_X1 U110 (.ZN(n70), 
	.A3(n75), 
	.A2(n76), 
	.A1(n74));
   NAND3_X1 U111 (.ZN(n71), 
	.A3(n168), 
	.A2(n169), 
	.A1(n167));
   XNOR2_X1 U113 (.ZN(DIFF[27]), 
	.B(n72), 
	.A(n16));
   XOR2_X1 U114 (.Z(n73), 
	.B(\B_not[20] ), 
	.A(A[20]));
   XOR2_X1 U115 (.Z(DIFF[20]), 
	.B(n73), 
	.A(n35));
   NAND2_X1 U116 (.ZN(n74), 
	.A2(A[20]), 
	.A1(\carry[20] ));
   NAND2_X1 U117 (.ZN(n75), 
	.A2(\B_not[20] ), 
	.A1(\carry[20] ));
   NAND2_X1 U118 (.ZN(n76), 
	.A2(\B_not[20] ), 
	.A1(A[20]));
   NAND3_X1 U119 (.ZN(\carry[21] ), 
	.A3(n76), 
	.A2(n75), 
	.A1(n74));
   XOR2_X1 U120 (.Z(n77), 
	.B(A[16]), 
	.A(\B_not[16] ));
   XOR2_X1 U121 (.Z(DIFF[16]), 
	.B(n77), 
	.A(\carry[16] ));
   NAND2_X1 U122 (.ZN(n78), 
	.A2(\B_not[16] ), 
	.A1(\carry[16] ));
   NAND2_X1 U123 (.ZN(n79), 
	.A2(A[16]), 
	.A1(\carry[16] ));
   XOR2_X1 U124 (.Z(n81), 
	.B(\B_not[28] ), 
	.A(A[28]));
   NAND2_X1 U125 (.ZN(n82), 
	.A2(A[28]), 
	.A1(\carry[28] ));
   NAND2_X1 U126 (.ZN(n83), 
	.A2(\B_not[28] ), 
	.A1(\carry[28] ));
   NAND2_X1 U127 (.ZN(n84), 
	.A2(\B_not[28] ), 
	.A1(A[28]));
   NAND3_X1 U128 (.ZN(\carry[29] ), 
	.A3(n84), 
	.A2(n83), 
	.A1(n82));
   NAND3_X1 U131 (.ZN(n87), 
	.A3(n1), 
	.A2(n140), 
	.A1(n139));
   NAND3_X1 U132 (.ZN(n88), 
	.A3(n147), 
	.A2(n148), 
	.A1(n146));
   NAND3_X1 U134 (.ZN(n90), 
	.A3(n125), 
	.A2(n123), 
	.A1(n2));
   XOR2_X1 U135 (.Z(n91), 
	.B(\B_not[21] ), 
	.A(A[21]));
   XOR2_X1 U136 (.Z(DIFF[21]), 
	.B(n91), 
	.A(n70));
   NAND2_X1 U137 (.ZN(n92), 
	.A2(A[21]), 
	.A1(\carry[21] ));
   NAND2_X1 U138 (.ZN(n93), 
	.A2(\B_not[21] ), 
	.A1(\carry[21] ));
   NAND2_X1 U139 (.ZN(n94), 
	.A2(\B_not[21] ), 
	.A1(A[21]));
   XOR2_X1 U140 (.Z(n95), 
	.B(A[1]), 
	.A(n177));
   XOR2_X1 U141 (.Z(DIFF[1]), 
	.B(n95), 
	.A(\carry[1] ));
   NAND2_X1 U142 (.ZN(n96), 
	.A2(n177), 
	.A1(\carry[1] ));
   NAND2_X1 U143 (.ZN(n97), 
	.A2(A[1]), 
	.A1(\carry[1] ));
   NAND2_X1 U144 (.ZN(n98), 
	.A2(A[1]), 
	.A1(n177));
   NAND3_X1 U145 (.ZN(\carry[2] ), 
	.A3(n96), 
	.A2(n98), 
	.A1(n97));
   NAND3_X1 U146 (.ZN(\carry[13] ), 
	.A3(n140), 
	.A2(n139), 
	.A1(n1));
   INV_X1 U150 (.ZN(\B_not[21] ), 
	.A(B[21]));
   OR2_X1 U151 (.ZN(\carry[1] ), 
	.A2(A[0]), 
	.A1(n165));
   NAND2_X1 U152 (.ZN(n162), 
	.A2(\B_not[7] ), 
	.A1(n56));
   XOR2_X1 U153 (.Z(n99), 
	.B(A[5]), 
	.A(\B_not[5] ));
   XOR2_X1 U154 (.Z(DIFF[5]), 
	.B(n99), 
	.A(\carry[5] ));
   NAND2_X1 U155 (.ZN(n100), 
	.A2(\B_not[5] ), 
	.A1(\carry[5] ));
   NAND2_X1 U156 (.ZN(n101), 
	.A2(A[5]), 
	.A1(\carry[5] ));
   NAND2_X1 U157 (.ZN(n102), 
	.A2(A[5]), 
	.A1(\B_not[5] ));
   XOR2_X1 U158 (.Z(n103), 
	.B(A[11]), 
	.A(\B_not[11] ));
   XOR2_X1 U159 (.Z(DIFF[11]), 
	.B(n103), 
	.A(n29));
   INV_X1 U161 (.ZN(\B_not[11] ), 
	.A(B[11]));
   XOR2_X1 U162 (.Z(n106), 
	.B(A[9]), 
	.A(\B_not[9] ));
   XOR2_X1 U163 (.Z(DIFF[9]), 
	.B(n106), 
	.A(\carry[9] ));
   NAND2_X1 U164 (.ZN(n107), 
	.A2(\B_not[9] ), 
	.A1(n9));
   NAND2_X1 U165 (.ZN(n108), 
	.A2(A[9]), 
	.A1(\carry[9] ));
   XOR2_X1 U166 (.Z(n110), 
	.B(A[10]), 
	.A(\B_not[10] ));
   XOR2_X1 U167 (.Z(DIFF[10]), 
	.B(n110), 
	.A(\carry[10] ));
   NAND2_X1 U168 (.ZN(n112), 
	.A2(A[10]), 
	.A1(\carry[10] ));
   XOR2_X1 U169 (.Z(n114), 
	.B(A[3]), 
	.A(n175));
   XOR2_X1 U170 (.Z(DIFF[3]), 
	.B(n114), 
	.A(n21));
   NAND2_X1 U171 (.ZN(n115), 
	.A2(n175), 
	.A1(n21));
   NAND2_X1 U173 (.ZN(n117), 
	.A2(A[3]), 
	.A1(n175));
   XOR2_X1 U174 (.Z(n118), 
	.B(\B_not[27] ), 
	.A(A[27]));
   NAND2_X1 U175 (.ZN(n119), 
	.A2(A[27]), 
	.A1(\carry[27] ));
   NAND2_X1 U176 (.ZN(n120), 
	.A2(\B_not[27] ), 
	.A1(n16));
   NAND2_X1 U177 (.ZN(n121), 
	.A2(\B_not[27] ), 
	.A1(A[27]));
   NAND3_X1 U178 (.ZN(\carry[28] ), 
	.A3(n121), 
	.A2(n120), 
	.A1(n119));
   XOR2_X1 U179 (.Z(n122), 
	.B(\B_not[24] ), 
	.A(A[24]));
   XOR2_X1 U180 (.Z(DIFF[24]), 
	.B(n122), 
	.A(\carry[24] ));
   XOR2_X1 U181 (.Z(n126), 
	.B(\B_not[25] ), 
	.A(A[25]));
   XOR2_X1 U182 (.Z(DIFF[25]), 
	.B(n90), 
	.A(n126));
   NAND2_X1 U183 (.ZN(n127), 
	.A2(\B_not[25] ), 
	.A1(A[25]));
   NAND2_X1 U184 (.ZN(n128), 
	.A2(A[25]), 
	.A1(n90));
   XOR2_X1 U187 (.Z(n130), 
	.B(A[2]), 
	.A(n176));
   XOR2_X1 U188 (.Z(DIFF[2]), 
	.B(n130), 
	.A(n27));
   NAND2_X1 U189 (.ZN(n131), 
	.A2(n176), 
	.A1(\carry[2] ));
   NAND2_X1 U190 (.ZN(n132), 
	.A2(A[2]), 
	.A1(n27));
   NAND2_X1 U191 (.ZN(n133), 
	.A2(A[2]), 
	.A1(n176));
   XOR2_X1 U192 (.Z(n134), 
	.B(\B_not[30] ), 
	.A(A[30]));
   NAND2_X1 U193 (.ZN(n135), 
	.A2(A[30]), 
	.A1(\carry[30] ));
   NAND2_X1 U194 (.ZN(n136), 
	.A2(\B_not[30] ), 
	.A1(\carry[30] ));
   NAND2_X1 U195 (.ZN(n137), 
	.A2(\B_not[30] ), 
	.A1(A[30]));
   NAND3_X1 U196 (.ZN(\carry[31] ), 
	.A3(n137), 
	.A2(n136), 
	.A1(n135));
   XOR2_X1 U197 (.Z(n138), 
	.B(A[12]), 
	.A(\B_not[12] ));
   XOR2_X1 U198 (.Z(DIFF[12]), 
	.B(n138), 
	.A(n64));
   NAND2_X1 U199 (.ZN(n139), 
	.A2(A[12]), 
	.A1(n64));
   XOR2_X1 U200 (.Z(n141), 
	.B(A[6]), 
	.A(\B_not[6] ));
   XOR2_X1 U201 (.Z(DIFF[6]), 
	.B(n141), 
	.A(\carry[6] ));
   NAND2_X1 U202 (.ZN(n142), 
	.A2(\B_not[6] ), 
	.A1(\carry[6] ));
   NAND2_X1 U203 (.ZN(n143), 
	.A2(A[6]), 
	.A1(\carry[6] ));
   INV_X1 U204 (.ZN(\B_not[30] ), 
	.A(B[30]));
   XOR2_X1 U205 (.Z(n145), 
	.B(A[13]), 
	.A(\B_not[13] ));
   XOR2_X1 U206 (.Z(DIFF[13]), 
	.B(n145), 
	.A(\carry[13] ));
   XOR2_X1 U207 (.Z(n149), 
	.B(\B_not[29] ), 
	.A(A[29]));
   XOR2_X1 U208 (.Z(DIFF[29]), 
	.B(n149), 
	.A(n61));
   NAND2_X1 U209 (.ZN(n150), 
	.A2(A[29]), 
	.A1(\carry[29] ));
   NAND2_X1 U210 (.ZN(n151), 
	.A2(\B_not[29] ), 
	.A1(\carry[29] ));
   NAND2_X1 U211 (.ZN(n152), 
	.A2(\B_not[29] ), 
	.A1(A[29]));
   NAND3_X1 U212 (.ZN(\carry[30] ), 
	.A3(n152), 
	.A2(n151), 
	.A1(n150));
   XOR2_X1 U213 (.Z(n153), 
	.B(A[14]), 
	.A(\B_not[14] ));
   XOR2_X1 U214 (.Z(DIFF[14]), 
	.B(n153), 
	.A(n88));
   NAND2_X1 U215 (.ZN(n154), 
	.A2(\B_not[14] ), 
	.A1(n14));
   NAND2_X1 U216 (.ZN(n155), 
	.A2(A[14]), 
	.A1(n14));
   NAND3_X1 U217 (.ZN(\carry[15] ), 
	.A3(n154), 
	.A2(n156), 
	.A1(n155));
   XOR2_X1 U218 (.Z(n157), 
	.B(A[8]), 
	.A(\B_not[8] ));
   XOR2_X1 U219 (.Z(DIFF[8]), 
	.B(n157), 
	.A(\carry[8] ));
   NAND2_X1 U220 (.ZN(n158), 
	.A2(\B_not[8] ), 
	.A1(\carry[8] ));
   NAND2_X1 U221 (.ZN(n159), 
	.A2(A[8]), 
	.A1(\carry[8] ));
   XOR2_X1 U222 (.Z(n161), 
	.B(A[7]), 
	.A(\B_not[7] ));
   XOR2_X1 U223 (.Z(DIFF[7]), 
	.B(n161), 
	.A(n56));
   NAND2_X1 U224 (.ZN(n163), 
	.A2(A[7]), 
	.A1(n56));
   INV_X1 U225 (.ZN(\B_not[29] ), 
	.A(B[29]));
   INV_X1 U226 (.ZN(n165), 
	.A(B[0]));
   XOR2_X1 U227 (.Z(n166), 
	.B(A[23]), 
	.A(\B_not[23] ));
   XOR2_X1 U228 (.Z(DIFF[23]), 
	.B(n166), 
	.A(\carry[23] ));
   NAND2_X1 U229 (.ZN(n167), 
	.A2(\B_not[23] ), 
	.A1(\carry[23] ));
   NAND2_X1 U230 (.ZN(n168), 
	.A2(A[23]), 
	.A1(\carry[23] ));
   NAND3_X1 U231 (.ZN(\carry[24] ), 
	.A3(n169), 
	.A2(n167), 
	.A1(n168));
   XOR2_X1 U232 (.Z(n170), 
	.B(A[17]), 
	.A(\B_not[17] ));
   XOR2_X1 U233 (.Z(DIFF[17]), 
	.B(n170), 
	.A(n54));
   NAND2_X1 U234 (.ZN(n171), 
	.A2(\B_not[17] ), 
	.A1(\carry[17] ));
   NAND2_X1 U235 (.ZN(n172), 
	.A2(A[17]), 
	.A1(\carry[17] ));
   NAND3_X1 U236 (.ZN(\carry[18] ), 
	.A3(n173), 
	.A2(n171), 
	.A1(n172));
   INV_X1 U237 (.ZN(n174), 
	.A(B[4]));
   INV_X1 U238 (.ZN(n175), 
	.A(B[3]));
   INV_X1 U239 (.ZN(n176), 
	.A(B[2]));
   INV_X1 U240 (.ZN(n177), 
	.A(B[1]));
   XNOR2_X1 U242 (.ZN(DIFF[0]), 
	.B(n165), 
	.A(A[0]));
   INV_X1 U243 (.ZN(\B_not[9] ), 
	.A(B[9]));
   INV_X1 U244 (.ZN(\B_not[8] ), 
	.A(B[8]));
   INV_X1 U245 (.ZN(\B_not[7] ), 
	.A(B[7]));
   INV_X1 U246 (.ZN(\B_not[6] ), 
	.A(B[6]));
   INV_X1 U247 (.ZN(\B_not[5] ), 
	.A(B[5]));
   INV_X1 U248 (.ZN(\B_not[31] ), 
	.A(B[31]));
   INV_X1 U249 (.ZN(\B_not[28] ), 
	.A(B[28]));
   INV_X1 U250 (.ZN(\B_not[27] ), 
	.A(B[27]));
   INV_X1 U251 (.ZN(\B_not[26] ), 
	.A(B[26]));
   INV_X1 U252 (.ZN(\B_not[25] ), 
	.A(B[25]));
   INV_X1 U253 (.ZN(\B_not[24] ), 
	.A(B[24]));
   INV_X1 U254 (.ZN(\B_not[23] ), 
	.A(B[23]));
   INV_X1 U255 (.ZN(\B_not[20] ), 
	.A(B[20]));
   INV_X1 U256 (.ZN(\B_not[19] ), 
	.A(B[19]));
   INV_X1 U257 (.ZN(\B_not[18] ), 
	.A(B[18]));
   INV_X1 U258 (.ZN(\B_not[17] ), 
	.A(B[17]));
   INV_X1 U259 (.ZN(\B_not[16] ), 
	.A(B[16]));
   INV_X1 U260 (.ZN(\B_not[15] ), 
	.A(B[15]));
   INV_X1 U261 (.ZN(\B_not[14] ), 
	.A(B[14]));
   INV_X1 U262 (.ZN(\B_not[13] ), 
	.A(B[13]));
   INV_X1 U263 (.ZN(\B_not[12] ), 
	.A(B[12]));
   INV_X1 U264 (.ZN(\B_not[10] ), 
	.A(B[10]));
endmodule

module up_island_DW01_cmp6_0 (
	A, 
	B, 
	TC, 
	LT, 
	GT, 
	EQ, 
	LE, 
	GE, 
	NE, 
	n6832);
   input [31:0] A;
   input [31:0] B;
   input TC;
   output LT;
   output GT;
   output EQ;
   output LE;
   output GE;
   output NE;
   input n6832;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;

   AND4_X1 U1 (.ZN(n6), 
	.A4(n4), 
	.A3(n3), 
	.A2(n2), 
	.A1(n1));
   AND4_X1 U2 (.ZN(n1), 
	.A4(n22), 
	.A3(n21), 
	.A2(n20), 
	.A1(n19));
   AND4_X1 U3 (.ZN(n2), 
	.A4(n18), 
	.A3(n17), 
	.A2(n16), 
	.A1(n15));
   AND4_X1 U4 (.ZN(n3), 
	.A4(n14), 
	.A3(n13), 
	.A2(n12), 
	.A1(n11));
   AND4_X1 U5 (.ZN(n4), 
	.A4(n10), 
	.A3(n9), 
	.A2(n8), 
	.A1(n7));
   INV_X1 U6 (.ZN(EQ), 
	.A(NE));
   NAND2_X1 U7 (.ZN(NE), 
	.A2(n6), 
	.A1(n5));
   XNOR2_X1 U8 (.ZN(n10), 
	.B(A[11]), 
	.A(B[11]));
   XNOR2_X1 U9 (.ZN(n9), 
	.B(A[12]), 
	.A(B[12]));
   XNOR2_X1 U10 (.ZN(n8), 
	.B(A[13]), 
	.A(B[13]));
   XNOR2_X1 U11 (.ZN(n7), 
	.B(A[14]), 
	.A(B[14]));
   XNOR2_X1 U12 (.ZN(n14), 
	.B(A[7]), 
	.A(B[7]));
   XNOR2_X1 U13 (.ZN(n13), 
	.B(A[8]), 
	.A(B[8]));
   XNOR2_X1 U14 (.ZN(n12), 
	.B(A[9]), 
	.A(B[9]));
   XNOR2_X1 U15 (.ZN(n11), 
	.B(A[10]), 
	.A(B[10]));
   XNOR2_X1 U16 (.ZN(n18), 
	.B(A[3]), 
	.A(B[3]));
   XNOR2_X1 U17 (.ZN(n17), 
	.B(A[4]), 
	.A(B[4]));
   XNOR2_X1 U18 (.ZN(n16), 
	.B(A[5]), 
	.A(B[5]));
   XNOR2_X1 U19 (.ZN(n15), 
	.B(A[6]), 
	.A(B[6]));
   OAI22_X1 U20 (.ZN(n22), 
	.B2(n23), 
	.B1(B[1]), 
	.A2(n24), 
	.A1(n23));
   INV_X1 U21 (.ZN(n24), 
	.A(A[1]));
   AND2_X1 U22 (.ZN(n23), 
	.A2(n6832), 
	.A1(B[0]));
   OAI22_X1 U23 (.ZN(n21), 
	.B2(n27), 
	.B1(n26), 
	.A2(n26), 
	.A1(A[1]));
   INV_X1 U24 (.ZN(n27), 
	.A(B[1]));
   NOR2_X1 U25 (.ZN(n26), 
	.A2(B[0]), 
	.A1(n6832));
   XNOR2_X1 U27 (.ZN(n20), 
	.B(A[31]), 
	.A(B[31]));
   XNOR2_X1 U28 (.ZN(n19), 
	.B(A[2]), 
	.A(B[2]));
   NOR4_X1 U29 (.ZN(n5), 
	.A4(n31), 
	.A3(n30), 
	.A2(n29), 
	.A1(n28));
   NAND4_X1 U30 (.ZN(n31), 
	.A4(n35), 
	.A3(n34), 
	.A2(n33), 
	.A1(n32));
   XNOR2_X1 U31 (.ZN(n35), 
	.B(A[27]), 
	.A(B[27]));
   XNOR2_X1 U32 (.ZN(n34), 
	.B(A[28]), 
	.A(B[28]));
   XNOR2_X1 U33 (.ZN(n33), 
	.B(A[29]), 
	.A(B[29]));
   XNOR2_X1 U34 (.ZN(n32), 
	.B(A[30]), 
	.A(B[30]));
   NAND4_X1 U35 (.ZN(n30), 
	.A4(n39), 
	.A3(n38), 
	.A2(n37), 
	.A1(n36));
   XNOR2_X1 U36 (.ZN(n39), 
	.B(A[23]), 
	.A(B[23]));
   XNOR2_X1 U37 (.ZN(n38), 
	.B(A[24]), 
	.A(B[24]));
   XNOR2_X1 U38 (.ZN(n37), 
	.B(A[25]), 
	.A(B[25]));
   XNOR2_X1 U39 (.ZN(n36), 
	.B(A[26]), 
	.A(B[26]));
   NAND4_X1 U40 (.ZN(n29), 
	.A4(n43), 
	.A3(n42), 
	.A2(n41), 
	.A1(n40));
   XNOR2_X1 U41 (.ZN(n43), 
	.B(A[19]), 
	.A(B[19]));
   XNOR2_X1 U42 (.ZN(n42), 
	.B(A[20]), 
	.A(B[20]));
   XNOR2_X1 U43 (.ZN(n41), 
	.B(A[21]), 
	.A(B[21]));
   XNOR2_X1 U44 (.ZN(n40), 
	.B(A[22]), 
	.A(B[22]));
   NAND4_X1 U45 (.ZN(n28), 
	.A4(n47), 
	.A3(n46), 
	.A2(n45), 
	.A1(n44));
   XNOR2_X1 U46 (.ZN(n47), 
	.B(A[15]), 
	.A(B[15]));
   XNOR2_X1 U47 (.ZN(n46), 
	.B(A[16]), 
	.A(B[16]));
   XNOR2_X1 U48 (.ZN(n45), 
	.B(A[17]), 
	.A(B[17]));
   XNOR2_X1 U49 (.ZN(n44), 
	.B(A[18]), 
	.A(B[18]));
endmodule

module up_island_DW01_add_2 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [24:0] A;
   input [24:0] B;
   input CI;
   output [24:0] SUM;
   output CO;

   // Internal wires
   wire \A[1] ;
   wire \A[0] ;
   wire \carry[23] ;
   wire \carry[22] ;
   wire \carry[21] ;
   wire \carry[20] ;
   wire \carry[19] ;
   wire \carry[18] ;
   wire \carry[17] ;
   wire \carry[16] ;
   wire \carry[15] ;
   wire \carry[14] ;
   wire \carry[13] ;
   wire \carry[12] ;
   wire \carry[11] ;
   wire \carry[10] ;
   wire \carry[9] ;
   wire \carry[8] ;
   wire \carry[7] ;
   wire \carry[6] ;
   wire \carry[5] ;
   wire \carry[4] ;
   wire \carry[3] ;

   assign SUM[1] = \A[1]  ;
   assign \A[1]  = A[1] ;
   assign SUM[0] = \A[0]  ;
   assign \A[0]  = A[0] ;
   assign \carry[3]  = A[2] ;

   XOR2_X1 U1 (.Z(SUM[20]), 
	.B(\carry[20] ), 
	.A(A[20]));
   XOR2_X1 U2 (.Z(SUM[17]), 
	.B(\carry[17] ), 
	.A(A[17]));
   XOR2_X1 U3 (.Z(SUM[22]), 
	.B(\carry[22] ), 
	.A(A[22]));
   XOR2_X1 U4 (.Z(SUM[19]), 
	.B(\carry[19] ), 
	.A(A[19]));
   XOR2_X1 U5 (.Z(SUM[21]), 
	.B(\carry[21] ), 
	.A(A[21]));
   XOR2_X1 U6 (.Z(SUM[15]), 
	.B(\carry[15] ), 
	.A(A[15]));
   XOR2_X1 U7 (.Z(SUM[23]), 
	.B(\carry[23] ), 
	.A(A[23]));
   AND2_X1 U8 (.ZN(\carry[23] ), 
	.A2(A[22]), 
	.A1(\carry[22] ));
   AND2_X1 U9 (.ZN(\carry[22] ), 
	.A2(A[21]), 
	.A1(\carry[21] ));
   AND2_X1 U10 (.ZN(\carry[21] ), 
	.A2(A[20]), 
	.A1(\carry[20] ));
   AND2_X1 U11 (.ZN(\carry[20] ), 
	.A2(A[19]), 
	.A1(\carry[19] ));
   AND2_X1 U12 (.ZN(\carry[19] ), 
	.A2(A[18]), 
	.A1(\carry[18] ));
   XOR2_X1 U13 (.Z(SUM[18]), 
	.B(\carry[18] ), 
	.A(A[18]));
   AND2_X1 U14 (.ZN(\carry[18] ), 
	.A2(A[17]), 
	.A1(\carry[17] ));
   AND2_X1 U15 (.ZN(\carry[17] ), 
	.A2(A[16]), 
	.A1(\carry[16] ));
   XOR2_X1 U16 (.Z(SUM[16]), 
	.B(\carry[16] ), 
	.A(A[16]));
   AND2_X1 U17 (.ZN(\carry[16] ), 
	.A2(A[15]), 
	.A1(\carry[15] ));
   AND2_X1 U18 (.ZN(\carry[15] ), 
	.A2(A[14]), 
	.A1(\carry[14] ));
   XOR2_X1 U19 (.Z(SUM[14]), 
	.B(\carry[14] ), 
	.A(A[14]));
   AND2_X1 U20 (.ZN(\carry[14] ), 
	.A2(A[13]), 
	.A1(\carry[13] ));
   XOR2_X1 U21 (.Z(SUM[13]), 
	.B(\carry[13] ), 
	.A(A[13]));
   AND2_X1 U22 (.ZN(\carry[13] ), 
	.A2(A[12]), 
	.A1(\carry[12] ));
   XOR2_X1 U23 (.Z(SUM[12]), 
	.B(\carry[12] ), 
	.A(A[12]));
   AND2_X1 U24 (.ZN(\carry[12] ), 
	.A2(A[11]), 
	.A1(\carry[11] ));
   XOR2_X1 U25 (.Z(SUM[11]), 
	.B(\carry[11] ), 
	.A(A[11]));
   AND2_X1 U26 (.ZN(\carry[11] ), 
	.A2(A[10]), 
	.A1(\carry[10] ));
   XOR2_X1 U27 (.Z(SUM[10]), 
	.B(\carry[10] ), 
	.A(A[10]));
   AND2_X1 U28 (.ZN(\carry[10] ), 
	.A2(A[9]), 
	.A1(\carry[9] ));
   XOR2_X1 U29 (.Z(SUM[9]), 
	.B(\carry[9] ), 
	.A(A[9]));
   AND2_X1 U30 (.ZN(\carry[9] ), 
	.A2(A[8]), 
	.A1(\carry[8] ));
   XOR2_X1 U31 (.Z(SUM[8]), 
	.B(\carry[8] ), 
	.A(A[8]));
   AND2_X1 U32 (.ZN(\carry[8] ), 
	.A2(A[7]), 
	.A1(\carry[7] ));
   XOR2_X1 U33 (.Z(SUM[7]), 
	.B(\carry[7] ), 
	.A(A[7]));
   AND2_X1 U34 (.ZN(\carry[7] ), 
	.A2(A[6]), 
	.A1(\carry[6] ));
   XOR2_X1 U35 (.Z(SUM[6]), 
	.B(\carry[6] ), 
	.A(A[6]));
   AND2_X1 U36 (.ZN(\carry[6] ), 
	.A2(A[5]), 
	.A1(\carry[5] ));
   XOR2_X1 U37 (.Z(SUM[5]), 
	.B(\carry[5] ), 
	.A(A[5]));
   AND2_X1 U38 (.ZN(\carry[5] ), 
	.A2(A[4]), 
	.A1(\carry[4] ));
   XOR2_X1 U39 (.Z(SUM[4]), 
	.B(\carry[4] ), 
	.A(A[4]));
   AND2_X1 U40 (.ZN(\carry[4] ), 
	.A2(A[3]), 
	.A1(\carry[3] ));
   XOR2_X1 U41 (.Z(SUM[3]), 
	.B(\carry[3] ), 
	.A(A[3]));
   INV_X1 U42 (.ZN(SUM[2]), 
	.A(\carry[3] ));
endmodule

module up_island_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [24:0] A;
   input [24:0] B;
   input CI;
   output [24:0] SUM;
   output CO;

   // Internal wires
   wire \carry[23] ;
   wire \carry[22] ;
   wire \carry[21] ;
   wire \carry[20] ;
   wire \carry[19] ;
   wire \carry[18] ;
   wire \carry[17] ;
   wire \carry[16] ;
   wire \carry[14] ;
   wire \carry[13] ;
   wire \carry[12] ;
   wire \carry[11] ;
   wire \carry[9] ;
   wire \carry[8] ;
   wire \carry[7] ;
   wire \carry[6] ;
   wire \carry[5] ;
   wire \carry[4] ;
   wire \carry[3] ;
   wire \carry[2] ;
   wire \carry[1] ;
   wire n1;
   wire n2;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;

   FA_X1 U1_23 (.S(SUM[23]), 
	.CI(\carry[23] ), 
	.B(B[23]), 
	.A(A[23]));
   FA_X1 U1_19 (.S(SUM[19]), 
	.CO(\carry[20] ), 
	.CI(\carry[19] ), 
	.B(B[19]), 
	.A(A[19]));
   FA_X1 U1_18 (.S(SUM[18]), 
	.CO(\carry[19] ), 
	.CI(\carry[18] ), 
	.B(B[18]), 
	.A(A[18]));
   FA_X1 U1_17 (.S(SUM[17]), 
	.CO(\carry[18] ), 
	.CI(\carry[17] ), 
	.B(B[17]), 
	.A(A[17]));
   FA_X1 U1_16 (.S(SUM[16]), 
	.CO(\carry[17] ), 
	.CI(\carry[16] ), 
	.B(B[16]), 
	.A(A[16]));
   FA_X1 U1_13 (.S(SUM[13]), 
	.CO(\carry[14] ), 
	.CI(\carry[13] ), 
	.B(B[13]), 
	.A(A[13]));
   FA_X1 U1_12 (.S(SUM[12]), 
	.CO(\carry[13] ), 
	.CI(\carry[12] ), 
	.B(B[12]), 
	.A(A[12]));
   FA_X1 U1_11 (.S(SUM[11]), 
	.CO(\carry[12] ), 
	.CI(\carry[11] ), 
	.B(B[11]), 
	.A(A[11]));
   FA_X1 U1_8 (.S(SUM[8]), 
	.CO(\carry[9] ), 
	.CI(\carry[8] ), 
	.B(B[8]), 
	.A(A[8]));
   FA_X1 U1_7 (.S(SUM[7]), 
	.CO(\carry[8] ), 
	.CI(\carry[7] ), 
	.B(B[7]), 
	.A(A[7]));
   FA_X1 U1_6 (.S(SUM[6]), 
	.CO(\carry[7] ), 
	.CI(\carry[6] ), 
	.B(B[6]), 
	.A(A[6]));
   FA_X1 U1_5 (.S(SUM[5]), 
	.CO(\carry[6] ), 
	.CI(\carry[5] ), 
	.B(B[5]), 
	.A(A[5]));
   FA_X1 U1_4 (.S(SUM[4]), 
	.CO(\carry[5] ), 
	.CI(\carry[4] ), 
	.B(B[4]), 
	.A(A[4]));
   FA_X1 U1_3 (.S(SUM[3]), 
	.CO(\carry[4] ), 
	.CI(\carry[3] ), 
	.B(B[3]), 
	.A(A[3]));
   NAND3_X1 U1 (.ZN(n1), 
	.A3(n20), 
	.A2(n19), 
	.A1(n18));
   NAND3_X1 U2 (.ZN(n2), 
	.A3(n28), 
	.A2(n27), 
	.A1(n26));
   XOR2_X1 U5 (.Z(n4), 
	.B(B[20]), 
	.A(A[20]));
   XOR2_X1 U6 (.Z(SUM[20]), 
	.B(\carry[20] ), 
	.A(n4));
   NAND2_X1 U7 (.ZN(n5), 
	.A2(B[20]), 
	.A1(A[20]));
   NAND2_X1 U8 (.ZN(n6), 
	.A2(\carry[20] ), 
	.A1(A[20]));
   NAND2_X1 U9 (.ZN(n7), 
	.A2(\carry[20] ), 
	.A1(B[20]));
   NAND3_X1 U10 (.ZN(\carry[21] ), 
	.A3(n7), 
	.A2(n6), 
	.A1(n5));
   XOR2_X1 U11 (.Z(n8), 
	.B(B[21]), 
	.A(A[21]));
   XOR2_X1 U12 (.Z(SUM[21]), 
	.B(\carry[21] ), 
	.A(n8));
   NAND2_X1 U13 (.ZN(n9), 
	.A2(B[21]), 
	.A1(A[21]));
   NAND2_X1 U14 (.ZN(n10), 
	.A2(\carry[21] ), 
	.A1(A[21]));
   NAND2_X1 U15 (.ZN(n11), 
	.A2(\carry[21] ), 
	.A1(B[21]));
   NAND3_X1 U16 (.ZN(\carry[22] ), 
	.A3(n11), 
	.A2(n10), 
	.A1(n9));
   XOR2_X1 U19 (.Z(n13), 
	.B(A[22]), 
	.A(B[22]));
   XOR2_X1 U20 (.Z(SUM[22]), 
	.B(n13), 
	.A(\carry[22] ));
   NAND2_X1 U21 (.ZN(n14), 
	.A2(B[22]), 
	.A1(\carry[22] ));
   NAND2_X1 U22 (.ZN(n15), 
	.A2(A[22]), 
	.A1(\carry[22] ));
   NAND2_X1 U23 (.ZN(n16), 
	.A2(A[22]), 
	.A1(B[22]));
   NAND3_X1 U24 (.ZN(\carry[23] ), 
	.A3(n15), 
	.A2(n16), 
	.A1(n14));
   XOR2_X1 U25 (.Z(n17), 
	.B(B[9]), 
	.A(A[9]));
   XOR2_X1 U26 (.Z(SUM[9]), 
	.B(\carry[9] ), 
	.A(n17));
   NAND2_X1 U27 (.ZN(n18), 
	.A2(B[9]), 
	.A1(A[9]));
   NAND2_X1 U28 (.ZN(n19), 
	.A2(\carry[9] ), 
	.A1(A[9]));
   NAND2_X1 U29 (.ZN(n20), 
	.A2(\carry[9] ), 
	.A1(B[9]));
   XOR2_X1 U30 (.Z(n21), 
	.B(B[10]), 
	.A(A[10]));
   XOR2_X1 U31 (.Z(SUM[10]), 
	.B(n1), 
	.A(n21));
   NAND2_X1 U32 (.ZN(n22), 
	.A2(B[10]), 
	.A1(A[10]));
   NAND2_X1 U33 (.ZN(n23), 
	.A2(n1), 
	.A1(A[10]));
   NAND2_X1 U34 (.ZN(n24), 
	.A2(n1), 
	.A1(B[10]));
   NAND3_X1 U35 (.ZN(\carry[11] ), 
	.A3(n24), 
	.A2(n23), 
	.A1(n22));
   AND2_X1 U36 (.ZN(\carry[1] ), 
	.A2(A[0]), 
	.A1(B[0]));
   XOR2_X1 U37 (.Z(n25), 
	.B(B[14]), 
	.A(A[14]));
   XOR2_X1 U38 (.Z(SUM[14]), 
	.B(\carry[14] ), 
	.A(n25));
   NAND2_X1 U39 (.ZN(n26), 
	.A2(B[14]), 
	.A1(A[14]));
   NAND2_X1 U40 (.ZN(n27), 
	.A2(\carry[14] ), 
	.A1(A[14]));
   NAND2_X1 U41 (.ZN(n28), 
	.A2(\carry[14] ), 
	.A1(B[14]));
   XOR2_X1 U42 (.Z(n29), 
	.B(B[15]), 
	.A(A[15]));
   XOR2_X1 U43 (.Z(SUM[15]), 
	.B(n2), 
	.A(n29));
   NAND2_X1 U44 (.ZN(n30), 
	.A2(B[15]), 
	.A1(A[15]));
   NAND2_X1 U45 (.ZN(n31), 
	.A2(n2), 
	.A1(A[15]));
   NAND2_X1 U46 (.ZN(n32), 
	.A2(n2), 
	.A1(B[15]));
   NAND3_X1 U47 (.ZN(\carry[16] ), 
	.A3(n30), 
	.A2(n31), 
	.A1(n32));
   XOR2_X1 U48 (.Z(n33), 
	.B(B[1]), 
	.A(A[1]));
   XOR2_X1 U49 (.Z(SUM[1]), 
	.B(\carry[1] ), 
	.A(n33));
   NAND2_X1 U50 (.ZN(n34), 
	.A2(B[1]), 
	.A1(A[1]));
   NAND2_X1 U51 (.ZN(n35), 
	.A2(\carry[1] ), 
	.A1(A[1]));
   NAND2_X1 U52 (.ZN(n36), 
	.A2(\carry[1] ), 
	.A1(B[1]));
   NAND3_X1 U53 (.ZN(\carry[2] ), 
	.A3(n36), 
	.A2(n35), 
	.A1(n34));
   XOR2_X1 U54 (.Z(n37), 
	.B(B[2]), 
	.A(A[2]));
   XOR2_X1 U55 (.Z(SUM[2]), 
	.B(\carry[2] ), 
	.A(n37));
   NAND2_X1 U56 (.ZN(n38), 
	.A2(B[2]), 
	.A1(A[2]));
   NAND2_X1 U57 (.ZN(n39), 
	.A2(\carry[2] ), 
	.A1(A[2]));
   NAND2_X1 U58 (.ZN(n40), 
	.A2(\carry[2] ), 
	.A1(B[2]));
   NAND3_X1 U59 (.ZN(\carry[3] ), 
	.A3(n40), 
	.A2(n39), 
	.A1(n38));
   XOR2_X1 U60 (.Z(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module up_island_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	FE_PT1_n380, 
	n806, 
	n769, 
	n555, 
	n529, 
	n746, 
	n402, 
	n632, 
	n454, 
	n580, 
	n599, 
	n577, 
	FE_PT1_n213, 
	n615, 
	n552, 
	n424, 
	n794, 
	n772, 
	n723, 
	n700, 
	n946, 
	n635, 
	n861);
   input [64:0] A;
   input [64:0] B;
   input CI;
   output [64:0] SUM;
   output CO;
   input FE_PT1_n380;
   input n806;
   input n769;
   input n555;
   input n529;
   input n746;
   input n402;
   input n632;
   input n454;
   input n580;
   input n599;
   input n577;
   input FE_PT1_n213;
   input n615;
   input n552;
   input n424;
   input n794;
   input n772;
   input n723;
   input n700;
   input n946;
   input n635;
   input n861;

   // Internal wires
   wire \carry[58] ;
   wire \carry[47] ;
   wire \carry[46] ;
   wire \carry[45] ;
   wire \carry[29] ;
   wire \carry[20] ;
   wire \carry[19] ;
   wire \carry[15] ;
   wire \carry[6] ;
   wire \carry[5] ;
   wire \carry[1] ;
   wire net55603;
   wire net55599;
   wire net55595;
   wire net55592;
   wire net55587;
   wire net55583;
   wire net55579;
   wire net55571;
   wire net55691;
   wire net55683;
   wire net55682;
   wire net55681;
   wire net55672;
   wire net55837;
   wire net55836;
   wire net55830;
   wire net55826;
   wire net55822;
   wire net55819;
   wire net55817;
   wire net55816;
   wire net55812;
   wire net55808;
   wire net55927;
   wire net55925;
   wire net55923;
   wire net55976;
   wire net55967;
   wire net55964;
   wire net56025;
   wire net56022;
   wire net56020;
   wire net56060;
   wire net56056;
   wire net56052;
   wire net56048;
   wire net56044;
   wire net56040;
   wire net56036;
   wire net56158;
   wire net56154;
   wire net56150;
   wire net56140;
   wire net56227;
   wire net56226;
   wire net56225;
   wire net56313;
   wire net56309;
   wire net56341;
   wire net56336;
   wire net56332;
   wire net56368;
   wire net56437;
   wire net56435;
   wire net56433;
   wire net56427;
   wire net56471;
   wire net56477;
   wire net56476;
   wire net56540;
   wire net56545;
   wire net56549;
   wire net56561;
   wire net56571;
   wire net56562;
   wire net56598;
   wire net56630;
   wire net56628;
   wire net56651;
   wire net56650;
   wire net56649;
   wire net56639;
   wire net56739;
   wire net56755;
   wire net56753;
   wire net56808;
   wire net56856;
   wire net56887;
   wire net56901;
   wire net57006;
   wire net57011;
   wire net57022;
   wire net57069;
   wire net57089;
   wire net57091;
   wire net58078;
   wire net58056;
   wire net58054;
   wire net58040;
   wire net58037;
   wire net58121;
   wire net58242;
   wire net58243;
   wire net58244;
   wire net58238;
   wire net58236;
   wire net58228;
   wire net58227;
   wire net58226;
   wire net58222;
   wire net58210;
   wire net58282;
   wire net58315;
   wire net58323;
   wire net58329;
   wire net58422;
   wire net58404;
   wire net58399;
   wire net58389;
   wire net58447;
   wire net59519;
   wire net59517;
   wire net60649;
   wire net60647;
   wire net60691;
   wire net60758;
   wire net60821;
   wire net60815;
   wire net60813;
   wire net60809;
   wire net60808;
   wire net60794;
   wire net60770;
   wire net60835;
   wire net60880;
   wire net62145;
   wire net62140;
   wire net62139;
   wire net62132;
   wire net62131;
   wire net62130;
   wire net62129;
   wire net62111;
   wire net62110;
   wire net62177;
   wire net62194;
   wire net62205;
   wire net62338;
   wire net62309;
   wire net59538;
   wire net59537;
   wire net56045;
   wire net64022;
   wire net64020;
   wire net64053;
   wire net65126;
   wire net65225;
   wire net65221;
   wire net65201;
   wire net65199;
   wire net65196;
   wire net65188;
   wire net65160;
   wire net65159;
   wire net65153;
   wire net65144;
   wire net65272;
   wire net65290;
   wire net65309;
   wire net65321;
   wire net65638;
   wire net65704;
   wire net65683;
   wire net67391;
   wire net67389;
   wire net67385;
   wire net67373;
   wire net67368;
   wire net67360;
   wire net67359;
   wire net67357;
   wire net67355;
   wire net67429;
   wire net67433;
   wire net67466;
   wire net60799;
   wire net69139;
   wire net69132;
   wire net69126;
   wire net69124;
   wire net69119;
   wire net69117;
   wire net69094;
   wire net69089;
   wire net69188;
   wire net69203;
   wire net70500;
   wire net70495;
   wire net70488;
   wire net70487;
   wire net70483;
   wire net70482;
   wire net70474;
   wire net70465;
   wire net70464;
   wire net70460;
   wire net70456;
   wire net70443;
   wire net70524;
   wire net70527;
   wire net72087;
   wire net72085;
   wire net65288;
   wire net65181;
   wire net73498;
   wire net73494;
   wire net73492;
   wire net73491;
   wire net73490;
   wire net73489;
   wire net73488;
   wire net73487;
   wire net73473;
   wire net73472;
   wire net73468;
   wire net73518;
   wire net73562;
   wire net73570;
   wire net73589;
   wire net73634;
   wire net73660;
   wire net73675;
   wire net65183;
   wire net65687;
   wire net65686;
   wire net65680;
   wire net65675;
   wire net57080;
   wire net56371;
   wire net56370;
   wire net75678;
   wire net75759;
   wire net75757;
   wire net75743;
   wire net75725;
   wire net75723;
   wire net75720;
   wire net75699;
   wire net75831;
   wire net56859;
   wire net77785;
   wire net77768;
   wire net77766;
   wire net77765;
   wire net77818;
   wire net77817;
   wire net77826;
   wire net56041;
   wire net58038;
   wire net56817;
   wire net56144;
   wire net79856;
   wire net79855;
   wire net79851;
   wire net79849;
   wire net79844;
   wire net79832;
   wire net79904;
   wire net56333;
   wire net73564;
   wire net65215;
   wire net64058;
   wire \carry[39] ;
   wire net67379;
   wire \carry[28] ;
   wire net82430;
   wire net82429;
   wire net82427;
   wire net82423;
   wire net82419;
   wire net82413;
   wire net82412;
   wire net82405;
   wire net82402;
   wire net82394;
   wire net82391;
   wire net82387;
   wire net82385;
   wire net82384;
   wire net82383;
   wire net82381;
   wire net82377;
   wire net82373;
   wire net82369;
   wire net82365;
   wire net82355;
   wire net82338;
   wire net82333;
   wire net82512;
   wire net82511;
   wire net82516;
   wire net82542;
   wire net84135;
   wire net84131;
   wire net84129;
   wire net84122;
   wire net84105;
   wire net84099;
   wire net73663;
   wire net73561;
   wire net73557;
   wire net73554;
   wire net65191;
   wire net64019;
   wire net64012;
   wire net57019;
   wire net62344;
   wire net62332;
   wire net62307;
   wire net56569;
   wire net56054;
   wire net65709;
   wire net65697;
   wire net65693;
   wire net65691;
   wire net65679;
   wire net65678;
   wire net65677;
   wire net65671;
   wire net65659;
   wire net65658;
   wire \carry[32] ;
   wire net58409;
   wire net58206;
   wire net58069;
   wire net58061;
   wire net58055;
   wire net84167;
   wire net75846;
   wire net82409;
   wire net82378;
   wire net73517;
   wire net58450;
   wire net58449;
   wire net58424;
   wire net58326;
   wire net58320;
   wire net58289;
   wire net58064;
   wire net58063;
   wire net58060;
   wire net58057;
   wire net56855;
   wire net56142;
   wire \carry[53] ;
   wire net70458;
   wire net69072;
   wire net67456;
   wire net67421;
   wire net55937;
   wire net67465;
   wire net67462;
   wire net56888;
   wire \carry[18] ;
   wire net82523;
   wire net82375;
   wire net70489;
   wire net69130;
   wire net69110;
   wire net84123;
   wire net84111;
   wire net75750;
   wire net75745;
   wire net75736;
   wire net75726;
   wire net75707;
   wire net55680;
   wire net58440;
   wire net58419;
   wire net58393;
   wire net58384;
   wire net58327;
   wire net65682;
   wire net59514;
   wire \carry[3] ;
   wire net79932;
   wire net79908;
   wire net75853;
   wire net60817;
   wire net60810;
   wire net60805;
   wire net60798;
   wire net60797;
   wire net60779;
   wire net60768;
   wire net57039;
   wire net55833;
   wire net87602;
   wire net87601;
   wire net87597;
   wire net87578;
   wire net87623;
   wire net73567;
   wire net73556;
   wire net65251;
   wire net65202;
   wire net65200;
   wire net65197;
   wire net65184;
   wire net75735;
   wire net75731;
   wire net62181;
   wire \carry[43] ;
   wire n2;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n19;
   wire n20;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n39;
   wire n40;
   wire n41;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n56;
   wire n57;
   wire n58;
   wire n60;
   wire n61;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n82;
   wire n83;
   wire n84;
   wire n86;
   wire n87;
   wire n88;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n111;
   wire n112;
   wire n114;
   wire n115;
   wire n116;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n153;
   wire n154;
   wire n155;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n230;
   wire n231;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n253;
   wire n254;
   wire n255;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n273;
   wire n274;
   wire n276;
   wire n277;
   wire n278;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n295;
   wire n296;
   wire n297;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n304;
   wire n305;
   wire n307;
   wire n308;
   wire n309;
   wire n311;
   wire n312;
   wire n313;
   wire n316;
   wire n319;
   wire n321;
   wire n322;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n337;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n352;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n359;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n372;
   wire n374;
   wire n376;
   wire n377;
   wire n378;
   wire n380;
   wire n382;
   wire n383;
   wire n384;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n391;
   wire n392;
   wire n395;

   NOR2_X1 net58124 (.ZN(net58315), 
	.A2(n402), 
	.A1(net58404));
   NAND3_X1 net57010 (.ZN(net56158), 
	.A3(n297), 
	.A2(net62111), 
	.A1(net62110));
   NAND2_X1 net62274 (.ZN(net60808), 
	.A2(net60815), 
	.A1(net62309));
   NAND2_X1 net62276 (.ZN(net60809), 
	.A2(net60813), 
	.A1(B[24]));
   NAND2_X1 net65122 (.ZN(net55817), 
	.A2(net65201), 
	.A1(net65144));
   NAND2_X1 syn338 (.ZN(net69094), 
	.A2(B[12]), 
	.A1(net70464));
   NAND3_X1 net56885 (.ZN(net56020), 
	.A3(net69094), 
	.A2(net55925), 
	.A1(net69089));
   NAND2_X1 net70438 (.ZN(net69132), 
	.A2(net70443), 
	.A1(n270));
   INV_X1 syn301 (.ZN(net56753), 
	.A(n265));
   INV_X1 syn271 (.ZN(net73490), 
	.A(net73468));
   INV_X1 syn371 (.ZN(net56336), 
	.A(net75757));
   NAND2_X1 net58346 (.ZN(net56041), 
	.A2(A[50]), 
	.A1(B[50]));
   NAND2_X1 syn194 (.ZN(net79844), 
	.A2(B[39]), 
	.A1(A[39]));
   INV_X1 syn454 (.ZN(n222), 
	.A(n223));
   NAND3_X1 net56021 (.ZN(net55976), 
	.A3(net67357), 
	.A2(net67391), 
	.A1(net67355));
   MUX2_X1 syn755 (.Z(n181), 
	.S(n200), 
	.B(n203), 
	.A(net82338));
   NAND2_X1 syn753 (.ZN(n203), 
	.A2(n580), 
	.A1(A[11]));
   XNOR2_X1 syn751 (.ZN(n201), 
	.B(n580), 
	.A(n199));
   INV_X1 syn750 (.ZN(net55967), 
	.A(n202));
   XNOR2_X1 syn749 (.ZN(n202), 
	.B(A[10]), 
	.A(B[10]));
   NAND2_X1 syn747 (.ZN(n182), 
	.A2(net82365), 
	.A1(n201));
   INV_X1 syn721 (.ZN(net82427), 
	.A(net82383));
   NAND2_X1 syn717 (.ZN(n192), 
	.A2(net82384), 
	.A1(net82381));
   INV_X1 syn704 (.ZN(net82387), 
	.A(net82381));
   NAND2_X1 syn687 (.ZN(n195), 
	.A2(net70500), 
	.A1(net82419));
   NAND2_X1 syn649 (.ZN(net82377), 
	.A2(net82365), 
	.A1(n580));
   INV_X1 syn643 (.ZN(net82419), 
	.A(net82338));
   INV_X1 syn640 (.ZN(n200), 
	.A(n199));
   OAI21_X1 syn638 (.ZN(n199), 
	.B2(n599), 
	.B1(net82413), 
	.A(n198));
   NAND2_X1 syn636 (.ZN(n198), 
	.A2(net77826), 
	.A1(A[10]));
   INV_X1 syn633 (.ZN(net82413), 
	.A(net82412));
   AND3_X1 syn502 (.ZN(n185), 
	.A3(n194), 
	.A2(n195), 
	.A1(n196));
   NAND2_X1 syn245 (.ZN(net82383), 
	.A2(net70500), 
	.A1(net82384));
   INV_X1 syn25 (.ZN(net82355), 
	.A(net56025));
   NAND2_X1 net82294 (.ZN(SUM[11]), 
	.A2(n182), 
	.A1(n181));
   NAND3_X1 net75835 (.ZN(net75831), 
	.A3(net62181), 
	.A2(net84167), 
	.A1(net56333));
   NAND2_X1 net84066 (.ZN(net75743), 
	.A2(net84105), 
	.A1(n162));
   NAND2_X1 net84042 (.ZN(net56476), 
	.A2(n161), 
	.A1(net62194));
   NAND2_X1 net84068 (.ZN(net75757), 
	.A2(n160), 
	.A1(net75725));
   AOI21_X1 net65125 (.ZN(net65126), 
	.B2(net65160), 
	.B1(net65159), 
	.A(n153));
   NAND2_X1 net62260 (.ZN(net60647), 
	.A2(net60794), 
	.A1(net60770));
   NAND2_X1 syn40 (.ZN(net65679), 
	.A2(net65671), 
	.A1(n946));
   NAND2_X1 net58373 (.ZN(net58236), 
	.A2(net58399), 
	.A1(net56041));
   NAND3_X1 net56627 (.ZN(net57006), 
	.A3(net58078), 
	.A2(net56041), 
	.A1(net58228));
   OAI21_X1 net73459 (.ZN(net72087), 
	.B2(B[7]), 
	.B1(A[7]), 
	.A(net73468));
   AOI21_X1 net70423 (.ZN(net56808), 
	.B2(net69094), 
	.B1(net70456), 
	.A(net70458));
   NAND2_X1 syn745 (.ZN(net82391), 
	.A2(net82423), 
	.A1(net82375));
   NOR2_X1 syn498 (.ZN(net82394), 
	.A2(net82369), 
	.A1(n105));
   NOR2_X1 syn520 (.ZN(net82402), 
	.A2(n105), 
	.A1(net82373));
   NAND2_X1 net70430 (.ZN(net69110), 
	.A2(net70443), 
	.A1(B[14]));
   NAND2_X1 syn515 (.ZN(n108), 
	.A2(net70489), 
	.A1(net82384));
   NAND2_X1 net55972 (.ZN(net82338), 
	.A2(A[11]), 
	.A1(B[11]));
   NAND3_X1 syn632 (.ZN(net82412), 
	.A3(net82523), 
	.A2(net82387), 
	.A1(n49));
   NAND3_X1 syn737 (.ZN(net82430), 
	.A3(net82387), 
	.A2(net82523), 
	.A1(net73517));
   NAND3_X1 syn739 (.ZN(net82405), 
	.A3(n111), 
	.A2(net73517), 
	.A1(net82523));
   INV_X1 syn653 (.ZN(n111), 
	.A(net82375));
   NOR2_X1 syn510 (.ZN(n107), 
	.A2(n105), 
	.A1(n104));
   NAND2_X1 net84036 (.ZN(\carry[45] ), 
	.A2(net84111), 
	.A1(net75726));
   NAND2_X1 net84060 (.ZN(net75725), 
	.A2(n577), 
	.A1(n103));
   NOR2_X1 syn164 (.ZN(net84123), 
	.A2(net75745), 
	.A1(A[43]));
   INV_X1 net84067 (.ZN(net75745), 
	.A(net75726));
   NAND3_X1 net58376 (.ZN(net58242), 
	.A3(net58389), 
	.A2(A[49]), 
	.A1(B[49]));
   NAND2_X1 net58374 (.ZN(net58238), 
	.A2(net58393), 
	.A1(net58384));
   NAND3_X1 net65644 (.ZN(net56628), 
	.A3(net65697), 
	.A2(net65704), 
	.A1(net59514));
   OAI21_X1 net60751 (.ZN(net56471), 
	.B2(net60805), 
	.B1(net75853), 
	.A(net60768));
   INV_X1 net62278 (.ZN(net60810), 
	.A(net60770));
   AND2_X1 net60757 (.ZN(net60758), 
	.A2(n73), 
	.A1(net69203));
   NAND2_X1 net62247 (.ZN(net55833), 
	.A2(A[24]), 
	.A1(B[24]));
   NOR2_X1 net62259 (.ZN(net57039), 
	.A2(net60779), 
	.A1(n75));
   NAND2_X1 syn223 (.ZN(net87578), 
	.A2(net87601), 
	.A1(net87602));
   INV_X1 net65132 (.ZN(net64012), 
	.A(A[37]));
   OAI21_X1 net65134 (.ZN(net64020), 
	.B2(B[37]), 
	.B1(A[37]), 
	.A(net65153));
   NAND3_X1 net84034 (.ZN(\carry[43] ), 
	.A3(net56333), 
	.A2(net84167), 
	.A1(net62181));
   INV_X1 net84062 (.ZN(net75731), 
	.A(net75723));
   INV_X1 syn283 (.ZN(n22), 
	.A(n35));
   NAND2_X1 syn282 (.ZN(n35), 
	.A2(n33), 
	.A1(n34));
   NAND2_X1 syn274 (.ZN(n34), 
	.A2(A[61]), 
	.A1(net87578));
   NAND2_X1 syn272 (.ZN(n33), 
	.A2(B[61]), 
	.A1(net87578));
   NAND2_X1 syn263 (.ZN(n26), 
	.A2(B[62]), 
	.A1(A[62]));
   NAND3_X1 syn261 (.ZN(n31), 
	.A3(net56649), 
	.A2(n26), 
	.A1(n27));
   NAND3_X1 syn234 (.ZN(n28), 
	.A3(net56540), 
	.A2(A[62]), 
	.A1(B[62]));
   OAI21_X1 syn197 (.ZN(n17), 
	.B2(n20), 
	.B1(n19), 
	.A(n28));
   NOR2_X1 syn190 (.ZN(n27), 
	.A2(B[62]), 
	.A1(A[62]));
   NAND3_X1 syn189 (.ZN(n25), 
	.A3(net56649), 
	.A2(n26), 
	.A1(n20));
   XNOR2_X1 syn182 (.ZN(net56477), 
	.B(n861), 
	.A(A[62]));
   XNOR2_X1 syn172 (.ZN(net87597), 
	.B(A[61]), 
	.A(B[61]));
   NOR2_X1 syn146 (.ZN(n23), 
	.A2(A[61]), 
	.A1(B[61]));
   NAND3_X1 syn141 (.ZN(net87623), 
	.A3(net56227), 
	.A2(net56225), 
	.A1(net56226));
   NAND2_X1 syn69 (.ZN(n20), 
	.A2(A[61]), 
	.A1(B[61]));
   INV_X1 syn46 (.ZN(n19), 
	.A(net87578));
   NOR2_X1 net88854 (.ZN(net56650), 
	.A2(n17), 
	.A1(n16));
   NAND2_X1 net88860 (.ZN(net87602), 
	.A2(B[62]), 
	.A1(net56540));
   NAND2_X1 net88859 (.ZN(net87601), 
	.A2(A[62]), 
	.A1(net56540));
   INV_X1 U1 (.ZN(net73561), 
	.A(net62131));
   INV_X1 U3 (.ZN(n58), 
	.A(n359));
   NAND2_X1 U5 (.ZN(n180), 
	.A2(n2), 
	.A1(net82430));
   AND2_X1 U6 (.ZN(n2), 
	.A2(net70488), 
	.A1(net82384));
   NAND2_X1 U8 (.ZN(n4), 
	.A2(B[17]), 
	.A1(n121));
   AND3_X1 U10 (.ZN(n5), 
	.A3(net73561), 
	.A2(net62139), 
	.A1(net73562));
   NAND3_X1 U11 (.ZN(n6), 
	.A3(n245), 
	.A2(n54), 
	.A1(n8));
   NAND3_X1 U12 (.ZN(n116), 
	.A3(n115), 
	.A2(n114), 
	.A1(net56888));
   NAND3_X1 U13 (.ZN(\carry[46] ), 
	.A3(net55682), 
	.A2(net55681), 
	.A1(net55680));
   NOR2_X1 U14 (.ZN(n7), 
	.A2(net56435), 
	.A1(net65680));
   NAND2_X1 U15 (.ZN(n8), 
	.A2(B[47]), 
	.A1(n61));
   NAND3_X1 U16 (.ZN(n9), 
	.A3(n388), 
	.A2(n389), 
	.A1(n319));
   NAND2_X1 U17 (.ZN(n389), 
	.A2(A[56]), 
	.A1(n321));
   NAND3_X1 U18 (.ZN(n337), 
	.A3(n368), 
	.A2(n369), 
	.A1(net57091));
   NAND3_X1 U20 (.ZN(n10), 
	.A3(n112), 
	.A2(n4), 
	.A1(net67462));
   NOR2_X1 U21 (.ZN(net65290), 
	.A2(net65309), 
	.A1(n41));
   NOR2_X1 U25 (.ZN(n24), 
	.A2(n23), 
	.A1(n36));
   NAND2_X1 U26 (.ZN(n11), 
	.A2(A[1]), 
	.A1(\carry[1] ));
   NAND3_X1 U28 (.ZN(n12), 
	.A3(n88), 
	.A2(n90), 
	.A1(n86));
   NAND2_X1 U29 (.ZN(n88), 
	.A2(n93), 
	.A1(n94));
   NAND2_X1 U30 (.ZN(net73517), 
	.A2(n145), 
	.A1(n146));
   NOR2_X1 U31 (.ZN(n16), 
	.A2(n22), 
	.A1(n37));
   NAND2_X1 U33 (.ZN(n14), 
	.A2(B[46]), 
	.A1(\carry[46] ));
   NAND3_X1 U34 (.ZN(n15), 
	.A3(n354), 
	.A2(n328), 
	.A1(net56549));
   AND3_X1 U35 (.ZN(n36), 
	.A3(net56225), 
	.A2(net56227), 
	.A1(net56226));
   OAI21_X1 U36 (.ZN(n32), 
	.B2(n36), 
	.B1(n23), 
	.A(n20));
   XNOR2_X1 U37 (.ZN(SUM[62]), 
	.B(net56598), 
	.A(n32));
   OAI21_X1 U38 (.ZN(n30), 
	.B2(n25), 
	.B1(n24), 
	.A(n31));
   INV_X1 U39 (.ZN(net56651), 
	.A(n30));
   INV_X1 U40 (.ZN(n37), 
	.A(net87623));
   NOR2_X1 U41 (.ZN(net75735), 
	.A2(n39), 
	.A1(n40));
   AOI21_X1 U42 (.ZN(net55680), 
	.B2(net75736), 
	.B1(net75735), 
	.A(net75707));
   NOR2_X1 U43 (.ZN(n40), 
	.A2(B[43]), 
	.A1(\carry[43] ));
   NAND2_X1 U44 (.ZN(n39), 
	.A2(B[45]), 
	.A1(net75731));
   NAND2_X1 U46 (.ZN(net84111), 
	.A2(net75731), 
	.A1(net84135));
   NAND2_X1 U48 (.ZN(net62181), 
	.A2(B[42]), 
	.A1(net79932));
   NAND2_X1 U49 (.ZN(net84122), 
	.A2(net75726), 
	.A1(net75723));
   NAND2_X1 U50 (.ZN(net84167), 
	.A2(A[42]), 
	.A1(net82512));
   OAI21_X1 U52 (.ZN(n41), 
	.B2(n43), 
	.B1(n46), 
	.A(n44));
   NAND2_X1 U53 (.ZN(n44), 
	.A2(B[38]), 
	.A1(net65202));
   INV_X1 U54 (.ZN(net65202), 
	.A(net65153));
   NAND2_X1 U55 (.ZN(n46), 
	.A2(net65196), 
	.A1(net65197));
   NAND2_X1 U56 (.ZN(n43), 
	.A2(net64019), 
	.A1(B[38]));
   INV_X1 U57 (.ZN(net65225), 
	.A(n43));
   NAND2_X1 U58 (.ZN(net65153), 
	.A2(A[37]), 
	.A1(B[37]));
   NAND2_X1 U59 (.ZN(net65197), 
	.A2(n45), 
	.A1(n5));
   INV_X1 U61 (.ZN(n45), 
	.A(net65251));
   AND2_X1 U62 (.ZN(net73567), 
	.A2(net65153), 
	.A1(n45));
   AND2_X1 U63 (.ZN(net73556), 
	.A2(net73557), 
	.A1(n45));
   NAND2_X1 U64 (.ZN(net65251), 
	.A2(net65184), 
	.A1(net65201));
   INV_X1 U65 (.ZN(net65184), 
	.A(A[36]));
   AOI21_X1 U66 (.ZN(net65196), 
	.B2(net65201), 
	.B1(net65200), 
	.A(n723));
   NOR2_X1 U68 (.ZN(net65200), 
	.A2(net65183), 
	.A1(A[36]));
   INV_X1 U69 (.ZN(net65215), 
	.A(net64019));
   NAND2_X1 U70 (.ZN(net73554), 
	.A2(net73556), 
	.A1(n5));
   NAND2_X1 U71 (.ZN(net73564), 
	.A2(net73567), 
	.A1(n5));
   XNOR2_X1 U72 (.ZN(net64022), 
	.B(A[36]), 
	.A(B[36]));
   NAND2_X1 U73 (.ZN(net65144), 
	.A2(net65288), 
	.A1(net65183));
   NAND2_X1 U74 (.ZN(net65191), 
	.A2(net65183), 
	.A1(A[36]));
   NAND2_X1 U75 (.ZN(n47), 
	.A2(net84099), 
	.A1(net75846));
   NOR2_X1 U76 (.ZN(net84099), 
	.A2(B[43]), 
	.A1(net75745));
   OAI21_X1 U77 (.ZN(net60797), 
	.B2(net60805), 
	.B1(net79908), 
	.A(net60817));
   NAND3_X1 U78 (.ZN(n48), 
	.A3(net79844), 
	.A2(n168), 
	.A1(n178));
   AND3_X1 U80 (.ZN(net70460), 
	.A3(n183), 
	.A2(n184), 
	.A1(n185));
   INV_X1 U81 (.ZN(n49), 
	.A(net82542));
   NAND2_X1 U82 (.ZN(n50), 
	.A2(A[48]), 
	.A1(n6));
   NAND2_X1 U83 (.ZN(n51), 
	.A2(net79856), 
	.A1(n48));
   OAI21_X1 U84 (.ZN(n264), 
	.B2(net73489), 
	.B1(net73494), 
	.A(net73468));
   AND2_X1 U85 (.ZN(net79904), 
	.A2(net79849), 
	.A1(n51));
   AND2_X1 U86 (.ZN(n52), 
	.A2(n78), 
	.A1(n77));
   NAND2_X1 U88 (.ZN(n53), 
	.A2(B[53]), 
	.A1(\carry[53] ));
   NAND2_X1 U89 (.ZN(n54), 
	.A2(A[47]), 
	.A1(\carry[47] ));
   NAND2_X1 U91 (.ZN(n56), 
	.A2(A[46]), 
	.A1(n333));
   NAND2_X1 U93 (.ZN(n57), 
	.A2(B[55]), 
	.A1(n171));
   XNOR2_X1 U94 (.ZN(SUM[60]), 
	.B(n350), 
	.A(n58));
   NAND2_X1 U97 (.ZN(n60), 
	.A2(net67360), 
	.A1(net67359));
   NAND3_X1 U98 (.ZN(n61), 
	.A3(n392), 
	.A2(n14), 
	.A1(n56));
   NOR2_X1 U100 (.ZN(n183), 
	.A2(n188), 
	.A1(net82385));
   INV_X1 U102 (.ZN(n64), 
	.A(n172));
   NAND2_X1 U103 (.ZN(n65), 
	.A2(net70500), 
	.A1(net82423));
   NAND2_X1 U104 (.ZN(n196), 
	.A2(n66), 
	.A1(net82429));
   INV_X1 U105 (.ZN(n66), 
	.A(n65));
   NAND2_X1 U106 (.ZN(net70500), 
	.A2(net70474), 
	.A1(n555));
   INV_X1 U107 (.ZN(net82423), 
	.A(n105));
   NAND2_X1 U109 (.ZN(n67), 
	.A2(B[48]), 
	.A1(n6));
   NAND2_X1 U110 (.ZN(n68), 
	.A2(B[26]), 
	.A1(n302));
   AOI21_X1 U111 (.ZN(n109), 
	.B2(n107), 
	.B1(net82405), 
	.A(n106));
   XNOR2_X1 U112 (.ZN(SUM[61]), 
	.B(net87597), 
	.A(net87623));
   AND2_X1 U113 (.ZN(n69), 
	.A2(n180), 
	.A1(n197));
   NAND3_X1 U114 (.ZN(n70), 
	.A3(net55833), 
	.A2(n71), 
	.A1(net57039));
   NAND2_X1 U115 (.ZN(net60691), 
	.A2(A[25]), 
	.A1(n70));
   NAND2_X1 U117 (.ZN(n71), 
	.A2(n74), 
	.A1(net60797));
   AND2_X1 U118 (.ZN(n74), 
	.A2(A[24]), 
	.A1(n73));
   INV_X1 U119 (.ZN(net60817), 
	.A(net60798));
   OAI21_X1 U120 (.ZN(net69203), 
	.B2(net60805), 
	.B1(net75853), 
	.A(net60817));
   NAND2_X1 U123 (.ZN(net60798), 
	.A2(net60794), 
	.A1(net60768));
   NOR2_X1 U124 (.ZN(net60805), 
	.A2(B[22]), 
	.A1(A[22]));
   NAND2_X1 U125 (.ZN(net60779), 
	.A2(net60809), 
	.A1(net60808));
   NOR2_X1 U126 (.ZN(n75), 
	.A2(net62307), 
	.A1(net75853));
   AND3_X1 U127 (.ZN(net75853), 
	.A3(net62332), 
	.A2(net56054), 
	.A1(net62344));
   NAND3_X1 U128 (.ZN(net82511), 
	.A3(net55833), 
	.A2(net65321), 
	.A1(net82516));
   NAND3_X1 U129 (.ZN(net60880), 
	.A3(net55833), 
	.A2(net65321), 
	.A1(net57039));
   NAND2_X1 U131 (.ZN(n73), 
	.A2(net60794), 
	.A1(net60810));
   XNOR2_X1 U133 (.ZN(net62338), 
	.B(A[24]), 
	.A(B[24]));
   AND3_X1 U134 (.ZN(net79908), 
	.A3(net62332), 
	.A2(net62344), 
	.A1(net56054));
   NOR2_X1 U135 (.ZN(net60799), 
	.A2(net62307), 
	.A1(net79908));
   NAND2_X1 U136 (.ZN(net60768), 
	.A2(B[22]), 
	.A1(A[22]));
   INV_X1 U137 (.ZN(net60815), 
	.A(net60768));
   NAND3_X1 U138 (.ZN(net79932), 
	.A3(net56371), 
	.A2(net79904), 
	.A1(n52));
   OR2_X1 U141 (.ZN(n78), 
	.A2(net79832), 
	.A1(n79));
   INV_X1 U142 (.ZN(n79), 
	.A(A[41]));
   NAND2_X1 U143 (.ZN(n77), 
	.A2(n80), 
	.A1(n48));
   AND2_X1 U144 (.ZN(n80), 
	.A2(A[41]), 
	.A1(net79855));
   NAND2_X1 U146 (.ZN(net56371), 
	.A2(A[41]), 
	.A1(B[41]));
   NAND2_X1 U148 (.ZN(net56630), 
	.A2(net79832), 
	.A1(n76));
   INV_X1 U149 (.ZN(net79851), 
	.A(net79832));
   NAND2_X1 U150 (.ZN(n76), 
	.A2(net79855), 
	.A1(n48));
   NAND2_X1 U152 (.ZN(\carry[3] ), 
	.A2(n83), 
	.A1(n82));
   NAND2_X1 U153 (.ZN(net62205), 
	.A2(B[3]), 
	.A1(\carry[3] ));
   NAND2_X1 U156 (.ZN(n83), 
	.A2(B[2]), 
	.A1(n92));
   AND2_X1 U158 (.ZN(net77765), 
	.A2(B[2]), 
	.A1(A[3]));
   XNOR2_X1 U159 (.ZN(net77785), 
	.B(A[2]), 
	.A(B[2]));
   NAND3_X1 U161 (.ZN(n92), 
	.A3(n91), 
	.A2(n11), 
	.A1(n90));
   NAND2_X1 U162 (.ZN(n82), 
	.A2(A[2]), 
	.A1(n87));
   NAND2_X1 U165 (.ZN(n90), 
	.A2(B[1]), 
	.A1(net57022));
   NAND2_X1 U168 (.ZN(n91), 
	.A2(A[1]), 
	.A1(B[1]));
   NAND2_X1 U173 (.ZN(n86), 
	.A2(A[1]), 
	.A1(net57022));
   NAND3_X1 U174 (.ZN(n87), 
	.A3(n86), 
	.A2(n90), 
	.A1(n88));
   NAND2_X1 U175 (.ZN(net77768), 
	.A2(net77766), 
	.A1(n12));
   NAND2_X1 U176 (.ZN(n93), 
	.A2(n84), 
	.A1(n772));
   INV_X1 U177 (.ZN(n84), 
	.A(A[1]));
   NAND2_X1 U178 (.ZN(n94), 
	.A2(n794), 
	.A1(n772));
   NOR2_X1 U180 (.ZN(n100), 
	.A2(net65682), 
	.A1(n101));
   AOI21_X1 U181 (.ZN(\carry[32] ), 
	.B2(net65697), 
	.B1(n100), 
	.A(net65659));
   AND2_X1 U182 (.ZN(n101), 
	.A2(A[30]), 
	.A1(net57011));
   NAND2_X1 U185 (.ZN(net65682), 
	.A2(net59514), 
	.A1(net65677));
   NOR2_X1 U186 (.ZN(net65658), 
	.A2(n101), 
	.A1(net65682));
   NAND2_X1 U187 (.ZN(net56435), 
	.A2(A[30]), 
	.A1(net57011));
   XNOR2_X1 U188 (.ZN(net59517), 
	.B(B[30]), 
	.A(A[30]));
   NAND2_X1 U189 (.ZN(net59514), 
	.A2(B[30]), 
	.A1(A[30]));
   NAND2_X1 U190 (.ZN(net65693), 
	.A2(net65677), 
	.A1(net65691));
   NOR2_X1 U191 (.ZN(net65678), 
	.A2(net65677), 
	.A1(net65675));
   NOR2_X1 U192 (.ZN(net65683), 
	.A2(net59514), 
	.A1(net65680));
   NAND2_X1 U193 (.ZN(net58327), 
	.A2(net58393), 
	.A1(n102));
   NAND2_X1 U194 (.ZN(net58057), 
	.A2(net58326), 
	.A1(net58327));
   NAND2_X1 U195 (.ZN(net58449), 
	.A2(net58409), 
	.A1(net58327));
   NAND2_X1 U197 (.ZN(n102), 
	.A2(net58384), 
	.A1(net58440));
   NAND2_X1 U198 (.ZN(net58393), 
	.A2(B[49]), 
	.A1(A[49]));
   NAND3_X1 U201 (.ZN(net58440), 
	.A3(net58226), 
	.A2(n50), 
	.A1(net58227));
   NAND2_X1 U203 (.ZN(net58384), 
	.A2(net58419), 
	.A1(n424));
   INV_X1 U204 (.ZN(net58222), 
	.A(net58384));
   INV_X1 U205 (.ZN(net58419), 
	.A(A[49]));
   AND3_X1 U208 (.ZN(net58329), 
	.A3(net58226), 
	.A2(n50), 
	.A1(n67));
   INV_X1 U209 (.ZN(net75707), 
	.A(net75750));
   NAND2_X1 U210 (.ZN(net75750), 
	.A2(B[45]), 
	.A1(net75745));
   NAND2_X1 U211 (.ZN(net75736), 
	.A2(n103), 
	.A1(net75846));
   INV_X1 U212 (.ZN(n103), 
	.A(A[43]));
   NAND3_X1 U213 (.ZN(net84105), 
	.A3(net84131), 
	.A2(n103), 
	.A1(net75726));
   NAND2_X1 U214 (.ZN(net75726), 
	.A2(B[44]), 
	.A1(A[44]));
   NAND2_X1 U215 (.ZN(net84129), 
	.A2(net84123), 
	.A1(net75846));
   INV_X1 U217 (.ZN(net75720), 
	.A(A[44]));
   XNOR2_X1 U218 (.ZN(net75759), 
	.B(B[44]), 
	.A(A[44]));
   OAI21_X1 U220 (.ZN(net82409), 
	.B2(n108), 
	.B1(net82413), 
	.A(n109));
   NOR2_X1 U221 (.ZN(n106), 
	.A2(net82338), 
	.A1(n104));
   INV_X1 U222 (.ZN(n104), 
	.A(net70489));
   NAND2_X1 U223 (.ZN(net82429), 
	.A2(n111), 
	.A1(net73517));
   NOR2_X1 U224 (.ZN(net82385), 
	.A2(net73517), 
	.A1(net82383));
   AND2_X1 U225 (.ZN(net70489), 
	.A2(net69130), 
	.A1(A[12]));
   NAND2_X1 U226 (.ZN(net70527), 
	.A2(net70489), 
	.A1(net70464));
   INV_X1 U227 (.ZN(net69130), 
	.A(net69110));
   NAND2_X1 U228 (.ZN(net69117), 
	.A2(net69130), 
	.A1(net69126));
   AND2_X1 U229 (.ZN(net70488), 
	.A2(B[12]), 
	.A1(net69130));
   NAND2_X1 U230 (.ZN(n105), 
	.A2(A[10]), 
	.A1(net82377));
   AND2_X1 U231 (.ZN(net82523), 
	.A2(n241), 
	.A1(n240));
   NAND2_X1 U233 (.ZN(net82375), 
	.A2(net56025), 
	.A1(net73518));
   NOR2_X1 U234 (.ZN(net82333), 
	.A2(net82375), 
	.A1(net82542));
   NAND2_X1 U235 (.ZN(net57091), 
	.A2(B[19]), 
	.A1(n116));
   NAND2_X1 U238 (.ZN(n114), 
	.A2(A[18]), 
	.A1(\carry[18] ));
   NAND2_X1 U239 (.ZN(net56888), 
	.A2(B[18]), 
	.A1(\carry[18] ));
   NAND2_X1 U240 (.ZN(n115), 
	.A2(A[18]), 
	.A1(B[18]));
   NAND3_X1 U241 (.ZN(\carry[19] ), 
	.A3(n115), 
	.A2(n114), 
	.A1(net67465));
   NAND3_X1 U242 (.ZN(\carry[18] ), 
	.A3(n112), 
	.A2(net67462), 
	.A1(n4));
   NAND2_X1 U244 (.ZN(net67462), 
	.A2(A[17]), 
	.A1(n60));
   NAND2_X1 U246 (.ZN(n121), 
	.A2(net67379), 
	.A1(net67421));
   XOR2_X1 U247 (.Z(net56887), 
	.B(A[18]), 
	.A(B[18]));
   NAND2_X1 U249 (.ZN(net67465), 
	.A2(B[18]), 
	.A1(n10));
   NAND2_X1 U253 (.ZN(n112), 
	.A2(B[17]), 
	.A1(A[17]));
   XOR2_X1 U254 (.Z(net55603), 
	.B(B[17]), 
	.A(A[17]));
   AND2_X1 U255 (.ZN(net67421), 
	.A2(n126), 
	.A1(n127));
   INV_X1 U256 (.ZN(n126), 
	.A(n123));
   AND2_X1 U257 (.ZN(net67359), 
	.A2(n126), 
	.A1(net67385));
   OAI21_X1 U258 (.ZN(n123), 
	.B2(net67355), 
	.B1(n124), 
	.A(n125));
   NAND2_X1 U259 (.ZN(n125), 
	.A2(A[16]), 
	.A1(B[16]));
   INV_X1 U260 (.ZN(n124), 
	.A(net67373));
   NAND2_X1 U261 (.ZN(n127), 
	.A2(n128), 
	.A1(net55937));
   INV_X1 U262 (.ZN(n128), 
	.A(n122));
   NAND2_X1 U263 (.ZN(net67360), 
	.A2(n128), 
	.A1(net67466));
   NAND2_X1 U264 (.ZN(n122), 
	.A2(B[15]), 
	.A1(net67373));
   NAND3_X1 U265 (.ZN(net55937), 
	.A3(net55837), 
	.A2(net69188), 
	.A1(net67456));
   NAND2_X1 U266 (.ZN(net67456), 
	.A2(A[14]), 
	.A1(net69072));
   AOI21_X1 U267 (.ZN(net69072), 
	.B2(n129), 
	.B1(net70460), 
	.A(net70458));
   INV_X1 U268 (.ZN(net70458), 
	.A(net70443));
   INV_X1 U270 (.ZN(n129), 
	.A(net70482));
   NOR2_X1 U271 (.ZN(net70465), 
	.A2(n129), 
	.A1(net70483));
   NAND3_X1 U272 (.ZN(n132), 
	.A3(net56144), 
	.A2(n134), 
	.A1(n53));
   NAND2_X1 U273 (.ZN(net55819), 
	.A2(B[54]), 
	.A1(n132));
   NAND3_X1 U278 (.ZN(\carry[53] ), 
	.A3(net56140), 
	.A2(net58289), 
	.A1(net56855));
   INV_X1 U279 (.ZN(net58289), 
	.A(net58320));
   OAI211_X1 U280 (.ZN(net58320), 
	.C2(net58061), 
	.C1(net58064), 
	.B(net58449), 
	.A(n135));
   NAND2_X1 U281 (.ZN(n135), 
	.A2(net58206), 
	.A1(net58327));
   INV_X1 U282 (.ZN(net58064), 
	.A(net58069));
   OAI211_X1 U283 (.ZN(net58063), 
	.C2(net58061), 
	.C1(net58064), 
	.B(n135), 
	.A(net58449));
   OAI21_X1 U284 (.ZN(net56855), 
	.B2(net58040), 
	.B1(n133), 
	.A(A[52]));
   NAND2_X1 U285 (.ZN(n133), 
	.A2(net58057), 
	.A1(net58060));
   NOR2_X1 U286 (.ZN(net58060), 
	.A2(net58450), 
	.A1(n136));
   INV_X1 U287 (.ZN(net58450), 
	.A(net58242));
   NOR2_X1 U288 (.ZN(n136), 
	.A2(net58329), 
	.A1(net58244));
   INV_X1 U289 (.ZN(net58326), 
	.A(net58424));
   NAND2_X1 U291 (.ZN(net58424), 
	.A2(net58054), 
	.A1(B[50]));
   NAND2_X1 U292 (.ZN(n134), 
	.A2(A[53]), 
	.A1(n131));
   NAND3_X1 U293 (.ZN(n131), 
	.A3(net56140), 
	.A2(n130), 
	.A1(net56142));
   INV_X1 U294 (.ZN(net56142), 
	.A(net58063));
   NAND2_X1 U297 (.ZN(n130), 
	.A2(A[52]), 
	.A1(net56817));
   NAND3_X1 U298 (.ZN(n141), 
	.A3(n138), 
	.A2(n139), 
	.A1(n140));
   NAND2_X1 U299 (.ZN(net56549), 
	.A2(B[58]), 
	.A1(n141));
   NAND2_X1 U302 (.ZN(n140), 
	.A2(B[57]), 
	.A1(n9));
   NAND3_X1 U303 (.ZN(\carry[58] ), 
	.A3(n140), 
	.A2(n138), 
	.A1(n139));
   NAND2_X1 U304 (.ZN(n139), 
	.A2(A[57]), 
	.A1(n9));
   NAND2_X1 U305 (.ZN(n138), 
	.A2(B[57]), 
	.A1(A[57]));
   XOR2_X1 U306 (.Z(net55571), 
	.B(B[57]), 
	.A(A[57]));
   INV_X1 U307 (.ZN(net82542), 
	.A(net73517));
   AND2_X1 U308 (.ZN(n145), 
	.A2(B[9]), 
	.A1(n144));
   NAND3_X1 U309 (.ZN(n146), 
	.A3(net73487), 
	.A2(net73488), 
	.A1(net56755));
   NAND2_X1 U311 (.ZN(n144), 
	.A2(n142), 
	.A1(n143));
   AND2_X1 U312 (.ZN(net77818), 
	.A2(A[9]), 
	.A1(n144));
   NAND2_X1 U313 (.ZN(net73473), 
	.A2(n144), 
	.A1(n146));
   NAND2_X1 U315 (.ZN(n142), 
	.A2(A[7]), 
	.A1(net73491));
   NAND2_X1 U316 (.ZN(n143), 
	.A2(B[7]), 
	.A1(net73491));
   NAND2_X1 U318 (.ZN(net56025), 
	.A2(A[9]), 
	.A1(B[9]));
   XOR2_X1 U319 (.Z(net56022), 
	.B(A[9]), 
	.A(B[9]));
   AOI21_X1 U321 (.ZN(net73472), 
	.B2(net73491), 
	.B1(net73490), 
	.A(net73492));
   NAND2_X1 U322 (.ZN(net73468), 
	.A2(B[7]), 
	.A1(A[7]));
   NOR2_X1 U323 (.ZN(net73489), 
	.A2(B[7]), 
	.A1(A[7]));
   INV_X1 U324 (.ZN(net69119), 
	.A(net82409));
   INV_X1 U325 (.ZN(net82384), 
	.A(net82378));
   NAND2_X1 U326 (.ZN(net82378), 
	.A2(B[10]), 
	.A1(net82377));
   AND3_X1 U328 (.ZN(net75846), 
	.A3(net56333), 
	.A2(net84167), 
	.A1(net62181));
   NAND2_X1 U329 (.ZN(net58061), 
	.A2(B[52]), 
	.A1(n147));
   NAND2_X1 U330 (.ZN(n147), 
	.A2(net56041), 
	.A1(net58056));
   AND3_X1 U331 (.ZN(net58206), 
	.A3(net58069), 
	.A2(B[52]), 
	.A1(A[50]));
   AND3_X1 U332 (.ZN(net58409), 
	.A3(net58069), 
	.A2(B[52]), 
	.A1(B[50]));
   NAND2_X1 U333 (.ZN(net58069), 
	.A2(net58056), 
	.A1(net58055));
   INV_X1 U334 (.ZN(net58055), 
	.A(net58054));
   OAI21_X1 U335 (.ZN(net58040), 
	.B2(net56041), 
	.B1(net58055), 
	.A(net58056));
   NAND2_X1 U336 (.ZN(net59537), 
	.A2(B[32]), 
	.A1(\carry[32] ));
   INV_X1 U337 (.ZN(net65659), 
	.A(net65693));
   AOI21_X1 U338 (.ZN(net65638), 
	.B2(net65697), 
	.B1(net65658), 
	.A(net65659));
   INV_X1 U340 (.ZN(net65691), 
	.A(net65679));
   INV_X1 U341 (.ZN(net65697), 
	.A(net65709));
   NAND2_X1 U343 (.ZN(net65677), 
	.A2(A[31]), 
	.A1(B[31]));
   NAND2_X1 U344 (.ZN(net65680), 
	.A2(net65679), 
	.A1(A[32]));
   INV_X1 U345 (.ZN(net65671), 
	.A(A[31]));
   AND2_X1 U346 (.ZN(net65709), 
	.A2(B[30]), 
	.A1(net57011));
   AOI21_X1 U347 (.ZN(net65686), 
	.B2(net65687), 
	.B1(net65709), 
	.A(net65678));
   XNOR2_X1 U348 (.ZN(net59519), 
	.B(A[31]), 
	.A(B[31]));
   NAND2_X1 U350 (.ZN(net62307), 
	.A2(net60770), 
	.A1(n149));
   NOR2_X1 U352 (.ZN(n149), 
	.A2(FE_PT1_n213), 
	.A1(n148));
   NOR2_X1 U354 (.ZN(n148), 
	.A2(A[22]), 
	.A1(B[22]));
   NAND2_X1 U355 (.ZN(net62344), 
	.A2(B[21]), 
	.A1(net56569));
   NAND3_X1 U356 (.ZN(net56569), 
	.A3(net55964), 
	.A2(net57089), 
	.A1(net56901));
   NAND2_X1 U357 (.ZN(net56054), 
	.A2(A[21]), 
	.A1(net56569));
   NAND2_X1 U358 (.ZN(net62332), 
	.A2(B[21]), 
	.A1(A[21]));
   AND2_X1 U361 (.ZN(net62309), 
	.A2(B[24]), 
	.A1(net60770));
   XNOR2_X1 U363 (.ZN(net60821), 
	.B(B[21]), 
	.A(A[21]));
   AOI21_X1 U367 (.ZN(net57019), 
	.B2(n155), 
	.B1(n154), 
	.A(n153));
   NAND2_X1 U368 (.ZN(net65272), 
	.A2(A[38]), 
	.A1(net57019));
   INV_X1 U369 (.ZN(n153), 
	.A(n157));
   NAND2_X1 U370 (.ZN(n157), 
	.A2(net65215), 
	.A1(net65153));
   NAND2_X1 U372 (.ZN(net64019), 
	.A2(n700), 
	.A1(net64012));
   NAND2_X1 U374 (.ZN(n155), 
	.A2(net65221), 
	.A1(n159));
   INV_X1 U375 (.ZN(net65221), 
	.A(net65191));
   NAND2_X1 U376 (.ZN(n159), 
	.A2(net73663), 
	.A1(net73570));
   AND2_X1 U377 (.ZN(net73663), 
	.A2(net73561), 
	.A1(net73562));
   NAND2_X1 U379 (.ZN(n154), 
	.A2(n158), 
	.A1(net73554));
   OR2_X1 U380 (.ZN(n158), 
	.A2(net65196), 
	.A1(net65199));
   INV_X1 U381 (.ZN(net73557), 
	.A(net65199));
   AND2_X1 U383 (.ZN(n162), 
	.A2(net84122), 
	.A1(n47));
   INV_X1 U384 (.ZN(n163), 
	.A(net75699));
   INV_X1 U385 (.ZN(net84131), 
	.A(net57080));
   NAND2_X1 U386 (.ZN(n160), 
	.A2(B[43]), 
	.A1(A[43]));
   NAND2_X1 U387 (.ZN(n161), 
	.A2(n163), 
	.A1(A[43]));
   NAND4_X1 U389 (.ZN(net84135), 
	.A4(net56333), 
	.A3(net84167), 
	.A2(n160), 
	.A1(net62181));
   AND3_X1 U390 (.ZN(net75678), 
	.A3(net84122), 
	.A2(net84129), 
	.A1(n47));
   NAND3_X1 U394 (.ZN(n167), 
	.A3(n168), 
	.A2(net79844), 
	.A1(n178));
   NAND2_X1 U395 (.ZN(n168), 
	.A2(A[39]), 
	.A1(\carry[39] ));
   NAND2_X1 U396 (.ZN(net70464), 
	.A2(n170), 
	.A1(n169));
   AND4_X1 U397 (.ZN(n169), 
	.A4(net82338), 
	.A3(n191), 
	.A2(n189), 
	.A1(n190));
   AND3_X1 U398 (.ZN(n170), 
	.A3(n193), 
	.A2(n192), 
	.A1(net82391));
   NAND3_X1 U400 (.ZN(n171), 
	.A3(n316), 
	.A2(n376), 
	.A1(net55819));
   NAND2_X1 U401 (.ZN(n189), 
	.A2(n172), 
	.A1(net82384));
   NAND2_X1 U402 (.ZN(n172), 
	.A2(n241), 
	.A1(n240));
   NAND2_X1 U403 (.ZN(n173), 
	.A2(B[27]), 
	.A1(n207));
   NAND2_X1 U404 (.ZN(n174), 
	.A2(A[27]), 
	.A1(n217));
   NOR2_X1 U406 (.ZN(net82516), 
	.A2(net60779), 
	.A1(net60799));
   NAND3_X1 U408 (.ZN(net82512), 
	.A3(net56371), 
	.A2(net56370), 
	.A1(net79904));
   NAND2_X1 U412 (.ZN(n190), 
	.A2(net82384), 
	.A1(net82542));
   NAND2_X1 U413 (.ZN(n193), 
	.A2(net82423), 
	.A1(net82542));
   NAND2_X1 U414 (.ZN(n191), 
	.A2(net82423), 
	.A1(n172));
   NAND2_X1 U415 (.ZN(n194), 
	.A2(net82394), 
	.A1(n172));
   NAND2_X1 U416 (.ZN(net77826), 
	.A2(n64), 
	.A1(net82333));
   NAND2_X1 U419 (.ZN(n178), 
	.A2(B[39]), 
	.A1(net56856));
   NAND2_X1 U420 (.ZN(n179), 
	.A2(B[28]), 
	.A1(\carry[28] ));
   AOI21_X1 U421 (.ZN(n197), 
	.B2(net82402), 
	.B1(net82405), 
	.A(n186));
   NAND2_X1 U422 (.ZN(n184), 
	.A2(n172), 
	.A1(net82427));
   AOI21_X1 U423 (.ZN(net55836), 
	.B2(n271), 
	.B1(net70464), 
	.A(net70465));
   INV_X1 U425 (.ZN(net82365), 
	.A(A[11]));
   INV_X1 U427 (.ZN(net82369), 
	.A(net70500));
   INV_X1 U428 (.ZN(net82373), 
	.A(net70488));
   NOR2_X1 U429 (.ZN(n186), 
	.A2(net82338), 
	.A1(net82373));
   NAND2_X1 U430 (.ZN(net82381), 
	.A2(net73518), 
	.A1(n187));
   NOR2_X1 U431 (.ZN(n188), 
	.A2(net82387), 
	.A1(net82383));
   NOR2_X1 U432 (.ZN(n187), 
	.A2(net82355), 
	.A1(A[10]));
   NAND3_X1 U433 (.ZN(n208), 
	.A3(n205), 
	.A2(n206), 
	.A1(n179));
   NAND2_X1 U434 (.ZN(net62177), 
	.A2(B[29]), 
	.A1(n208));
   NAND2_X1 U436 (.ZN(n206), 
	.A2(A[28]), 
	.A1(n209));
   NAND3_X1 U437 (.ZN(n209), 
	.A3(n204), 
	.A2(n173), 
	.A1(n174));
   NAND3_X1 U439 (.ZN(\carry[29] ), 
	.A3(n205), 
	.A2(n179), 
	.A1(n206));
   NAND3_X1 U440 (.ZN(\carry[28] ), 
	.A3(n204), 
	.A2(n174), 
	.A1(n173));
   NAND3_X1 U442 (.ZN(n217), 
	.A3(net55592), 
	.A2(net73589), 
	.A1(n68));
   NAND2_X1 U444 (.ZN(n205), 
	.A2(B[28]), 
	.A1(A[28]));
   XOR2_X1 U445 (.Z(net56060), 
	.B(B[28]), 
	.A(A[28]));
   NAND3_X1 U451 (.ZN(n207), 
	.A3(net55592), 
	.A2(n68), 
	.A1(net73589));
   NAND2_X1 U452 (.ZN(n204), 
	.A2(B[27]), 
	.A1(A[27]));
   XOR2_X1 U453 (.Z(net55595), 
	.B(B[27]), 
	.A(A[27]));
   NAND2_X1 U456 (.ZN(net67379), 
	.A2(n218), 
	.A1(net70524));
   AND2_X1 U457 (.ZN(n218), 
	.A2(net67373), 
	.A1(A[15]));
   XNOR2_X1 U459 (.ZN(net67389), 
	.B(A[16]), 
	.A(B[16]));
   NAND3_X1 U465 (.ZN(\carry[39] ), 
	.A3(net56739), 
	.A2(n219), 
	.A1(net65272));
   NAND2_X1 U466 (.ZN(n219), 
	.A2(B[38]), 
	.A1(net64058));
   AOI21_X1 U467 (.ZN(net64058), 
	.B2(n221), 
	.B1(n220), 
	.A(n222));
   NAND2_X1 U468 (.ZN(n223), 
	.A2(net65153), 
	.A1(net65215));
   NAND2_X1 U469 (.ZN(n221), 
	.A2(n224), 
	.A1(net73564));
   OR2_X1 U470 (.ZN(n224), 
	.A2(net65196), 
	.A1(net65202));
   NAND2_X1 U472 (.ZN(n220), 
	.A2(n226), 
	.A1(n225));
   OR2_X1 U473 (.ZN(n226), 
	.A2(net65221), 
	.A1(n227));
   INV_X1 U474 (.ZN(n227), 
	.A(net65188));
   NAND2_X1 U475 (.ZN(n225), 
	.A2(net73675), 
	.A1(net73663));
   NAND2_X1 U478 (.ZN(net56333), 
	.A2(B[42]), 
	.A1(A[42]));
   XOR2_X1 U479 (.Z(net56332), 
	.B(B[42]), 
	.A(A[42]));
   NAND3_X1 U481 (.ZN(net56427), 
	.A3(net79904), 
	.A2(net56371), 
	.A1(n52));
   AND2_X1 U482 (.ZN(net56370), 
	.A2(n78), 
	.A1(n230));
   NAND2_X1 U483 (.ZN(n230), 
	.A2(n80), 
	.A1(n167));
   INV_X1 U487 (.ZN(n231), 
	.A(A[40]));
   NAND2_X1 U489 (.ZN(net79832), 
	.A2(B[40]), 
	.A1(A[40]));
   NAND2_X1 U490 (.ZN(n233), 
	.A2(A[40]), 
	.A1(B[41]));
   NAND2_X1 U491 (.ZN(n234), 
	.A2(B[40]), 
	.A1(B[41]));
   NAND2_X1 U492 (.ZN(net79849), 
	.A2(B[41]), 
	.A1(net79851));
   NAND2_X1 U493 (.ZN(net79855), 
	.A2(n231), 
	.A1(n632));
   NAND2_X1 U494 (.ZN(net79856), 
	.A2(n233), 
	.A1(n234));
   XNOR2_X1 U495 (.ZN(n235), 
	.B(B[39]), 
	.A(A[39]));
   INV_X1 U496 (.ZN(net56639), 
	.A(n235));
   XNOR2_X1 U497 (.ZN(n236), 
	.B(B[40]), 
	.A(A[40]));
   INV_X1 U498 (.ZN(net56562), 
	.A(n236));
   NAND2_X1 U499 (.ZN(net56817), 
	.A2(net58057), 
	.A1(n237));
   AND2_X1 U500 (.ZN(n237), 
	.A2(n238), 
	.A1(net58447));
   AND2_X1 U501 (.ZN(n238), 
	.A2(net58242), 
	.A1(net58038));
   INV_X1 U502 (.ZN(net58038), 
	.A(net58040));
   NAND2_X1 U503 (.ZN(net58121), 
	.A2(net58038), 
	.A1(net58037));
   NAND2_X1 U504 (.ZN(net56144), 
	.A2(B[53]), 
	.A1(A[53]));
   AND2_X1 U507 (.ZN(n239), 
	.A2(n243), 
	.A1(net77768));
   NAND2_X1 U508 (.ZN(n240), 
	.A2(net77818), 
	.A1(n146));
   OR2_X1 U509 (.ZN(n241), 
	.A2(net73472), 
	.A1(net77817));
   INV_X1 U510 (.ZN(net77817), 
	.A(A[9]));
   AND2_X1 U511 (.ZN(net77766), 
	.A2(A[3]), 
	.A1(A[2]));
   INV_X1 U512 (.ZN(net55812), 
	.A(net77785));
   INV_X1 U513 (.ZN(net55808), 
	.A(n244));
   XNOR2_X1 U514 (.ZN(n244), 
	.B(B[1]), 
	.A(A[1]));
   NOR2_X1 U515 (.ZN(n242), 
	.A2(A[1]), 
	.A1(\carry[1] ));
   OAI21_X1 U516 (.ZN(net56545), 
	.B2(n242), 
	.B1(n794), 
	.A(net56561));
   NAND2_X1 U518 (.ZN(n243), 
	.A2(n92), 
	.A1(net77765));
   NAND3_X1 U519 (.ZN(net56859), 
	.A3(n245), 
	.A2(n8), 
	.A1(n54));
   NAND2_X1 U520 (.ZN(net58227), 
	.A2(B[48]), 
	.A1(net56859));
   NAND2_X1 U525 (.ZN(n245), 
	.A2(B[47]), 
	.A1(A[47]));
   XOR2_X1 U526 (.Z(net55579), 
	.B(B[47]), 
	.A(A[47]));
   NOR2_X1 U528 (.ZN(n248), 
	.A2(net65683), 
	.A1(n7));
   NAND2_X1 U530 (.ZN(n249), 
	.A2(A[45]), 
	.A1(net75678));
   INV_X1 U531 (.ZN(net57080), 
	.A(net75846));
   NAND2_X1 U532 (.ZN(net75723), 
	.A2(net75725), 
	.A1(n250));
   INV_X1 U533 (.ZN(net57069), 
	.A(net75743));
   NAND2_X1 U534 (.ZN(n250), 
	.A2(n552), 
	.A1(net75720));
   INV_X1 U535 (.ZN(net55822), 
	.A(net75759));
   NOR2_X1 U536 (.ZN(net75699), 
	.A2(B[43]), 
	.A1(net75831));
   AND2_X1 U537 (.ZN(net67433), 
	.A2(A[15]), 
	.A1(net70524));
   AND2_X1 U538 (.ZN(net67429), 
	.A2(A[15]), 
	.A1(net67373));
   XOR2_X1 U539 (.Z(net56368), 
	.B(A[41]), 
	.A(B[41]));
   AND2_X1 U540 (.ZN(net59538), 
	.A2(net65686), 
	.A1(n248));
   AND2_X1 U541 (.ZN(net73660), 
	.A2(n248), 
	.A1(net65686));
   INV_X1 U542 (.ZN(net65675), 
	.A(A[32]));
   INV_X1 U543 (.ZN(net65687), 
	.A(net65680));
   XOR2_X1 U544 (.Z(net56044), 
	.B(B[32]), 
	.A(A[32]));
   NAND2_X1 U545 (.ZN(net56045), 
	.A2(B[32]), 
	.A1(A[32]));
   NAND2_X1 U546 (.ZN(net65183), 
	.A2(n746), 
	.A1(net65181));
   AND2_X1 U547 (.ZN(net73675), 
	.A2(net65188), 
	.A1(net73570));
   NAND3_X1 U548 (.ZN(n251), 
	.A3(n386), 
	.A2(net60691), 
	.A1(n313));
   INV_X1 U549 (.ZN(net73634), 
	.A(net73494));
   AND2_X1 U551 (.ZN(n253), 
	.A2(n292), 
	.A1(net56739));
   NAND2_X1 U552 (.ZN(n292), 
	.A2(net65225), 
	.A1(n227));
   NAND3_X1 U553 (.ZN(n254), 
	.A3(n346), 
	.A2(n239), 
	.A1(net62205));
   NAND2_X1 U555 (.ZN(net73589), 
	.A2(A[26]), 
	.A1(n251));
   NAND3_X1 U556 (.ZN(n255), 
	.A3(net56045), 
	.A2(net59537), 
	.A1(net73660));
   AND2_X1 U558 (.ZN(n266), 
	.A2(net65196), 
	.A1(net65197));
   NAND2_X1 U559 (.ZN(n257), 
	.A2(net65197), 
	.A1(net65196));
   NAND2_X1 U560 (.ZN(net73570), 
	.A2(net62140), 
	.A1(n284));
   NAND2_X1 U561 (.ZN(net73562), 
	.A2(n267), 
	.A1(n268));
   NAND3_X1 U562 (.ZN(n258), 
	.A3(n330), 
	.A2(n331), 
	.A1(n332));
   NAND2_X1 U563 (.ZN(n259), 
	.A2(B[4]), 
	.A1(n254));
   NAND3_X1 U564 (.ZN(\carry[6] ), 
	.A3(n331), 
	.A2(n330), 
	.A1(n332));
   NAND2_X1 U565 (.ZN(n260), 
	.A2(net70488), 
	.A1(net70464));
   OR2_X1 U570 (.ZN(net73518), 
	.A2(net73472), 
	.A1(n615));
   NAND2_X1 U571 (.ZN(net56341), 
	.A2(net73472), 
	.A1(net73473));
   INV_X1 U572 (.ZN(net73494), 
	.A(n146));
   NAND2_X1 U573 (.ZN(net73488), 
	.A2(B[6]), 
	.A1(\carry[6] ));
   INV_X1 U574 (.ZN(n263), 
	.A(A[8]));
   XNOR2_X1 U575 (.ZN(net72085), 
	.B(B[8]), 
	.A(A[8]));
   NAND2_X1 U577 (.ZN(net73491), 
	.A2(n635), 
	.A1(n263));
   NAND2_X1 U578 (.ZN(net73498), 
	.A2(B[8]), 
	.A1(A[8]));
   INV_X1 U579 (.ZN(net73492), 
	.A(net73498));
   NAND2_X1 U580 (.ZN(net73487), 
	.A2(B[6]), 
	.A1(A[6]));
   XNOR2_X1 U581 (.ZN(n265), 
	.B(A[6]), 
	.A(B[6]));
   NAND2_X1 U582 (.ZN(net65288), 
	.A2(net73570), 
	.A1(net73663));
   INV_X1 U585 (.ZN(net65181), 
	.A(A[35]));
   INV_X1 U587 (.ZN(n267), 
	.A(n295));
   NAND3_X1 U588 (.ZN(n268), 
	.A3(net56045), 
	.A2(net59538), 
	.A1(net59537));
   INV_X1 U590 (.ZN(net56313), 
	.A(net72085));
   INV_X1 U591 (.ZN(net56309), 
	.A(net72087));
   AND3_X1 U593 (.ZN(n269), 
	.A3(n278), 
	.A2(net70527), 
	.A1(n260));
   NAND3_X1 U594 (.ZN(net70524), 
	.A3(net55837), 
	.A2(net55836), 
	.A1(n269));
   INV_X1 U595 (.ZN(net70474), 
	.A(A[12]));
   INV_X1 U597 (.ZN(n273), 
	.A(A[13]));
   NAND2_X1 U599 (.ZN(net70482), 
	.A2(n270), 
	.A1(net69089));
   NAND2_X1 U600 (.ZN(net70483), 
	.A2(net70443), 
	.A1(A[14]));
   NOR2_X1 U601 (.ZN(n274), 
	.A2(n555), 
	.A1(net70483));
   NOR2_X1 U602 (.ZN(net69139), 
	.A2(net70474), 
	.A1(net70487));
   AOI21_X1 U604 (.ZN(net70456), 
	.B2(net70464), 
	.B1(A[12]), 
	.A(net70482));
   NAND2_X1 U605 (.ZN(n270), 
	.A2(B[13]), 
	.A1(A[13]));
   INV_X1 U606 (.ZN(net69124), 
	.A(n270));
   INV_X1 U607 (.ZN(net70487), 
	.A(net70464));
   NAND2_X1 U608 (.ZN(net70443), 
	.A2(n529), 
	.A1(n273));
   INV_X1 U609 (.ZN(net70495), 
	.A(net70483));
   NAND2_X1 U610 (.ZN(n276), 
	.A2(A[12]), 
	.A1(net70495));
   INV_X1 U611 (.ZN(n277), 
	.A(n274));
   NAND2_X1 U612 (.ZN(n271), 
	.A2(n276), 
	.A1(n277));
   AND2_X1 U614 (.ZN(n278), 
	.A2(n280), 
	.A1(net69117));
   AND3_X1 U615 (.ZN(net69188), 
	.A3(n278), 
	.A2(n69), 
	.A1(net69119));
   NAND2_X1 U616 (.ZN(n280), 
	.A2(B[14]), 
	.A1(net69124));
   INV_X1 U617 (.ZN(net55925), 
	.A(net69139));
   NAND2_X1 U618 (.ZN(net69089), 
	.A2(B[12]), 
	.A1(A[12]));
   INV_X1 U620 (.ZN(net69126), 
	.A(net69089));
   INV_X1 U621 (.ZN(net55927), 
	.A(net69132));
   XNOR2_X1 U622 (.ZN(n281), 
	.B(A[12]), 
	.A(B[12]));
   INV_X1 U623 (.ZN(net55923), 
	.A(n281));
   NAND2_X1 U624 (.ZN(n282), 
	.A2(B[25]), 
	.A1(net82511));
   NAND3_X1 U625 (.ZN(net67466), 
	.A3(net55837), 
	.A2(n269), 
	.A1(net67456));
   NAND2_X1 U626 (.ZN(n297), 
	.A2(A[33]), 
	.A1(n284));
   NAND2_X1 U628 (.ZN(net67357), 
	.A2(B[15]), 
	.A1(net67466));
   INV_X1 U630 (.ZN(net67368), 
	.A(A[16]));
   NAND2_X1 U631 (.ZN(net67355), 
	.A2(B[15]), 
	.A1(A[15]));
   NAND2_X1 U632 (.ZN(net67373), 
	.A2(net67368), 
	.A1(n454));
   XNOR2_X1 U633 (.ZN(n283), 
	.B(B[15]), 
	.A(A[15]));
   INV_X1 U634 (.ZN(net55691), 
	.A(n283));
   INV_X1 U635 (.ZN(net55599), 
	.A(net67389));
   INV_X1 U636 (.ZN(net67391), 
	.A(net67433));
   NAND2_X1 U637 (.ZN(net67385), 
	.A2(net67429), 
	.A1(\carry[15] ));
   NAND3_X1 U639 (.ZN(n284), 
	.A3(net56045), 
	.A2(net73660), 
	.A1(net59537));
   INV_X1 U641 (.ZN(net65704), 
	.A(n101));
   NAND2_X1 U642 (.ZN(net65321), 
	.A2(n74), 
	.A1(net69203));
   NAND2_X1 U645 (.ZN(net65160), 
	.A2(net65288), 
	.A1(net65221));
   NAND2_X1 U647 (.ZN(net65309), 
	.A2(n253), 
	.A1(n291));
   NAND2_X1 U649 (.ZN(net65201), 
	.A2(B[35]), 
	.A1(A[35]));
   AND3_X1 U650 (.ZN(net64053), 
	.A3(net65160), 
	.A2(n257), 
	.A1(net65188));
   NOR2_X1 U651 (.ZN(net65159), 
	.A2(net65199), 
	.A1(n266));
   NAND2_X1 U652 (.ZN(net56856), 
	.A2(net65272), 
	.A1(net65290));
   NAND2_X1 U654 (.ZN(net65188), 
	.A2(A[36]), 
	.A1(n290));
   NAND2_X1 U655 (.ZN(net65199), 
	.A2(net65153), 
	.A1(net65188));
   INV_X1 U656 (.ZN(n290), 
	.A(net65201));
   NAND3_X1 U658 (.ZN(n291), 
	.A3(net65221), 
	.A2(net65225), 
	.A1(net65288));
   XNOR2_X1 U659 (.ZN(n293), 
	.B(B[35]), 
	.A(A[35]));
   INV_X1 U660 (.ZN(net55683), 
	.A(n293));
   NAND2_X1 U665 (.ZN(net62110), 
	.A2(n268), 
	.A1(B[33]));
   INV_X1 U667 (.ZN(net55587), 
	.A(net64020));
   INV_X1 U668 (.ZN(net55583), 
	.A(net64022));
   INV_X1 U669 (.ZN(net55672), 
	.A(net64053));
   NAND2_X1 U670 (.ZN(n295), 
	.A2(B[33]), 
	.A1(net62130));
   INV_X1 U672 (.ZN(net62132), 
	.A(net62130));
   NAND2_X1 U673 (.ZN(net62129), 
	.A2(A[33]), 
	.A1(net62130));
   NAND2_X1 U674 (.ZN(net62111), 
	.A2(A[33]), 
	.A1(B[33]));
   XNOR2_X1 U675 (.ZN(net62145), 
	.B(A[33]), 
	.A(B[33]));
   INV_X1 U676 (.ZN(net55830), 
	.A(net62338));
   NAND2_X1 U679 (.ZN(n296), 
	.A2(A[4]), 
	.A1(n254));
   NAND2_X1 U682 (.ZN(net62194), 
	.A2(B[43]), 
	.A1(net57080));
   NAND2_X1 U683 (.ZN(net62139), 
	.A2(net62140), 
	.A1(n255));
   OR2_X1 U685 (.ZN(net58447), 
	.A2(net58244), 
	.A1(net58329));
   INV_X1 U687 (.ZN(n299), 
	.A(A[34]));
   OAI21_X1 U688 (.ZN(net62131), 
	.B2(net62111), 
	.B1(net62132), 
	.A(n300));
   NAND2_X1 U689 (.ZN(net62130), 
	.A2(n769), 
	.A1(n299));
   NAND2_X1 U690 (.ZN(n300), 
	.A2(B[34]), 
	.A1(A[34]));
   INV_X1 U691 (.ZN(net62140), 
	.A(net62129));
   INV_X1 U692 (.ZN(net56048), 
	.A(net62145));
   XNOR2_X1 U693 (.ZN(n301), 
	.B(B[34]), 
	.A(A[34]));
   INV_X1 U694 (.ZN(net55826), 
	.A(n301));
   NAND3_X1 U695 (.ZN(n302), 
	.A3(n386), 
	.A2(n282), 
	.A1(net60691));
   INV_X1 U698 (.ZN(net60835), 
	.A(net75853));
   INV_X1 U700 (.ZN(n304), 
	.A(A[23]));
   NAND2_X1 U701 (.ZN(net60794), 
	.A2(B[23]), 
	.A1(A[23]));
   NAND2_X1 U702 (.ZN(net60770), 
	.A2(n304), 
	.A1(n806));
   XNOR2_X1 U706 (.ZN(net60649), 
	.B(B[22]), 
	.A(A[22]));
   INV_X1 U708 (.ZN(net60813), 
	.A(net60794));
   INV_X1 U710 (.ZN(net56052), 
	.A(net60821));
   INV_X1 U712 (.ZN(net56437), 
	.A(net60647));
   INV_X1 U713 (.ZN(net56056), 
	.A(net60649));
   INV_X1 U715 (.ZN(net58404), 
	.A(net58327));
   INV_X1 U716 (.ZN(net56433), 
	.A(net59517));
   INV_X1 U717 (.ZN(net56154), 
	.A(net59519));
   AND2_X1 U718 (.ZN(n305), 
	.A2(net58242), 
	.A1(net58447));
   INV_X1 U720 (.ZN(net58422), 
	.A(A[50]));
   INV_X1 U721 (.ZN(net58389), 
	.A(net58243));
   NAND2_X1 U722 (.ZN(net58399), 
	.A2(n402), 
	.A1(net58422));
   INV_X1 U723 (.ZN(net58323), 
	.A(net58329));
   NAND2_X1 U725 (.ZN(n307), 
	.A2(A[55]), 
	.A1(n171));
   NAND2_X1 U727 (.ZN(net58282), 
	.A2(n305), 
	.A1(net58057));
   INV_X1 U728 (.ZN(net58037), 
	.A(net58282));
   NAND2_X1 U729 (.ZN(net58228), 
	.A2(net58327), 
	.A1(A[50]));
   AND2_X1 U730 (.ZN(net58210), 
	.A2(net58054), 
	.A1(A[50]));
   XNOR2_X1 U732 (.ZN(n308), 
	.B(B[48]), 
	.A(A[48]));
   INV_X1 U733 (.ZN(net56150), 
	.A(n308));
   INV_X1 U734 (.ZN(net56040), 
	.A(net58236));
   INV_X1 U735 (.ZN(net56036), 
	.A(net58238));
   NAND2_X1 U736 (.ZN(net58226), 
	.A2(B[48]), 
	.A1(A[48]));
   OR2_X1 U737 (.ZN(net58244), 
	.A2(net58243), 
	.A1(net58222));
   INV_X1 U738 (.ZN(net58243), 
	.A(net58210));
   NAND2_X1 U739 (.ZN(n309), 
	.A2(A[52]), 
	.A1(net58121));
   INV_X1 U741 (.ZN(n311), 
	.A(A[51]));
   NAND2_X1 U742 (.ZN(net58054), 
	.A2(FE_PT1_n380), 
	.A1(n311));
   NAND2_X1 U743 (.ZN(net58056), 
	.A2(B[51]), 
	.A1(A[51]));
   XNOR2_X1 U744 (.ZN(n312), 
	.B(B[51]), 
	.A(A[51]));
   INV_X1 U745 (.ZN(net56571), 
	.A(n312));
   INV_X1 U747 (.ZN(net58078), 
	.A(net58315));
   NAND2_X1 U748 (.ZN(n313), 
	.A2(B[25]), 
	.A1(net60880));
   NAND2_X1 U750 (.ZN(net57089), 
	.A2(A[20]), 
	.A1(\carry[20] ));
   NAND2_X1 U753 (.ZN(net55681), 
	.A2(A[45]), 
	.A1(\carry[45] ));
   NAND2_X1 U754 (.ZN(n357), 
	.A2(A[59]), 
	.A1(n15));
   NAND2_X1 U755 (.ZN(n316), 
	.A2(A[54]), 
	.A1(n132));
   NAND2_X1 U759 (.ZN(n319), 
	.A2(B[56]), 
	.A1(n321));
   NAND3_X1 U764 (.ZN(n321), 
	.A3(n382), 
	.A2(n307), 
	.A1(n57));
   AND2_X1 U765 (.ZN(net57022), 
	.A2(A[0]), 
	.A1(B[0]));
   NAND3_X1 U766 (.ZN(n322), 
	.A3(n348), 
	.A2(n296), 
	.A1(n259));
   NAND3_X1 U768 (.ZN(\carry[5] ), 
	.A3(n296), 
	.A2(n348), 
	.A1(n259));
   NAND3_X1 U769 (.ZN(net57011), 
	.A3(n364), 
	.A2(n365), 
	.A1(net62177));
   NAND2_X1 U772 (.ZN(net56901), 
	.A2(B[20]), 
	.A1(n337));
   NAND2_X1 U774 (.ZN(n324), 
	.A2(B[45]), 
	.A1(net57069));
   XOR2_X1 U775 (.Z(SUM[18]), 
	.B(net56887), 
	.A(n10));
   NAND3_X1 U776 (.ZN(n325), 
	.A3(net56140), 
	.A2(n309), 
	.A1(net56142));
   NAND2_X1 U777 (.ZN(n326), 
	.A2(B[59]), 
	.A1(n15));
   NAND3_X1 U779 (.ZN(n327), 
	.A3(n356), 
	.A2(n357), 
	.A1(n326));
   NAND3_X1 U780 (.ZN(\carry[15] ), 
	.A3(net55837), 
	.A2(net55836), 
	.A1(net69188));
   NAND2_X1 U781 (.ZN(n328), 
	.A2(A[58]), 
	.A1(\carry[58] ));
   XOR2_X1 U783 (.Z(n329), 
	.B(B[5]), 
	.A(A[5]));
   XOR2_X1 U784 (.Z(SUM[5]), 
	.B(n322), 
	.A(n329));
   NAND2_X1 U785 (.ZN(n330), 
	.A2(B[5]), 
	.A1(A[5]));
   NAND2_X1 U786 (.ZN(n331), 
	.A2(A[5]), 
	.A1(\carry[5] ));
   NAND2_X1 U787 (.ZN(n332), 
	.A2(B[5]), 
	.A1(n322));
   XOR2_X1 U788 (.Z(SUM[6]), 
	.B(n258), 
	.A(net56753));
   NAND2_X1 U789 (.ZN(net56755), 
	.A2(A[6]), 
	.A1(n258));
   NAND3_X1 U790 (.ZN(n334), 
	.A3(n324), 
	.A2(net55682), 
	.A1(n249));
   NAND3_X1 U791 (.ZN(n333), 
	.A3(net55680), 
	.A2(net55682), 
	.A1(n249));
   XOR2_X1 U792 (.Z(n335), 
	.B(A[38]), 
	.A(B[38]));
   XOR2_X1 U793 (.Z(SUM[38]), 
	.B(n335), 
	.A(net65126));
   NAND2_X1 U794 (.ZN(net56739), 
	.A2(A[38]), 
	.A1(B[38]));
   XOR2_X1 U796 (.Z(SUM[39]), 
	.B(net56639), 
	.A(net56856));
   NAND2_X1 U797 (.ZN(SUM[63]), 
	.A2(net56650), 
	.A1(net56651));
   INV_X1 U798 (.ZN(net56649), 
	.A(net56540));
   INV_X1 U799 (.ZN(net56540), 
	.A(net55816));
   NAND3_X1 U801 (.ZN(\carry[20] ), 
	.A3(n368), 
	.A2(net57091), 
	.A1(n369));
   INV_X1 U802 (.ZN(net56598), 
	.A(net56477));
   XOR2_X1 U803 (.Z(SUM[40]), 
	.B(net56562), 
	.A(n48));
   XOR2_X1 U804 (.Z(SUM[51]), 
	.B(net56571), 
	.A(net57006));
   NAND2_X1 U805 (.ZN(net56561), 
	.A2(\carry[1] ), 
	.A1(A[1]));
   XOR2_X1 U812 (.Z(SUM[30]), 
	.B(net56433), 
	.A(net57011));
   XOR2_X1 U813 (.Z(SUM[23]), 
	.B(net56437), 
	.A(net56471));
   XOR2_X1 U816 (.Z(SUM[41]), 
	.B(net56368), 
	.A(net56630));
   XOR2_X1 U817 (.Z(SUM[42]), 
	.B(net56427), 
	.A(net56332));
   XOR2_X1 U818 (.Z(SUM[43]), 
	.B(net57080), 
	.A(net56336));
   XOR2_X1 U819 (.Z(SUM[7]), 
	.B(net73634), 
	.A(net56309));
   XOR2_X1 U820 (.Z(SUM[8]), 
	.B(n264), 
	.A(net56313));
   XOR2_X1 U823 (.Z(n345), 
	.B(B[3]), 
	.A(A[3]));
   XOR2_X1 U824 (.Z(SUM[3]), 
	.B(\carry[3] ), 
	.A(n345));
   NAND2_X1 U825 (.ZN(n346), 
	.A2(B[3]), 
	.A1(A[3]));
   XOR2_X1 U826 (.Z(n347), 
	.B(B[4]), 
	.A(A[4]));
   XOR2_X1 U827 (.Z(SUM[4]), 
	.B(n254), 
	.A(n347));
   NAND2_X1 U828 (.ZN(n348), 
	.A2(B[4]), 
	.A1(A[4]));
   NAND3_X1 U829 (.ZN(n349), 
	.A3(n328), 
	.A2(n354), 
	.A1(net56549));
   NAND3_X1 U830 (.ZN(n350), 
	.A3(n356), 
	.A2(n326), 
	.A1(n357));
   XOR2_X1 U832 (.Z(n352), 
	.B(A[58]), 
	.A(B[58]));
   XOR2_X1 U833 (.Z(SUM[58]), 
	.B(n352), 
	.A(n141));
   NAND2_X1 U834 (.ZN(n354), 
	.A2(A[58]), 
	.A1(B[58]));
   XOR2_X1 U836 (.Z(n355), 
	.B(B[59]), 
	.A(A[59]));
   XOR2_X1 U837 (.Z(SUM[59]), 
	.B(n349), 
	.A(n355));
   NAND2_X1 U838 (.ZN(n356), 
	.A2(B[59]), 
	.A1(A[59]));
   XOR2_X1 U839 (.Z(n359), 
	.B(B[60]), 
	.A(A[60]));
   NAND2_X1 U840 (.ZN(net56225), 
	.A2(B[60]), 
	.A1(A[60]));
   NAND2_X1 U841 (.ZN(net56226), 
	.A2(A[60]), 
	.A1(n327));
   NAND2_X1 U842 (.ZN(net56227), 
	.A2(B[60]), 
	.A1(n327));
   XOR2_X1 U844 (.Z(n361), 
	.B(B[52]), 
	.A(A[52]));
   XOR2_X1 U845 (.Z(SUM[52]), 
	.B(n361), 
	.A(net58121));
   NAND2_X1 U846 (.ZN(net56140), 
	.A2(B[52]), 
	.A1(A[52]));
   XOR2_X1 U847 (.Z(n362), 
	.B(B[53]), 
	.A(A[53]));
   XOR2_X1 U848 (.Z(SUM[53]), 
	.B(n362), 
	.A(n325));
   XOR2_X1 U849 (.Z(SUM[48]), 
	.B(net56150), 
	.A(n6));
   XOR2_X1 U850 (.Z(SUM[31]), 
	.B(net56154), 
	.A(net56628));
   XOR2_X1 U851 (.Z(SUM[49]), 
	.B(net56036), 
	.A(net58323));
   XOR2_X1 U852 (.Z(SUM[50]), 
	.B(net58327), 
	.A(net56040));
   XOR2_X1 U853 (.Z(SUM[32]), 
	.B(net65638), 
	.A(net56044));
   XOR2_X1 U854 (.Z(SUM[33]), 
	.B(n284), 
	.A(net56048));
   XOR2_X1 U855 (.Z(SUM[21]), 
	.B(net56569), 
	.A(net56052));
   XOR2_X1 U856 (.Z(SUM[22]), 
	.B(net60835), 
	.A(net56056));
   XOR2_X1 U857 (.Z(SUM[28]), 
	.B(n209), 
	.A(net56060));
   XOR2_X1 U858 (.Z(n363), 
	.B(B[29]), 
	.A(A[29]));
   XOR2_X1 U859 (.Z(SUM[29]), 
	.B(n208), 
	.A(n363));
   NAND2_X1 U860 (.ZN(n364), 
	.A2(B[29]), 
	.A1(A[29]));
   NAND2_X1 U861 (.ZN(n365), 
	.A2(A[29]), 
	.A1(\carry[29] ));
   XOR2_X1 U864 (.Z(SUM[9]), 
	.B(net56022), 
	.A(net56341));
   XOR2_X1 U865 (.Z(n367), 
	.B(B[19]), 
	.A(A[19]));
   XOR2_X1 U866 (.Z(SUM[19]), 
	.B(n116), 
	.A(n367));
   NAND2_X1 U867 (.ZN(n368), 
	.A2(B[19]), 
	.A1(A[19]));
   NAND2_X1 U868 (.ZN(n369), 
	.A2(A[19]), 
	.A1(\carry[19] ));
   XOR2_X1 U869 (.Z(n370), 
	.B(B[20]), 
	.A(A[20]));
   XOR2_X1 U870 (.Z(SUM[20]), 
	.B(n337), 
	.A(n370));
   NAND2_X1 U871 (.ZN(net55964), 
	.A2(B[20]), 
	.A1(A[20]));
   XOR2_X1 U874 (.Z(SUM[10]), 
	.B(net77826), 
	.A(net55967));
   XOR2_X1 U876 (.Z(SUM[12]), 
	.B(net70464), 
	.A(net55923));
   XOR2_X1 U877 (.Z(SUM[13]), 
	.B(net56020), 
	.A(net55927));
   NAND3_X1 U878 (.ZN(n372), 
	.A3(n57), 
	.A2(n382), 
	.A1(n307));
   XOR2_X1 U881 (.Z(SUM[1]), 
	.B(\carry[1] ), 
	.A(net55808));
   XOR2_X1 U882 (.Z(SUM[2]), 
	.B(net56545), 
	.A(net55812));
   XOR2_X1 U883 (.Z(net55816), 
	.B(A[63]), 
	.A(B[63]));
   XOR2_X1 U884 (.Z(n374), 
	.B(A[54]), 
	.A(B[54]));
   XOR2_X1 U885 (.Z(SUM[54]), 
	.B(n374), 
	.A(n132));
   NAND2_X1 U886 (.ZN(n376), 
	.A2(A[54]), 
	.A1(B[54]));
   XOR2_X1 U887 (.Z(SUM[44]), 
	.B(net55822), 
	.A(net56476));
   XOR2_X1 U888 (.Z(SUM[34]), 
	.B(net55826), 
	.A(net56158));
   XOR2_X1 U889 (.Z(SUM[24]), 
	.B(net55830), 
	.A(net60758));
   XOR2_X1 U890 (.Z(n377), 
	.B(A[14]), 
	.A(B[14]));
   XOR2_X1 U891 (.Z(SUM[14]), 
	.B(n377), 
	.A(net56808));
   NAND2_X1 U892 (.ZN(net55837), 
	.A2(A[14]), 
	.A1(B[14]));
   NAND3_X1 U893 (.ZN(n378), 
	.A3(n319), 
	.A2(n388), 
	.A1(n389));
   XOR2_X1 U895 (.Z(n380), 
	.B(A[55]), 
	.A(B[55]));
   XOR2_X1 U896 (.Z(SUM[55]), 
	.B(n380), 
	.A(n171));
   NAND2_X1 U897 (.ZN(n382), 
	.A2(A[55]), 
	.A1(B[55]));
   XOR2_X1 U898 (.Z(n383), 
	.B(A[45]), 
	.A(B[45]));
   XOR2_X1 U899 (.Z(SUM[45]), 
	.B(n383), 
	.A(net57069));
   NAND2_X1 U900 (.ZN(net55682), 
	.A2(A[45]), 
	.A1(B[45]));
   XOR2_X1 U901 (.Z(SUM[35]), 
	.B(net55683), 
	.A(net65288));
   XOR2_X1 U902 (.Z(n384), 
	.B(A[25]), 
	.A(B[25]));
   XOR2_X1 U903 (.Z(SUM[25]), 
	.B(n384), 
	.A(net60880));
   NAND2_X1 U905 (.ZN(n386), 
	.A2(A[25]), 
	.A1(B[25]));
   XOR2_X1 U906 (.Z(SUM[15]), 
	.B(net55691), 
	.A(net67466));
   NAND3_X1 U908 (.ZN(\carry[47] ), 
	.A3(n392), 
	.A2(n56), 
	.A1(n14));
   AND2_X1 U909 (.ZN(\carry[1] ), 
	.A2(B[0]), 
	.A1(A[0]));
   XOR2_X1 U910 (.Z(n387), 
	.B(B[56]), 
	.A(A[56]));
   XOR2_X1 U911 (.Z(SUM[56]), 
	.B(n372), 
	.A(n387));
   NAND2_X1 U912 (.ZN(n388), 
	.A2(B[56]), 
	.A1(A[56]));
   XOR2_X1 U914 (.Z(SUM[57]), 
	.B(n378), 
	.A(net55571));
   XOR2_X1 U915 (.Z(n391), 
	.B(B[46]), 
	.A(A[46]));
   XOR2_X1 U916 (.Z(SUM[46]), 
	.B(n391), 
	.A(n334));
   NAND2_X1 U917 (.ZN(n392), 
	.A2(B[46]), 
	.A1(A[46]));
   XOR2_X1 U919 (.Z(SUM[47]), 
	.B(n61), 
	.A(net55579));
   XOR2_X1 U920 (.Z(SUM[36]), 
	.B(net55817), 
	.A(net55583));
   XOR2_X1 U921 (.Z(SUM[37]), 
	.B(net55672), 
	.A(net55587));
   XOR2_X1 U922 (.Z(n395), 
	.B(B[26]), 
	.A(A[26]));
   XOR2_X1 U923 (.Z(SUM[26]), 
	.B(n302), 
	.A(n395));
   NAND2_X1 U924 (.ZN(net55592), 
	.A2(B[26]), 
	.A1(A[26]));
   XOR2_X1 U925 (.Z(SUM[27]), 
	.B(n207), 
	.A(net55595));
   XOR2_X1 U926 (.Z(SUM[16]), 
	.B(net55976), 
	.A(net55599));
   XOR2_X1 U927 (.Z(SUM[17]), 
	.B(n60), 
	.A(net55603));
   XOR2_X1 U928 (.Z(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module up_island (
	CLK, 
	reset, 
	BUS_NREADY, 
	BUS_BUSY, 
	BUS_MR, 
	BUS_MW, 
	BUS_ADDR_OUTBUS, 
	BUS_DATA_INBUS, 
	BUS_DATA_OUTBUS);
   input CLK;
   input reset;
   input BUS_NREADY;
   output BUS_BUSY;
   output BUS_MR;
   output BUS_MW;
   output [31:0] BUS_ADDR_OUTBUS;
   input [31:0] BUS_DATA_INBUS;
   output [31:0] BUS_DATA_OUTBUS;

   // Internal wires
   wire FE_OFCN208_FE_OFN7_n312;
   wire FE_OFCN207_n316;
   wire FE_OFCN206_FE_OFN186_n546;
   wire FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_;
   wire FE_OFCN204_FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_;
   wire FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_;
   wire FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_;
   wire FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_;
   wire FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_;
   wire FE_OFCN199_UUT_rs1_addr_3_;
   wire FE_OFCN198_UUT_Mpath_out_regA_2_;
   wire FE_OFN197_n741;
   wire FE_OFN196_n764;
   wire FE_OFN195_n5438;
   wire FE_OFN194_n5429;
   wire FE_OFN193_n5522;
   wire FE_OFN192_n208;
   wire FE_OFN191_n5435;
   wire FE_OFN190_n5447;
   wire FE_OFN189_n5459;
   wire FE_OFN188_n5492;
   wire FE_OFN187_UUT_branch_rega_1_;
   wire FE_OFN186_n546;
   wire FE_OFN185_UUT_Mpath_out_regB_0_;
   wire FE_OFN184_UUT_Mpath_out_regB_0_;
   wire FE_OFN182_UUT_Mpath_out_regB_0_;
   wire FE_OFN177_UUT_Mpath_the_mult_x_operand1_31_;
   wire FE_OFN176_UUT_Mpath_out_regB_1_;
   wire FE_OFN175_UUT_Mpath_out_regB_1_;
   wire FE_OFN173_UUT_Mpath_the_mult_x_operand1_23_;
   wire FE_OFN171_UUT_Mpath_the_mult_x_operand1_1_;
   wire FE_OFN170_UUT_Mpath_the_mult_x_operand2_1_;
   wire FE_OFN169_UUT_Mpath_out_regB_2_;
   wire FE_OFN168_UUT_Mpath_out_regB_2_;
   wire FE_OFN167_UUT_Mpath_the_mult_x_operand2_2_;
   wire FE_OFN165_UUT_Mpath_the_mult_x_operand1_3_;
   wire FE_OFN164_UUT_Mpath_out_regB_3_;
   wire FE_OFN163_UUT_Mpath_out_regB_3_;
   wire FE_OFN162_UUT_Mpath_out_regB_3_;
   wire FE_OFN160_UUT_Mpath_out_regB_4_;
   wire FE_OFN159_UUT_Mpath_out_regB_4_;
   wire FE_OFN156_UUT_Mpath_the_mult_x_operand1_5_;
   wire FE_OFN152_UUT_Mpath_the_mult_x_operand1_7_;
   wire FE_OFN149_UUT_Mpath_the_mult_x_operand1_9_;
   wire FE_OFN146_UUT_Mpath_the_mult_x_operand1_11_;
   wire FE_OFN142_UUT_Mpath_the_mult_x_operand1_13_;
   wire FE_OFN140_UUT_Mpath_the_mult_x_operand2_14_;
   wire FE_OFN138_UUT_Mpath_the_mult_x_operand1_15_;
   wire FE_OFN137_UUT_Mpath_the_mult_x_operand2_15_;
   wire FE_OFN136_UUT_Mpath_the_mult_x_operand2_16_;
   wire FE_OFN134_UUT_Mpath_the_mult_x_operand1_17_;
   wire FE_OFN133_UUT_Mpath_the_mult_x_operand2_17_;
   wire FE_OFN130_UUT_Mpath_the_mult_x_operand1_19_;
   wire FE_OFN129_UUT_Mpath_the_mult_x_operand2_19_;
   wire FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_;
   wire FE_OFN121_UUT_Mpath_the_mult_x_operand1_25_;
   wire FE_OFN120_UUT_Mpath_the_mult_x_operand2_25_;
   wire FE_OFN117_UUT_Mpath_the_mult_x_operand1_27_;
   wire FE_OFN113_UUT_Mpath_the_mult_x_operand1_29_;
   wire FE_OFN105_UUT_Mpath_the_mult_x_operand2_0_;
   wire FE_OFN104_UUT_Mpath_out_regA_0_;
   wire FE_OFN103_UUT_Mcontrol_Nextpc_decoding_N255;
   wire FE_OFN102_n117;
   wire FE_OFN101_n292;
   wire FE_OFN100_n327;
   wire FE_OFN99_n348;
   wire FE_OFN98_UUT_rs1_addr_1_;
   wire FE_OFN97_n5529;
   wire FE_OFN96_n5530;
   wire FE_OFN95_n2409;
   wire FE_OFN94_n2455;
   wire FE_OFN93_n1878;
   wire FE_OFN92_n5780;
   wire FE_OFN91_n285;
   wire FE_OFN90_n325;
   wire FE_OFN89_n290;
   wire FE_OFN88_n6201;
   wire FE_OFN87_n1211;
   wire FE_OFN86_n1214;
   wire FE_OFN85_n2173;
   wire FE_OFN84_n1498;
   wire FE_OFN83_n2340;
   wire FE_OFN82_n1718;
   wire FE_OFN80_n2581;
   wire FE_OFN79_n1778;
   wire FE_OFN77_n2547;
   wire FE_OFN76_n1798;
   wire FE_OFN74_n2525;
   wire FE_OFN73_n1818;
   wire FE_OFN71_n2501;
   wire FE_OFN69_n2478;
   wire FE_OFN68_n1858;
   wire FE_OFN63_n2386;
   wire FE_OFN62_n1318;
   wire FE_OFN60_n2363;
   wire FE_OFN59_n1338;
   wire FE_OFN57_n2313;
   wire FE_OFN56_n1358;
   wire FE_OFN54_n2293;
   wire FE_OFN53_n1378;
   wire FE_OFN50_n2253;
   wire FE_OFN49_n1418;
   wire FE_OFN30_n5450;
   wire FE_OFN26_n180;
   wire FE_OFN25_n859;
   wire FE_OFN24_n128;
   wire FE_OFN23_n152;
   wire FE_OFN22_n164;
   wire FE_OFN21_n193;
   wire FE_OFN18_n5441;
   wire FE_OFN17_n5444;
   wire FE_OFN13_n953;
   wire FE_OFN12_net54953;
   wire FE_OFN11_net54953;
   wire FE_OFN10_net54953;
   wire FE_OFN9_n986;
   wire FE_OFN8_n73;
   wire FE_OFN7_n312;
   wire FE_OFN6_n314;
   wire FE_OFN5_n318;
   wire FE_OFN4_n319;
   wire FE_OFN3_n202;
   wire FE_OFN1_n189;
   wire FE_OFN0_n173;
   wire FE_UNCONNECTED_1;
   wire FE_UNCONNECTED_0;
   wire I_BUSY;
   wire dmem_read;
   wire dmem_write;
   wire dmem_isbyte;
   wire dmem_ishalf;
   wire dram_mr;
   wire dram_mw;
   wire iram_rd;
   wire N22;
   wire N27;
   wire N31;
   wire N35;
   wire N42;
   wire N43;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N174;
   wire N178;
   wire \UUT/m_mem_command[SIGN] ;
   wire \UUT/m_mem_command[MR] ;
   wire \UUT/m_we ;
   wire \UUT/x_we ;
   wire \UUT/Alu_command[OP][0] ;
   wire \UUT/Alu_command[OP][1] ;
   wire \UUT/Alu_command[OP][2] ;
   wire \UUT/Alu_command[OP][3] ;
   wire \UUT/Alu_command[OP][4] ;
   wire \UUT/Alu_command[OP][5] ;
   wire \UUT/byp_controlB[0] ;
   wire \UUT/byp_controlB[2] ;
   wire \UUT/byp_controlA[0] ;
   wire \UUT/byp_controlA[2] ;
   wire \UUT/break_code[0] ;
   wire \UUT/break_code[1] ;
   wire \UUT/break_code[2] ;
   wire \UUT/break_code[3] ;
   wire \UUT/break_code[4] ;
   wire \UUT/break_code[5] ;
   wire \UUT/break_code[6] ;
   wire \UUT/break_code[7] ;
   wire \UUT/break_code[8] ;
   wire \UUT/break_code[9] ;
   wire \UUT/break_code[10] ;
   wire \UUT/break_code[11] ;
   wire \UUT/break_code[12] ;
   wire \UUT/break_code[13] ;
   wire \UUT/break_code[14] ;
   wire \UUT/break_code[15] ;
   wire \UUT/break_code[16] ;
   wire \UUT/break_code[17] ;
   wire \UUT/break_code[18] ;
   wire \UUT/break_code[19] ;
   wire \UUT/break_code[20] ;
   wire \UUT/break_code[21] ;
   wire \UUT/break_code[22] ;
   wire \UUT/break_code[23] ;
   wire \UUT/N3 ;
   wire \UUT/regfile/N455 ;
   wire \UUT/regfile/N439 ;
   wire \UUT/regfile/N415 ;
   wire \UUT/regfile/N414 ;
   wire \UUT/regfile/N391 ;
   wire \UUT/regfile/N367 ;
   wire \UUT/regfile/N366 ;
   wire \UUT/regfile/N358 ;
   wire \UUT/regfile/N342 ;
   wire \UUT/regfile/N318 ;
   wire \UUT/regfile/N317 ;
   wire \UUT/regfile/N315 ;
   wire \UUT/regfile/N293 ;
   wire \UUT/regfile/N290 ;
   wire \UUT/regfile/N273 ;
   wire \UUT/regfile/N272 ;
   wire \UUT/regfile/N269 ;
   wire \UUT/regfile/N267 ;
   wire \UUT/regfile/N266 ;
   wire \UUT/regfile/N265 ;
   wire \UUT/regfile/N262 ;
   wire \UUT/regfile/N261 ;
   wire \UUT/regfile/N260 ;
   wire \UUT/regfile/reg_out[18][0] ;
   wire \UUT/regfile/reg_out[18][1] ;
   wire \UUT/regfile/reg_out[18][2] ;
   wire \UUT/regfile/reg_out[18][3] ;
   wire \UUT/regfile/reg_out[18][4] ;
   wire \UUT/regfile/reg_out[18][5] ;
   wire \UUT/regfile/reg_out[18][6] ;
   wire \UUT/regfile/reg_out[18][7] ;
   wire \UUT/regfile/reg_out[18][8] ;
   wire \UUT/regfile/reg_out[18][9] ;
   wire \UUT/regfile/reg_out[18][10] ;
   wire \UUT/regfile/reg_out[18][11] ;
   wire \UUT/regfile/reg_out[18][12] ;
   wire \UUT/regfile/reg_out[18][13] ;
   wire \UUT/regfile/reg_out[18][14] ;
   wire \UUT/regfile/reg_out[18][15] ;
   wire \UUT/regfile/reg_out[18][16] ;
   wire \UUT/regfile/reg_out[18][17] ;
   wire \UUT/regfile/reg_out[18][18] ;
   wire \UUT/regfile/reg_out[18][19] ;
   wire \UUT/regfile/reg_out[18][20] ;
   wire \UUT/regfile/reg_out[18][21] ;
   wire \UUT/regfile/reg_out[18][22] ;
   wire \UUT/regfile/reg_out[18][23] ;
   wire \UUT/regfile/reg_out[18][24] ;
   wire \UUT/regfile/reg_out[18][25] ;
   wire \UUT/regfile/reg_out[18][26] ;
   wire \UUT/regfile/reg_out[18][27] ;
   wire \UUT/regfile/reg_out[18][28] ;
   wire \UUT/regfile/reg_out[18][29] ;
   wire \UUT/regfile/reg_out[18][30] ;
   wire \UUT/regfile/reg_out[18][31] ;
   wire \UUT/regfile/reg_out[19][0] ;
   wire \UUT/regfile/reg_out[19][1] ;
   wire \UUT/regfile/reg_out[19][2] ;
   wire \UUT/regfile/reg_out[19][3] ;
   wire \UUT/regfile/reg_out[19][4] ;
   wire \UUT/regfile/reg_out[19][5] ;
   wire \UUT/regfile/reg_out[19][6] ;
   wire \UUT/regfile/reg_out[19][7] ;
   wire \UUT/regfile/reg_out[19][8] ;
   wire \UUT/regfile/reg_out[19][9] ;
   wire \UUT/regfile/reg_out[19][10] ;
   wire \UUT/regfile/reg_out[19][11] ;
   wire \UUT/regfile/reg_out[19][12] ;
   wire \UUT/regfile/reg_out[19][13] ;
   wire \UUT/regfile/reg_out[19][14] ;
   wire \UUT/regfile/reg_out[19][15] ;
   wire \UUT/regfile/reg_out[19][16] ;
   wire \UUT/regfile/reg_out[19][17] ;
   wire \UUT/regfile/reg_out[19][18] ;
   wire \UUT/regfile/reg_out[19][19] ;
   wire \UUT/regfile/reg_out[19][20] ;
   wire \UUT/regfile/reg_out[19][21] ;
   wire \UUT/regfile/reg_out[19][22] ;
   wire \UUT/regfile/reg_out[19][23] ;
   wire \UUT/regfile/reg_out[19][24] ;
   wire \UUT/regfile/reg_out[19][25] ;
   wire \UUT/regfile/reg_out[19][26] ;
   wire \UUT/regfile/reg_out[19][27] ;
   wire \UUT/regfile/reg_out[19][28] ;
   wire \UUT/regfile/reg_out[19][29] ;
   wire \UUT/regfile/reg_out[19][30] ;
   wire \UUT/regfile/reg_out[19][31] ;
   wire \UUT/regfile/reg_out[20][0] ;
   wire \UUT/regfile/reg_out[20][1] ;
   wire \UUT/regfile/reg_out[20][2] ;
   wire \UUT/regfile/reg_out[20][3] ;
   wire \UUT/regfile/reg_out[20][4] ;
   wire \UUT/regfile/reg_out[20][5] ;
   wire \UUT/regfile/reg_out[20][6] ;
   wire \UUT/regfile/reg_out[20][7] ;
   wire \UUT/regfile/reg_out[20][8] ;
   wire \UUT/regfile/reg_out[20][9] ;
   wire \UUT/regfile/reg_out[20][10] ;
   wire \UUT/regfile/reg_out[20][11] ;
   wire \UUT/regfile/reg_out[20][12] ;
   wire \UUT/regfile/reg_out[20][13] ;
   wire \UUT/regfile/reg_out[20][14] ;
   wire \UUT/regfile/reg_out[20][15] ;
   wire \UUT/regfile/reg_out[20][16] ;
   wire \UUT/regfile/reg_out[20][17] ;
   wire \UUT/regfile/reg_out[20][18] ;
   wire \UUT/regfile/reg_out[20][19] ;
   wire \UUT/regfile/reg_out[20][20] ;
   wire \UUT/regfile/reg_out[20][21] ;
   wire \UUT/regfile/reg_out[20][22] ;
   wire \UUT/regfile/reg_out[20][23] ;
   wire \UUT/regfile/reg_out[20][24] ;
   wire \UUT/regfile/reg_out[20][25] ;
   wire \UUT/regfile/reg_out[20][26] ;
   wire \UUT/regfile/reg_out[20][27] ;
   wire \UUT/regfile/reg_out[20][28] ;
   wire \UUT/regfile/reg_out[20][29] ;
   wire \UUT/regfile/reg_out[20][30] ;
   wire \UUT/regfile/reg_out[20][31] ;
   wire \UUT/regfile/reg_out[21][0] ;
   wire \UUT/regfile/reg_out[21][1] ;
   wire \UUT/regfile/reg_out[21][2] ;
   wire \UUT/regfile/reg_out[21][3] ;
   wire \UUT/regfile/reg_out[21][4] ;
   wire \UUT/regfile/reg_out[21][5] ;
   wire \UUT/regfile/reg_out[21][6] ;
   wire \UUT/regfile/reg_out[21][7] ;
   wire \UUT/regfile/reg_out[21][8] ;
   wire \UUT/regfile/reg_out[21][9] ;
   wire \UUT/regfile/reg_out[21][10] ;
   wire \UUT/regfile/reg_out[21][11] ;
   wire \UUT/regfile/reg_out[21][12] ;
   wire \UUT/regfile/reg_out[21][13] ;
   wire \UUT/regfile/reg_out[21][14] ;
   wire \UUT/regfile/reg_out[21][15] ;
   wire \UUT/regfile/reg_out[21][16] ;
   wire \UUT/regfile/reg_out[21][17] ;
   wire \UUT/regfile/reg_out[21][18] ;
   wire \UUT/regfile/reg_out[21][19] ;
   wire \UUT/regfile/reg_out[21][20] ;
   wire \UUT/regfile/reg_out[21][21] ;
   wire \UUT/regfile/reg_out[21][22] ;
   wire \UUT/regfile/reg_out[21][23] ;
   wire \UUT/regfile/reg_out[21][24] ;
   wire \UUT/regfile/reg_out[21][25] ;
   wire \UUT/regfile/reg_out[21][26] ;
   wire \UUT/regfile/reg_out[21][27] ;
   wire \UUT/regfile/reg_out[21][28] ;
   wire \UUT/regfile/reg_out[21][29] ;
   wire \UUT/regfile/reg_out[21][30] ;
   wire \UUT/regfile/reg_out[21][31] ;
   wire \UUT/regfile/reg_out[24][0] ;
   wire \UUT/regfile/reg_out[24][1] ;
   wire \UUT/regfile/reg_out[24][2] ;
   wire \UUT/regfile/reg_out[24][3] ;
   wire \UUT/regfile/reg_out[24][4] ;
   wire \UUT/regfile/reg_out[24][5] ;
   wire \UUT/regfile/reg_out[24][6] ;
   wire \UUT/regfile/reg_out[24][7] ;
   wire \UUT/regfile/reg_out[24][8] ;
   wire \UUT/regfile/reg_out[24][9] ;
   wire \UUT/regfile/reg_out[24][10] ;
   wire \UUT/regfile/reg_out[24][11] ;
   wire \UUT/regfile/reg_out[24][12] ;
   wire \UUT/regfile/reg_out[24][13] ;
   wire \UUT/regfile/reg_out[24][14] ;
   wire \UUT/regfile/reg_out[24][15] ;
   wire \UUT/regfile/reg_out[24][16] ;
   wire \UUT/regfile/reg_out[24][17] ;
   wire \UUT/regfile/reg_out[24][18] ;
   wire \UUT/regfile/reg_out[24][19] ;
   wire \UUT/regfile/reg_out[24][20] ;
   wire \UUT/regfile/reg_out[24][21] ;
   wire \UUT/regfile/reg_out[24][22] ;
   wire \UUT/regfile/reg_out[24][23] ;
   wire \UUT/regfile/reg_out[24][24] ;
   wire \UUT/regfile/reg_out[24][25] ;
   wire \UUT/regfile/reg_out[24][26] ;
   wire \UUT/regfile/reg_out[24][27] ;
   wire \UUT/regfile/reg_out[24][28] ;
   wire \UUT/regfile/reg_out[24][29] ;
   wire \UUT/regfile/reg_out[24][30] ;
   wire \UUT/regfile/reg_out[24][31] ;
   wire \UUT/regfile/reg_out[25][0] ;
   wire \UUT/regfile/reg_out[25][1] ;
   wire \UUT/regfile/reg_out[25][2] ;
   wire \UUT/regfile/reg_out[25][3] ;
   wire \UUT/regfile/reg_out[25][4] ;
   wire \UUT/regfile/reg_out[25][5] ;
   wire \UUT/regfile/reg_out[25][6] ;
   wire \UUT/regfile/reg_out[25][7] ;
   wire \UUT/regfile/reg_out[25][8] ;
   wire \UUT/regfile/reg_out[25][9] ;
   wire \UUT/regfile/reg_out[25][10] ;
   wire \UUT/regfile/reg_out[25][11] ;
   wire \UUT/regfile/reg_out[25][12] ;
   wire \UUT/regfile/reg_out[25][13] ;
   wire \UUT/regfile/reg_out[25][14] ;
   wire \UUT/regfile/reg_out[25][15] ;
   wire \UUT/regfile/reg_out[25][16] ;
   wire \UUT/regfile/reg_out[25][17] ;
   wire \UUT/regfile/reg_out[25][18] ;
   wire \UUT/regfile/reg_out[25][19] ;
   wire \UUT/regfile/reg_out[25][20] ;
   wire \UUT/regfile/reg_out[25][21] ;
   wire \UUT/regfile/reg_out[25][22] ;
   wire \UUT/regfile/reg_out[25][23] ;
   wire \UUT/regfile/reg_out[25][24] ;
   wire \UUT/regfile/reg_out[25][25] ;
   wire \UUT/regfile/reg_out[25][26] ;
   wire \UUT/regfile/reg_out[25][27] ;
   wire \UUT/regfile/reg_out[25][28] ;
   wire \UUT/regfile/reg_out[25][29] ;
   wire \UUT/regfile/reg_out[25][30] ;
   wire \UUT/regfile/reg_out[25][31] ;
   wire \UUT/regfile/reg_out[28][0] ;
   wire \UUT/regfile/reg_out[28][1] ;
   wire \UUT/regfile/reg_out[28][2] ;
   wire \UUT/regfile/reg_out[28][3] ;
   wire \UUT/regfile/reg_out[28][4] ;
   wire \UUT/regfile/reg_out[28][5] ;
   wire \UUT/regfile/reg_out[28][6] ;
   wire \UUT/regfile/reg_out[28][7] ;
   wire \UUT/regfile/reg_out[28][8] ;
   wire \UUT/regfile/reg_out[28][9] ;
   wire \UUT/regfile/reg_out[28][10] ;
   wire \UUT/regfile/reg_out[28][11] ;
   wire \UUT/regfile/reg_out[28][12] ;
   wire \UUT/regfile/reg_out[28][13] ;
   wire \UUT/regfile/reg_out[28][14] ;
   wire \UUT/regfile/reg_out[28][15] ;
   wire \UUT/regfile/reg_out[28][16] ;
   wire \UUT/regfile/reg_out[28][17] ;
   wire \UUT/regfile/reg_out[28][18] ;
   wire \UUT/regfile/reg_out[28][19] ;
   wire \UUT/regfile/reg_out[28][20] ;
   wire \UUT/regfile/reg_out[28][21] ;
   wire \UUT/regfile/reg_out[28][22] ;
   wire \UUT/regfile/reg_out[28][23] ;
   wire \UUT/regfile/reg_out[28][24] ;
   wire \UUT/regfile/reg_out[28][25] ;
   wire \UUT/regfile/reg_out[28][26] ;
   wire \UUT/regfile/reg_out[28][27] ;
   wire \UUT/regfile/reg_out[28][28] ;
   wire \UUT/regfile/reg_out[28][29] ;
   wire \UUT/regfile/reg_out[28][30] ;
   wire \UUT/regfile/reg_out[28][31] ;
   wire \UUT/regfile/reg_out[29][0] ;
   wire \UUT/regfile/reg_out[29][1] ;
   wire \UUT/regfile/reg_out[29][2] ;
   wire \UUT/regfile/reg_out[29][3] ;
   wire \UUT/regfile/reg_out[29][4] ;
   wire \UUT/regfile/reg_out[29][5] ;
   wire \UUT/regfile/reg_out[29][6] ;
   wire \UUT/regfile/reg_out[29][7] ;
   wire \UUT/regfile/reg_out[29][8] ;
   wire \UUT/regfile/reg_out[29][9] ;
   wire \UUT/regfile/reg_out[29][10] ;
   wire \UUT/regfile/reg_out[29][11] ;
   wire \UUT/regfile/reg_out[29][12] ;
   wire \UUT/regfile/reg_out[29][13] ;
   wire \UUT/regfile/reg_out[29][14] ;
   wire \UUT/regfile/reg_out[29][15] ;
   wire \UUT/regfile/reg_out[29][16] ;
   wire \UUT/regfile/reg_out[29][17] ;
   wire \UUT/regfile/reg_out[29][18] ;
   wire \UUT/regfile/reg_out[29][19] ;
   wire \UUT/regfile/reg_out[29][20] ;
   wire \UUT/regfile/reg_out[29][21] ;
   wire \UUT/regfile/reg_out[29][22] ;
   wire \UUT/regfile/reg_out[29][23] ;
   wire \UUT/regfile/reg_out[29][24] ;
   wire \UUT/regfile/reg_out[29][25] ;
   wire \UUT/regfile/reg_out[29][26] ;
   wire \UUT/regfile/reg_out[29][27] ;
   wire \UUT/regfile/reg_out[29][28] ;
   wire \UUT/regfile/reg_out[29][29] ;
   wire \UUT/regfile/reg_out[29][30] ;
   wire \UUT/regfile/reg_out[29][31] ;
   wire \UUT/regfile/reg_out[4][0] ;
   wire \UUT/regfile/reg_out[4][1] ;
   wire \UUT/regfile/reg_out[4][2] ;
   wire \UUT/regfile/reg_out[4][3] ;
   wire \UUT/regfile/reg_out[4][4] ;
   wire \UUT/regfile/reg_out[4][5] ;
   wire \UUT/regfile/reg_out[4][6] ;
   wire \UUT/regfile/reg_out[4][7] ;
   wire \UUT/regfile/reg_out[4][8] ;
   wire \UUT/regfile/reg_out[4][9] ;
   wire \UUT/regfile/reg_out[4][10] ;
   wire \UUT/regfile/reg_out[4][11] ;
   wire \UUT/regfile/reg_out[4][12] ;
   wire \UUT/regfile/reg_out[4][13] ;
   wire \UUT/regfile/reg_out[4][14] ;
   wire \UUT/regfile/reg_out[4][15] ;
   wire \UUT/regfile/reg_out[4][16] ;
   wire \UUT/regfile/reg_out[4][17] ;
   wire \UUT/regfile/reg_out[4][18] ;
   wire \UUT/regfile/reg_out[4][19] ;
   wire \UUT/regfile/reg_out[4][20] ;
   wire \UUT/regfile/reg_out[4][21] ;
   wire \UUT/regfile/reg_out[4][22] ;
   wire \UUT/regfile/reg_out[4][23] ;
   wire \UUT/regfile/reg_out[4][24] ;
   wire \UUT/regfile/reg_out[4][25] ;
   wire \UUT/regfile/reg_out[4][26] ;
   wire \UUT/regfile/reg_out[4][27] ;
   wire \UUT/regfile/reg_out[4][28] ;
   wire \UUT/regfile/reg_out[4][29] ;
   wire \UUT/regfile/reg_out[4][30] ;
   wire \UUT/regfile/reg_out[4][31] ;
   wire \UUT/regfile/reg_out[5][0] ;
   wire \UUT/regfile/reg_out[5][1] ;
   wire \UUT/regfile/reg_out[5][2] ;
   wire \UUT/regfile/reg_out[5][3] ;
   wire \UUT/regfile/reg_out[5][4] ;
   wire \UUT/regfile/reg_out[5][5] ;
   wire \UUT/regfile/reg_out[5][6] ;
   wire \UUT/regfile/reg_out[5][7] ;
   wire \UUT/regfile/reg_out[5][8] ;
   wire \UUT/regfile/reg_out[5][9] ;
   wire \UUT/regfile/reg_out[5][10] ;
   wire \UUT/regfile/reg_out[5][11] ;
   wire \UUT/regfile/reg_out[5][12] ;
   wire \UUT/regfile/reg_out[5][13] ;
   wire \UUT/regfile/reg_out[5][14] ;
   wire \UUT/regfile/reg_out[5][15] ;
   wire \UUT/regfile/reg_out[5][16] ;
   wire \UUT/regfile/reg_out[5][17] ;
   wire \UUT/regfile/reg_out[5][18] ;
   wire \UUT/regfile/reg_out[5][19] ;
   wire \UUT/regfile/reg_out[5][20] ;
   wire \UUT/regfile/reg_out[5][21] ;
   wire \UUT/regfile/reg_out[5][22] ;
   wire \UUT/regfile/reg_out[5][23] ;
   wire \UUT/regfile/reg_out[5][24] ;
   wire \UUT/regfile/reg_out[5][25] ;
   wire \UUT/regfile/reg_out[5][26] ;
   wire \UUT/regfile/reg_out[5][27] ;
   wire \UUT/regfile/reg_out[5][28] ;
   wire \UUT/regfile/reg_out[5][29] ;
   wire \UUT/regfile/reg_out[5][30] ;
   wire \UUT/regfile/reg_out[5][31] ;
   wire \UUT/Mcontrol/x_sampled_dmem_command[SIGN] ;
   wire \UUT/Mcontrol/x_sampled_dmem_command[MW] ;
   wire \UUT/Mcontrol/x_sampled_dmem_command[MR] ;
   wire \UUT/Mcontrol/x_sampled_dmem_command[MH] ;
   wire \UUT/Mcontrol/x_sampled_dmem_command[MB] ;
   wire \UUT/Mcontrol/m_sampled_xrd[0] ;
   wire \UUT/Mcontrol/m_sampled_xrd[1] ;
   wire \UUT/Mcontrol/m_sampled_xrd[2] ;
   wire \UUT/Mcontrol/m_sampled_xrd[3] ;
   wire \UUT/Mcontrol/m_sampled_xrd[4] ;
   wire \UUT/Mcontrol/x_rd[0] ;
   wire \UUT/Mcontrol/x_rd[1] ;
   wire \UUT/Mcontrol/x_rd[2] ;
   wire \UUT/Mcontrol/x_rd[3] ;
   wire \UUT/Mcontrol/x_rd[4] ;
   wire \UUT/Mcontrol/d_jump_type[0] ;
   wire \UUT/Mcontrol/d_jump_type[1] ;
   wire \UUT/Mcontrol/d_jump_type[2] ;
   wire \UUT/Mcontrol/d_jump_type[3] ;
   wire \UUT/Mcontrol/int_reset ;
   wire \UUT/Mcontrol/Program_counter/N24 ;
   wire \UUT/Mcontrol/Program_counter/N22 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2086 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2085 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2084 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2083 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2079 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2071 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2070 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2066 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2061 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2060 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2059 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2054 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2047 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2046 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2045 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2043 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2041 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2040 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2039 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2037 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2036 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2030 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2029 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2025 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2023 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2022 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2020 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2019 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2007 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2005 ;
   wire \UUT/Mcontrol/Operation_decoding32/N2001 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1995 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1994 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1993 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1992 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1991 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1989 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1987 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1981 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1980 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1976 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1975 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1974 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1973 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1972 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1970 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1969 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1964 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1963 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1962 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1958 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1957 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1952 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1951 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1950 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1949 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1948 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1945 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1940 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1939 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1938 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1934 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1933 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1928 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1927 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1926 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1925 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1924 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1923 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1922 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1921 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1915 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1914 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1913 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1912 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1911 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1910 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1909 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1908 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1907 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1906 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1905 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1904 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1903 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1902 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1901 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1900 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1889 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1888 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1887 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1886 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1885 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1884 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1883 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1882 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1881 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1880 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1879 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1877 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1876 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1875 ;
   wire \UUT/Mcontrol/Operation_decoding32/N1871 ;
   wire \UUT/Mcontrol/Operation_decoding32/N89 ;
   wire \UUT/Mcontrol/Operation_decoding32/N62 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N266 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N264 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N262 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N255 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N252 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N247 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N242 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N241 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N224 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N222 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N160 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N159 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N125 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N116 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N114 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N32 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N27 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N25 ;
   wire \UUT/Mcontrol/Nextpc_decoding/N22 ;
   wire \UUT/Mcontrol/bp_logicA/N16 ;
   wire \UUT/Mcontrol/bp_logicA/N15 ;
   wire \UUT/Mcontrol/bp_logicA/N9 ;
   wire \UUT/Mcontrol/bp_logicA/memory_main ;
   wire \UUT/Mcontrol/bp_logicA/N3 ;
   wire \UUT/Mcontrol/bp_logicA/exec_main ;
   wire \UUT/Mcontrol/bp_logicA/N2 ;
   wire \UUT/Mcontrol/bp_logicB/N16 ;
   wire \UUT/Mcontrol/bp_logicB/N15 ;
   wire \UUT/Mcontrol/bp_logicB/N14 ;
   wire \UUT/Mcontrol/bp_logicB/N13 ;
   wire \UUT/Mcontrol/bp_logicB/N12 ;
   wire \UUT/Mcontrol/bp_logicB/N11 ;
   wire \UUT/Mcontrol/bp_logicB/N10 ;
   wire \UUT/Mcontrol/bp_logicB/N9 ;
   wire \UUT/Mcontrol/bp_logicB/N8 ;
   wire \UUT/Mcontrol/bp_logicB/N7 ;
   wire \UUT/Mcontrol/bp_logicB/N6 ;
   wire \UUT/Mcontrol/bp_logicB/N5 ;
   wire \UUT/Mcontrol/bp_logicB/memory_main ;
   wire \UUT/Mcontrol/bp_logicB/N3 ;
   wire \UUT/Mcontrol/bp_logicB/exec_main ;
   wire \UUT/Mcontrol/bp_logicB/N2 ;
   wire \UUT/Mcontrol/st_logic/N120 ;
   wire \UUT/Mcontrol/st_logic/N119 ;
   wire \UUT/Mcontrol/st_logic/N118 ;
   wire \UUT/Mcontrol/st_logic/N117 ;
   wire \UUT/Mcontrol/st_logic/N116 ;
   wire \UUT/Mcontrol/st_logic/N115 ;
   wire \UUT/Mcontrol/st_logic/N114 ;
   wire \UUT/Mcontrol/st_logic/N113 ;
   wire \UUT/Mcontrol/st_logic/N112 ;
   wire \UUT/Mcontrol/st_logic/N111 ;
   wire \UUT/Mcontrol/st_logic/N110 ;
   wire \UUT/Mcontrol/st_logic/N109 ;
   wire \UUT/Mcontrol/st_logic/N106 ;
   wire \UUT/Mcontrol/st_logic/N103 ;
   wire \UUT/Mcontrol/st_logic/N102 ;
   wire \UUT/Mcontrol/st_logic/N101 ;
   wire \UUT/Mcontrol/st_logic/N100 ;
   wire \UUT/Mcontrol/st_logic/N96 ;
   wire \UUT/Mcontrol/st_logic/N95 ;
   wire \UUT/Mcontrol/st_logic/N94 ;
   wire \UUT/Mcontrol/st_logic/N89 ;
   wire \UUT/Mcontrol/st_logic/N88 ;
   wire \UUT/Mcontrol/st_logic/N86 ;
   wire \UUT/Mcontrol/st_logic/N71 ;
   wire \UUT/Mcontrol/st_logic/N70 ;
   wire \UUT/Mcontrol/st_logic/N65 ;
   wire \UUT/Mcontrol/st_logic/N63 ;
   wire \UUT/Mcontrol/st_logic/N61 ;
   wire \UUT/Mcontrol/st_logic/N58 ;
   wire \UUT/Mcontrol/st_logic/N55 ;
   wire \UUT/Mcontrol/st_logic/N52 ;
   wire \UUT/Mcontrol/st_logic/N50 ;
   wire \UUT/Mcontrol/st_logic/N49 ;
   wire \UUT/Mcontrol/st_logic/N47 ;
   wire \UUT/Mcontrol/st_logic/N45 ;
   wire \UUT/Mcontrol/st_logic/N44 ;
   wire \UUT/Mcontrol/st_logic/N42 ;
   wire \UUT/Mcontrol/st_logic/N40 ;
   wire \UUT/Mcontrol/st_logic/N39 ;
   wire \UUT/Mcontrol/st_logic/N34 ;
   wire \UUT/Mcontrol/st_logic/N33 ;
   wire \UUT/Mcontrol/st_logic/N32 ;
   wire \UUT/Mcontrol/st_logic/N31 ;
   wire \UUT/Mcontrol/st_logic/N30 ;
   wire \UUT/Mcontrol/st_logic/N29 ;
   wire \UUT/Mcontrol/st_logic/N28 ;
   wire \UUT/Mcontrol/st_logic/N27 ;
   wire \UUT/Mcontrol/st_logic/N26 ;
   wire \UUT/Mcontrol/st_logic/N24 ;
   wire \UUT/Mcontrol/st_logic/N23 ;
   wire \UUT/Mcontrol/st_logic/N22 ;
   wire \UUT/Mcontrol/st_logic/N19 ;
   wire \UUT/Mcontrol/st_logic/N18 ;
   wire \UUT/Mcontrol/st_logic/N10 ;
   wire \UUT/Mcontrol/st_logic/N8 ;
   wire \UUT/Mcontrol/st_logic/N7 ;
   wire \UUT/Mcontrol/st_logic/N6 ;
   wire \UUT/Mcontrol/st_logic/N5 ;
   wire \UUT/Mcontrol/st_logic/N3 ;
   wire \UUT/Mcontrol/st_logic/N2 ;
   wire \UUT/Mpath/N125 ;
   wire \UUT/Mpath/N124 ;
   wire \UUT/Mpath/N119 ;
   wire \UUT/Mpath/N118 ;
   wire \UUT/Mpath/N117 ;
   wire \UUT/Mpath/N116 ;
   wire \UUT/Mpath/N115 ;
   wire \UUT/Mpath/N114 ;
   wire \UUT/Mpath/N113 ;
   wire \UUT/Mpath/N112 ;
   wire \UUT/Mpath/N111 ;
   wire \UUT/Mpath/out_jar[0] ;
   wire \UUT/Mpath/out_jar[1] ;
   wire \UUT/Mpath/out_jar[2] ;
   wire \UUT/Mpath/out_jar[3] ;
   wire \UUT/Mpath/out_jar[4] ;
   wire \UUT/Mpath/out_jar[5] ;
   wire \UUT/Mpath/out_jar[6] ;
   wire \UUT/Mpath/out_jar[7] ;
   wire \UUT/Mpath/out_jar[8] ;
   wire \UUT/Mpath/out_jar[9] ;
   wire \UUT/Mpath/out_jar[10] ;
   wire \UUT/Mpath/out_jar[11] ;
   wire \UUT/Mpath/out_jar[12] ;
   wire \UUT/Mpath/out_jar[13] ;
   wire \UUT/Mpath/out_jar[14] ;
   wire \UUT/Mpath/out_jar[15] ;
   wire \UUT/Mpath/out_jar[16] ;
   wire \UUT/Mpath/out_jar[17] ;
   wire \UUT/Mpath/out_jar[18] ;
   wire \UUT/Mpath/out_jar[19] ;
   wire \UUT/Mpath/out_jar[20] ;
   wire \UUT/Mpath/out_jar[21] ;
   wire \UUT/Mpath/out_jar[22] ;
   wire \UUT/Mpath/out_jar[23] ;
   wire \UUT/Mpath/out_regB[0] ;
   wire \UUT/Mpath/out_regB[1] ;
   wire \UUT/Mpath/out_regB[2] ;
   wire \UUT/Mpath/out_regB[3] ;
   wire \UUT/Mpath/out_regB[4] ;
   wire \UUT/Mpath/out_regB[5] ;
   wire \UUT/Mpath/out_regB[6] ;
   wire \UUT/Mpath/out_regB[7] ;
   wire \UUT/Mpath/out_regB[8] ;
   wire \UUT/Mpath/out_regB[9] ;
   wire \UUT/Mpath/out_regB[10] ;
   wire \UUT/Mpath/out_regB[11] ;
   wire \UUT/Mpath/out_regB[12] ;
   wire \UUT/Mpath/out_regB[13] ;
   wire \UUT/Mpath/out_regB[14] ;
   wire \UUT/Mpath/out_regB[15] ;
   wire \UUT/Mpath/out_regB[16] ;
   wire \UUT/Mpath/out_regB[17] ;
   wire \UUT/Mpath/out_regB[18] ;
   wire \UUT/Mpath/out_regB[19] ;
   wire \UUT/Mpath/out_regB[20] ;
   wire \UUT/Mpath/out_regB[21] ;
   wire \UUT/Mpath/out_regB[22] ;
   wire \UUT/Mpath/out_regB[23] ;
   wire \UUT/Mpath/out_regB[24] ;
   wire \UUT/Mpath/out_regB[25] ;
   wire \UUT/Mpath/out_regB[26] ;
   wire \UUT/Mpath/out_regB[27] ;
   wire \UUT/Mpath/out_regB[28] ;
   wire \UUT/Mpath/out_regB[29] ;
   wire \UUT/Mpath/out_regB[30] ;
   wire \UUT/Mpath/out_regB[31] ;
   wire \UUT/Mpath/out_regA[0] ;
   wire \UUT/Mpath/out_regA[1] ;
   wire \UUT/Mpath/out_regA[2] ;
   wire \UUT/Mpath/out_regA[3] ;
   wire \UUT/Mpath/out_regA[4] ;
   wire \UUT/Mpath/out_regA[5] ;
   wire \UUT/Mpath/out_regA[6] ;
   wire \UUT/Mpath/out_regA[7] ;
   wire \UUT/Mpath/out_regA[8] ;
   wire \UUT/Mpath/out_regA[9] ;
   wire \UUT/Mpath/out_regA[10] ;
   wire \UUT/Mpath/out_regA[11] ;
   wire \UUT/Mpath/out_regA[12] ;
   wire \UUT/Mpath/out_regA[13] ;
   wire \UUT/Mpath/out_regA[14] ;
   wire \UUT/Mpath/out_regA[15] ;
   wire \UUT/Mpath/out_regA[16] ;
   wire \UUT/Mpath/out_regA[17] ;
   wire \UUT/Mpath/out_regA[18] ;
   wire \UUT/Mpath/out_regA[19] ;
   wire \UUT/Mpath/out_regA[20] ;
   wire \UUT/Mpath/out_regA[21] ;
   wire \UUT/Mpath/out_regA[22] ;
   wire \UUT/Mpath/out_regA[23] ;
   wire \UUT/Mpath/out_regA[24] ;
   wire \UUT/Mpath/out_regA[25] ;
   wire \UUT/Mpath/out_regA[26] ;
   wire \UUT/Mpath/out_regA[27] ;
   wire \UUT/Mpath/out_regA[28] ;
   wire \UUT/Mpath/out_regA[29] ;
   wire \UUT/Mpath/out_regA[30] ;
   wire \UUT/Mpath/out_regA[31] ;
   wire \UUT/Mpath/the_alu/N520 ;
   wire \UUT/Mpath/the_alu/N519 ;
   wire \UUT/Mpath/the_alu/N518 ;
   wire \UUT/Mpath/the_alu/N517 ;
   wire \UUT/Mpath/the_alu/N515 ;
   wire \UUT/Mpath/the_alu/N509 ;
   wire \UUT/Mpath/the_alu/N508 ;
   wire \UUT/Mpath/the_alu/N507 ;
   wire \UUT/Mpath/the_alu/N506 ;
   wire \UUT/Mpath/the_alu/N505 ;
   wire \UUT/Mpath/the_alu/N503 ;
   wire \UUT/Mpath/the_alu/N498 ;
   wire \UUT/Mpath/the_alu/N497 ;
   wire \UUT/Mpath/the_alu/N496 ;
   wire \UUT/Mpath/the_alu/N495 ;
   wire \UUT/Mpath/the_alu/N494 ;
   wire \UUT/Mpath/the_alu/N493 ;
   wire \UUT/Mpath/the_alu/N492 ;
   wire \UUT/Mpath/the_alu/N491 ;
   wire \UUT/Mpath/the_alu/N486 ;
   wire \UUT/Mpath/the_alu/N485 ;
   wire \UUT/Mpath/the_alu/N484 ;
   wire \UUT/Mpath/the_alu/N480 ;
   wire \UUT/Mpath/the_alu/N479 ;
   wire \UUT/Mpath/the_alu/N474 ;
   wire \UUT/Mpath/the_alu/N473 ;
   wire \UUT/Mpath/the_alu/N472 ;
   wire \UUT/Mpath/the_alu/N471 ;
   wire \UUT/Mpath/the_alu/N470 ;
   wire \UUT/Mpath/the_alu/N469 ;
   wire \UUT/Mpath/the_alu/N468 ;
   wire \UUT/Mpath/the_alu/N467 ;
   wire \UUT/Mpath/the_alu/N466 ;
   wire \UUT/Mpath/the_alu/N453 ;
   wire \UUT/Mpath/the_alu/N221 ;
   wire \UUT/Mpath/the_alu/N219 ;
   wire \UUT/Mpath/the_alu/N218 ;
   wire \UUT/Mpath/the_alu/N217 ;
   wire \UUT/Mpath/the_alu/N216 ;
   wire \UUT/Mpath/the_alu/N215 ;
   wire \UUT/Mpath/the_alu/N214 ;
   wire \UUT/Mpath/the_alu/N213 ;
   wire \UUT/Mpath/the_alu/N212 ;
   wire \UUT/Mpath/the_alu/N211 ;
   wire \UUT/Mpath/the_alu/N210 ;
   wire \UUT/Mpath/the_alu/N209 ;
   wire \UUT/Mpath/the_alu/N208 ;
   wire \UUT/Mpath/the_alu/N207 ;
   wire \UUT/Mpath/the_alu/N206 ;
   wire \UUT/Mpath/the_alu/N205 ;
   wire \UUT/Mpath/the_alu/N204 ;
   wire \UUT/Mpath/the_alu/N203 ;
   wire \UUT/Mpath/the_alu/N202 ;
   wire \UUT/Mpath/the_alu/N201 ;
   wire \UUT/Mpath/the_alu/N200 ;
   wire \UUT/Mpath/the_alu/N199 ;
   wire \UUT/Mpath/the_alu/N198 ;
   wire \UUT/Mpath/the_alu/N197 ;
   wire \UUT/Mpath/the_alu/N196 ;
   wire \UUT/Mpath/the_alu/N195 ;
   wire \UUT/Mpath/the_alu/N194 ;
   wire \UUT/Mpath/the_alu/N193 ;
   wire \UUT/Mpath/the_alu/N192 ;
   wire \UUT/Mpath/the_alu/N191 ;
   wire \UUT/Mpath/the_alu/N190 ;
   wire \UUT/Mpath/the_alu/N189 ;
   wire \UUT/Mpath/the_alu/N187 ;
   wire \UUT/Mpath/the_alu/N186 ;
   wire \UUT/Mpath/the_alu/N185 ;
   wire \UUT/Mpath/the_alu/N184 ;
   wire \UUT/Mpath/the_alu/N183 ;
   wire \UUT/Mpath/the_alu/N182 ;
   wire \UUT/Mpath/the_alu/N181 ;
   wire \UUT/Mpath/the_alu/N180 ;
   wire \UUT/Mpath/the_alu/N179 ;
   wire \UUT/Mpath/the_alu/N178 ;
   wire \UUT/Mpath/the_alu/N177 ;
   wire \UUT/Mpath/the_alu/N176 ;
   wire \UUT/Mpath/the_alu/N175 ;
   wire \UUT/Mpath/the_alu/N174 ;
   wire \UUT/Mpath/the_alu/N173 ;
   wire \UUT/Mpath/the_alu/N172 ;
   wire \UUT/Mpath/the_alu/N171 ;
   wire \UUT/Mpath/the_alu/N170 ;
   wire \UUT/Mpath/the_alu/N169 ;
   wire \UUT/Mpath/the_alu/N168 ;
   wire \UUT/Mpath/the_alu/N167 ;
   wire \UUT/Mpath/the_alu/N166 ;
   wire \UUT/Mpath/the_alu/N165 ;
   wire \UUT/Mpath/the_alu/N164 ;
   wire \UUT/Mpath/the_alu/N163 ;
   wire \UUT/Mpath/the_alu/N162 ;
   wire \UUT/Mpath/the_alu/N161 ;
   wire \UUT/Mpath/the_alu/N160 ;
   wire \UUT/Mpath/the_alu/N159 ;
   wire \UUT/Mpath/the_alu/N158 ;
   wire \UUT/Mpath/the_alu/N157 ;
   wire \UUT/Mpath/the_alu/N155 ;
   wire \UUT/Mpath/the_alu/N154 ;
   wire \UUT/Mpath/the_alu/N153 ;
   wire \UUT/Mpath/the_alu/N152 ;
   wire \UUT/Mpath/the_alu/N151 ;
   wire \UUT/Mpath/the_alu/N150 ;
   wire \UUT/Mpath/the_alu/N149 ;
   wire \UUT/Mpath/the_alu/N148 ;
   wire \UUT/Mpath/the_alu/N147 ;
   wire \UUT/Mpath/the_alu/N146 ;
   wire \UUT/Mpath/the_alu/N145 ;
   wire \UUT/Mpath/the_alu/N144 ;
   wire \UUT/Mpath/the_alu/N143 ;
   wire \UUT/Mpath/the_alu/N142 ;
   wire \UUT/Mpath/the_alu/N141 ;
   wire \UUT/Mpath/the_alu/N140 ;
   wire \UUT/Mpath/the_alu/N139 ;
   wire \UUT/Mpath/the_alu/N138 ;
   wire \UUT/Mpath/the_alu/N137 ;
   wire \UUT/Mpath/the_alu/N136 ;
   wire \UUT/Mpath/the_alu/N135 ;
   wire \UUT/Mpath/the_alu/N134 ;
   wire \UUT/Mpath/the_alu/N133 ;
   wire \UUT/Mpath/the_alu/N132 ;
   wire \UUT/Mpath/the_alu/N131 ;
   wire \UUT/Mpath/the_alu/N130 ;
   wire \UUT/Mpath/the_alu/N129 ;
   wire \UUT/Mpath/the_alu/N128 ;
   wire \UUT/Mpath/the_alu/N127 ;
   wire \UUT/Mpath/the_alu/N126 ;
   wire \UUT/Mpath/the_alu/N125 ;
   wire \UUT/Mpath/the_alu/N123 ;
   wire \UUT/Mpath/the_alu/N122 ;
   wire \UUT/Mpath/the_alu/N121 ;
   wire \UUT/Mpath/the_alu/N120 ;
   wire \UUT/Mpath/the_alu/N119 ;
   wire \UUT/Mpath/the_alu/N118 ;
   wire \UUT/Mpath/the_alu/N117 ;
   wire \UUT/Mpath/the_alu/N116 ;
   wire \UUT/Mpath/the_alu/N115 ;
   wire \UUT/Mpath/the_alu/N114 ;
   wire \UUT/Mpath/the_alu/N113 ;
   wire \UUT/Mpath/the_alu/N112 ;
   wire \UUT/Mpath/the_alu/N111 ;
   wire \UUT/Mpath/the_alu/N110 ;
   wire \UUT/Mpath/the_alu/N109 ;
   wire \UUT/Mpath/the_alu/N108 ;
   wire \UUT/Mpath/the_alu/N107 ;
   wire \UUT/Mpath/the_alu/N106 ;
   wire \UUT/Mpath/the_alu/N105 ;
   wire \UUT/Mpath/the_alu/N104 ;
   wire \UUT/Mpath/the_alu/N103 ;
   wire \UUT/Mpath/the_alu/N102 ;
   wire \UUT/Mpath/the_alu/N101 ;
   wire \UUT/Mpath/the_alu/N100 ;
   wire \UUT/Mpath/the_alu/N99 ;
   wire \UUT/Mpath/the_alu/N98 ;
   wire \UUT/Mpath/the_alu/N97 ;
   wire \UUT/Mpath/the_alu/N96 ;
   wire \UUT/Mpath/the_alu/N95 ;
   wire \UUT/Mpath/the_alu/N94 ;
   wire \UUT/Mpath/the_alu/N93 ;
   wire \UUT/Mpath/the_alu/N91 ;
   wire \UUT/Mpath/the_alu/diff[0] ;
   wire \UUT/Mpath/the_alu/diff[1] ;
   wire \UUT/Mpath/the_alu/diff[2] ;
   wire \UUT/Mpath/the_alu/diff[3] ;
   wire \UUT/Mpath/the_alu/diff[4] ;
   wire \UUT/Mpath/the_alu/diff[5] ;
   wire \UUT/Mpath/the_alu/diff[6] ;
   wire \UUT/Mpath/the_alu/diff[7] ;
   wire \UUT/Mpath/the_alu/diff[8] ;
   wire \UUT/Mpath/the_alu/diff[9] ;
   wire \UUT/Mpath/the_alu/diff[10] ;
   wire \UUT/Mpath/the_alu/diff[11] ;
   wire \UUT/Mpath/the_alu/diff[12] ;
   wire \UUT/Mpath/the_alu/diff[13] ;
   wire \UUT/Mpath/the_alu/diff[14] ;
   wire \UUT/Mpath/the_alu/diff[15] ;
   wire \UUT/Mpath/the_alu/diff[16] ;
   wire \UUT/Mpath/the_alu/diff[17] ;
   wire \UUT/Mpath/the_alu/diff[18] ;
   wire \UUT/Mpath/the_alu/diff[19] ;
   wire \UUT/Mpath/the_alu/diff[20] ;
   wire \UUT/Mpath/the_alu/diff[21] ;
   wire \UUT/Mpath/the_alu/diff[22] ;
   wire \UUT/Mpath/the_alu/diff[23] ;
   wire \UUT/Mpath/the_alu/diff[24] ;
   wire \UUT/Mpath/the_alu/diff[25] ;
   wire \UUT/Mpath/the_alu/diff[26] ;
   wire \UUT/Mpath/the_alu/diff[27] ;
   wire \UUT/Mpath/the_alu/diff[28] ;
   wire \UUT/Mpath/the_alu/diff[29] ;
   wire \UUT/Mpath/the_alu/diff[30] ;
   wire \UUT/Mpath/the_alu/diff[31] ;
   wire \UUT/Mpath/the_alu/sum[0] ;
   wire \UUT/Mpath/the_alu/sum[1] ;
   wire \UUT/Mpath/the_alu/sum[2] ;
   wire \UUT/Mpath/the_alu/sum[3] ;
   wire \UUT/Mpath/the_alu/sum[4] ;
   wire \UUT/Mpath/the_alu/sum[5] ;
   wire \UUT/Mpath/the_alu/sum[6] ;
   wire \UUT/Mpath/the_alu/sum[7] ;
   wire \UUT/Mpath/the_alu/sum[8] ;
   wire \UUT/Mpath/the_alu/sum[9] ;
   wire \UUT/Mpath/the_alu/sum[10] ;
   wire \UUT/Mpath/the_alu/sum[11] ;
   wire \UUT/Mpath/the_alu/sum[12] ;
   wire \UUT/Mpath/the_alu/sum[13] ;
   wire \UUT/Mpath/the_alu/sum[14] ;
   wire \UUT/Mpath/the_alu/sum[15] ;
   wire \UUT/Mpath/the_alu/sum[16] ;
   wire \UUT/Mpath/the_alu/sum[17] ;
   wire \UUT/Mpath/the_alu/sum[18] ;
   wire \UUT/Mpath/the_alu/sum[19] ;
   wire \UUT/Mpath/the_alu/sum[20] ;
   wire \UUT/Mpath/the_alu/sum[21] ;
   wire \UUT/Mpath/the_alu/sum[22] ;
   wire \UUT/Mpath/the_alu/sum[23] ;
   wire \UUT/Mpath/the_alu/sum[24] ;
   wire \UUT/Mpath/the_alu/sum[25] ;
   wire \UUT/Mpath/the_alu/sum[26] ;
   wire \UUT/Mpath/the_alu/sum[27] ;
   wire \UUT/Mpath/the_alu/sum[28] ;
   wire \UUT/Mpath/the_alu/sum[29] ;
   wire \UUT/Mpath/the_alu/sum[30] ;
   wire \UUT/Mpath/the_alu/sum[31] ;
   wire \UUT/Mpath/the_alu/N84 ;
   wire \UUT/Mpath/the_alu/N83 ;
   wire \UUT/Mpath/the_alu/N82 ;
   wire \UUT/Mpath/the_alu/N81 ;
   wire \UUT/Mpath/the_alu/N80 ;
   wire \UUT/Mpath/the_alu/N79 ;
   wire \UUT/Mpath/the_alu/N78 ;
   wire \UUT/Mpath/the_alu/N77 ;
   wire \UUT/Mpath/the_alu/N76 ;
   wire \UUT/Mpath/the_alu/N75 ;
   wire \UUT/Mpath/the_alu/N74 ;
   wire \UUT/Mpath/the_alu/N73 ;
   wire \UUT/Mpath/the_alu/N72 ;
   wire \UUT/Mpath/the_alu/N71 ;
   wire \UUT/Mpath/the_alu/N70 ;
   wire \UUT/Mpath/the_alu/N69 ;
   wire \UUT/Mpath/the_alu/N68 ;
   wire \UUT/Mpath/the_alu/N67 ;
   wire \UUT/Mpath/the_alu/N66 ;
   wire \UUT/Mpath/the_alu/N65 ;
   wire \UUT/Mpath/the_alu/N64 ;
   wire \UUT/Mpath/the_alu/N63 ;
   wire \UUT/Mpath/the_alu/N62 ;
   wire \UUT/Mpath/the_alu/N61 ;
   wire \UUT/Mpath/the_alu/N60 ;
   wire \UUT/Mpath/the_alu/N59 ;
   wire \UUT/Mpath/the_alu/N58 ;
   wire \UUT/Mpath/the_alu/N57 ;
   wire \UUT/Mpath/the_alu/N56 ;
   wire \UUT/Mpath/the_alu/N55 ;
   wire \UUT/Mpath/the_alu/N54 ;
   wire \UUT/Mpath/the_alu/N53 ;
   wire \UUT/Mpath/the_alu/N52 ;
   wire \UUT/Mpath/the_alu/N51 ;
   wire \UUT/Mpath/the_alu/N50 ;
   wire \UUT/Mpath/the_alu/N49 ;
   wire \UUT/Mpath/the_alu/N48 ;
   wire \UUT/Mpath/the_alu/N47 ;
   wire \UUT/Mpath/the_alu/N46 ;
   wire \UUT/Mpath/the_alu/N45 ;
   wire \UUT/Mpath/the_alu/N44 ;
   wire \UUT/Mpath/the_alu/N43 ;
   wire \UUT/Mpath/the_alu/N42 ;
   wire \UUT/Mpath/the_alu/N41 ;
   wire \UUT/Mpath/the_alu/N40 ;
   wire \UUT/Mpath/the_alu/N39 ;
   wire \UUT/Mpath/the_alu/N38 ;
   wire \UUT/Mpath/the_alu/N37 ;
   wire \UUT/Mpath/the_alu/N36 ;
   wire \UUT/Mpath/the_alu/N35 ;
   wire \UUT/Mpath/the_alu/N34 ;
   wire \UUT/Mpath/the_alu/N33 ;
   wire \UUT/Mpath/the_alu/N32 ;
   wire \UUT/Mpath/the_alu/N31 ;
   wire \UUT/Mpath/the_alu/N30 ;
   wire \UUT/Mpath/the_alu/N29 ;
   wire \UUT/Mpath/the_alu/N28 ;
   wire \UUT/Mpath/the_alu/N27 ;
   wire \UUT/Mpath/the_alu/N26 ;
   wire \UUT/Mpath/the_alu/N25 ;
   wire \UUT/Mpath/the_alu/N24 ;
   wire \UUT/Mpath/the_alu/N23 ;
   wire \UUT/Mpath/the_alu/N22 ;
   wire \UUT/Mpath/the_alu/N21 ;
   wire \UUT/Mpath/the_shift/N118 ;
   wire \UUT/Mpath/the_shift/N117 ;
   wire \UUT/Mpath/the_shift/N116 ;
   wire \UUT/Mpath/the_shift/N115 ;
   wire \UUT/Mpath/the_shift/N114 ;
   wire \UUT/Mpath/the_shift/N113 ;
   wire \UUT/Mpath/the_shift/N112 ;
   wire \UUT/Mpath/the_shift/N111 ;
   wire \UUT/Mpath/the_shift/N110 ;
   wire \UUT/Mpath/the_shift/N108 ;
   wire \UUT/Mpath/the_shift/N107 ;
   wire \UUT/Mpath/the_shift/N106 ;
   wire \UUT/Mpath/the_shift/N105 ;
   wire \UUT/Mpath/the_shift/N104 ;
   wire \UUT/Mpath/the_mult/N312 ;
   wire \UUT/Mpath/the_mult/N311 ;
   wire \UUT/Mpath/the_mult/N285 ;
   wire \UUT/Mpath/the_mult/N280 ;
   wire \UUT/Mpath/the_mult/N279 ;
   wire \UUT/Mpath/the_mult/N274 ;
   wire \UUT/Mpath/the_mult/N273 ;
   wire \UUT/Mpath/the_mult/N272 ;
   wire \UUT/Mpath/the_mult/N271 ;
   wire \UUT/Mpath/the_mult/N268 ;
   wire \UUT/Mpath/the_mult/N267 ;
   wire \UUT/Mpath/the_mult/N262 ;
   wire \UUT/Mpath/the_mult/N261 ;
   wire \UUT/Mpath/the_mult/N260 ;
   wire \UUT/Mpath/the_mult/N259 ;
   wire \UUT/Mpath/the_mult/N258 ;
   wire \UUT/Mpath/the_mult/N255 ;
   wire \UUT/Mpath/the_mult/N254 ;
   wire \UUT/Mpath/the_mult/N253 ;
   wire \UUT/Mpath/the_mult/N252 ;
   wire \UUT/Mpath/the_mult/N251 ;
   wire \UUT/Mpath/the_mult/N244 ;
   wire \UUT/Mpath/the_mult/N231 ;
   wire \UUT/Mpath/the_mult/N230 ;
   wire \UUT/Mpath/the_mult/N229 ;
   wire \UUT/Mpath/the_mult/N227 ;
   wire \UUT/Mpath/the_mult/N226 ;
   wire \UUT/Mpath/the_mult/N225 ;
   wire \UUT/Mpath/the_mult/N224 ;
   wire \UUT/Mpath/the_mult/N223 ;
   wire \UUT/Mpath/the_mult/N222 ;
   wire \UUT/Mpath/the_mult/N221 ;
   wire \UUT/Mpath/the_mult/N220 ;
   wire \UUT/Mpath/the_mult/N216 ;
   wire \UUT/Mpath/the_mult/N198 ;
   wire \UUT/Mpath/the_mult/N197 ;
   wire \UUT/Mpath/the_mult/N196 ;
   wire \UUT/Mpath/the_mult/N195 ;
   wire \UUT/Mpath/the_mult/N194 ;
   wire \UUT/Mpath/the_mult/N193 ;
   wire \UUT/Mpath/the_mult/N192 ;
   wire \UUT/Mpath/the_mult/acc_out[0] ;
   wire \UUT/Mpath/the_mult/acc_out[1] ;
   wire \UUT/Mpath/the_mult/acc_out[2] ;
   wire \UUT/Mpath/the_mult/acc_out[3] ;
   wire \UUT/Mpath/the_mult/acc_out[4] ;
   wire \UUT/Mpath/the_mult/acc_out[5] ;
   wire \UUT/Mpath/the_mult/acc_out[6] ;
   wire \UUT/Mpath/the_mult/acc_out[7] ;
   wire \UUT/Mpath/the_mult/acc_out[8] ;
   wire \UUT/Mpath/the_mult/acc_out[9] ;
   wire \UUT/Mpath/the_mult/acc_out[10] ;
   wire \UUT/Mpath/the_mult/acc_out[11] ;
   wire \UUT/Mpath/the_mult/acc_out[12] ;
   wire \UUT/Mpath/the_mult/acc_out[13] ;
   wire \UUT/Mpath/the_mult/acc_out[14] ;
   wire \UUT/Mpath/the_mult/acc_out[15] ;
   wire \UUT/Mpath/the_mult/acc_out[16] ;
   wire \UUT/Mpath/the_mult/acc_out[17] ;
   wire \UUT/Mpath/the_mult/acc_out[18] ;
   wire \UUT/Mpath/the_mult/acc_out[19] ;
   wire \UUT/Mpath/the_mult/acc_out[20] ;
   wire \UUT/Mpath/the_mult/acc_out[21] ;
   wire \UUT/Mpath/the_mult/acc_out[22] ;
   wire \UUT/Mpath/the_mult/acc_out[23] ;
   wire \UUT/Mpath/the_mult/acc_out[24] ;
   wire \UUT/Mpath/the_mult/acc_out[25] ;
   wire \UUT/Mpath/the_mult/acc_out[26] ;
   wire \UUT/Mpath/the_mult/acc_out[27] ;
   wire \UUT/Mpath/the_mult/acc_out[28] ;
   wire \UUT/Mpath/the_mult/acc_out[29] ;
   wire \UUT/Mpath/the_mult/acc_out[30] ;
   wire \UUT/Mpath/the_mult/acc_out[31] ;
   wire \UUT/Mpath/the_mult/acc_out[32] ;
   wire \UUT/Mpath/the_mult/acc_out[33] ;
   wire \UUT/Mpath/the_mult/acc_out[34] ;
   wire \UUT/Mpath/the_mult/acc_out[35] ;
   wire \UUT/Mpath/the_mult/acc_out[36] ;
   wire \UUT/Mpath/the_mult/acc_out[37] ;
   wire \UUT/Mpath/the_mult/acc_out[38] ;
   wire \UUT/Mpath/the_mult/acc_out[39] ;
   wire \UUT/Mpath/the_mult/acc_out[40] ;
   wire \UUT/Mpath/the_mult/acc_out[41] ;
   wire \UUT/Mpath/the_mult/acc_out[42] ;
   wire \UUT/Mpath/the_mult/acc_out[43] ;
   wire \UUT/Mpath/the_mult/acc_out[44] ;
   wire \UUT/Mpath/the_mult/acc_out[45] ;
   wire \UUT/Mpath/the_mult/acc_out[46] ;
   wire \UUT/Mpath/the_mult/acc_out[47] ;
   wire \UUT/Mpath/the_mult/acc_out[48] ;
   wire \UUT/Mpath/the_mult/acc_out[49] ;
   wire \UUT/Mpath/the_mult/acc_out[50] ;
   wire \UUT/Mpath/the_mult/acc_out[51] ;
   wire \UUT/Mpath/the_mult/acc_out[52] ;
   wire \UUT/Mpath/the_mult/acc_out[53] ;
   wire \UUT/Mpath/the_mult/acc_out[54] ;
   wire \UUT/Mpath/the_mult/acc_out[55] ;
   wire \UUT/Mpath/the_mult/acc_out[56] ;
   wire \UUT/Mpath/the_mult/acc_out[57] ;
   wire \UUT/Mpath/the_mult/acc_out[58] ;
   wire \UUT/Mpath/the_mult/acc_out[59] ;
   wire \UUT/Mpath/the_mult/acc_out[60] ;
   wire \UUT/Mpath/the_mult/acc_out[61] ;
   wire \UUT/Mpath/the_mult/acc_out[62] ;
   wire \UUT/Mpath/the_mult/acc_out[63] ;
   wire \UUT/Mpath/the_mult/Mult_out[0] ;
   wire \UUT/Mpath/the_mult/Mult_out[1] ;
   wire \UUT/Mpath/the_mult/Mult_out[2] ;
   wire \UUT/Mpath/the_mult/Mult_out[3] ;
   wire \UUT/Mpath/the_mult/Mult_out[4] ;
   wire \UUT/Mpath/the_mult/Mult_out[5] ;
   wire \UUT/Mpath/the_mult/Mult_out[6] ;
   wire \UUT/Mpath/the_mult/Mult_out[7] ;
   wire \UUT/Mpath/the_mult/Mult_out[8] ;
   wire \UUT/Mpath/the_mult/Mult_out[9] ;
   wire \UUT/Mpath/the_mult/Mult_out[10] ;
   wire \UUT/Mpath/the_mult/Mult_out[11] ;
   wire \UUT/Mpath/the_mult/Mult_out[12] ;
   wire \UUT/Mpath/the_mult/Mult_out[13] ;
   wire \UUT/Mpath/the_mult/Mult_out[14] ;
   wire \UUT/Mpath/the_mult/Mult_out[15] ;
   wire \UUT/Mpath/the_mult/Mult_out[16] ;
   wire \UUT/Mpath/the_mult/Mult_out[17] ;
   wire \UUT/Mpath/the_mult/Mult_out[18] ;
   wire \UUT/Mpath/the_mult/Mult_out[19] ;
   wire \UUT/Mpath/the_mult/Mult_out[20] ;
   wire \UUT/Mpath/the_mult/Mult_out[21] ;
   wire \UUT/Mpath/the_mult/Mult_out[22] ;
   wire \UUT/Mpath/the_mult/Mult_out[23] ;
   wire \UUT/Mpath/the_mult/Mult_out[24] ;
   wire \UUT/Mpath/the_mult/Mult_out[25] ;
   wire \UUT/Mpath/the_mult/Mult_out[26] ;
   wire \UUT/Mpath/the_mult/Mult_out[27] ;
   wire \UUT/Mpath/the_mult/Mult_out[28] ;
   wire \UUT/Mpath/the_mult/Mult_out[29] ;
   wire \UUT/Mpath/the_mult/Mult_out[30] ;
   wire \UUT/Mpath/the_mult/Mult_out[31] ;
   wire \UUT/Mpath/the_mult/Mult_out[32] ;
   wire \UUT/Mpath/the_mult/Mult_out[33] ;
   wire \UUT/Mpath/the_mult/Mult_out[34] ;
   wire \UUT/Mpath/the_mult/Mult_out[35] ;
   wire \UUT/Mpath/the_mult/Mult_out[36] ;
   wire \UUT/Mpath/the_mult/Mult_out[37] ;
   wire \UUT/Mpath/the_mult/Mult_out[38] ;
   wire \UUT/Mpath/the_mult/Mult_out[39] ;
   wire \UUT/Mpath/the_mult/Mult_out[40] ;
   wire \UUT/Mpath/the_mult/Mult_out[41] ;
   wire \UUT/Mpath/the_mult/Mult_out[42] ;
   wire \UUT/Mpath/the_mult/Mult_out[43] ;
   wire \UUT/Mpath/the_mult/Mult_out[44] ;
   wire \UUT/Mpath/the_mult/Mult_out[45] ;
   wire \UUT/Mpath/the_mult/Mult_out[46] ;
   wire \UUT/Mpath/the_mult/Mult_out[47] ;
   wire \UUT/Mpath/the_mult/Mult_out[48] ;
   wire \UUT/Mpath/the_mult/Mult_out[49] ;
   wire \UUT/Mpath/the_mult/Mult_out[50] ;
   wire \UUT/Mpath/the_mult/Mult_out[51] ;
   wire \UUT/Mpath/the_mult/Mult_out[52] ;
   wire \UUT/Mpath/the_mult/Mult_out[53] ;
   wire \UUT/Mpath/the_mult/Mult_out[54] ;
   wire \UUT/Mpath/the_mult/Mult_out[55] ;
   wire \UUT/Mpath/the_mult/Mult_out[56] ;
   wire \UUT/Mpath/the_mult/Mult_out[57] ;
   wire \UUT/Mpath/the_mult/Mult_out[58] ;
   wire \UUT/Mpath/the_mult/Mult_out[59] ;
   wire \UUT/Mpath/the_mult/Mult_out[60] ;
   wire \UUT/Mpath/the_mult/Mult_out[61] ;
   wire \UUT/Mpath/the_mult/Mult_out[62] ;
   wire \UUT/Mpath/the_mult/Mult_out[63] ;
   wire \UUT/Mpath/the_mult/m_mul_command[0] ;
   wire \UUT/Mpath/the_mult/m_mul_command[1] ;
   wire \UUT/Mpath/the_mult/m_mul_command[2] ;
   wire \UUT/Mpath/the_mult/m_mul_command[3] ;
   wire \UUT/Mpath/the_mult/m_mul_command[4] ;
   wire \UUT/Mpath/the_mult/m_mul_command[5] ;
   wire \UUT/Mpath/the_mult/x_mult_out[0] ;
   wire \UUT/Mpath/the_mult/x_mult_out[1] ;
   wire \UUT/Mpath/the_mult/x_mult_out[2] ;
   wire \UUT/Mpath/the_mult/x_mult_out[3] ;
   wire \UUT/Mpath/the_mult/x_mult_out[4] ;
   wire \UUT/Mpath/the_mult/x_mult_out[5] ;
   wire \UUT/Mpath/the_mult/x_mult_out[6] ;
   wire \UUT/Mpath/the_mult/x_mult_out[7] ;
   wire \UUT/Mpath/the_mult/x_mult_out[8] ;
   wire \UUT/Mpath/the_mult/x_mult_out[9] ;
   wire \UUT/Mpath/the_mult/x_mult_out[10] ;
   wire \UUT/Mpath/the_mult/x_mult_out[11] ;
   wire \UUT/Mpath/the_mult/x_mult_out[12] ;
   wire \UUT/Mpath/the_mult/x_mult_out[13] ;
   wire \UUT/Mpath/the_mult/x_mult_out[14] ;
   wire \UUT/Mpath/the_mult/x_mult_out[15] ;
   wire \UUT/Mpath/the_mult/x_mult_out[16] ;
   wire \UUT/Mpath/the_mult/x_mult_out[17] ;
   wire \UUT/Mpath/the_mult/x_mult_out[18] ;
   wire \UUT/Mpath/the_mult/x_mult_out[19] ;
   wire \UUT/Mpath/the_mult/x_mult_out[20] ;
   wire \UUT/Mpath/the_mult/x_mult_out[21] ;
   wire \UUT/Mpath/the_mult/x_mult_out[22] ;
   wire \UUT/Mpath/the_mult/x_mult_out[23] ;
   wire \UUT/Mpath/the_mult/x_mult_out[24] ;
   wire \UUT/Mpath/the_mult/x_mult_out[25] ;
   wire \UUT/Mpath/the_mult/x_mult_out[26] ;
   wire \UUT/Mpath/the_mult/x_mult_out[27] ;
   wire \UUT/Mpath/the_mult/x_mult_out[28] ;
   wire \UUT/Mpath/the_mult/x_mult_out[29] ;
   wire \UUT/Mpath/the_mult/x_mult_out[30] ;
   wire \UUT/Mpath/the_mult/x_mult_out[31] ;
   wire \UUT/Mpath/the_mult/x_mult_out[32] ;
   wire \UUT/Mpath/the_mult/x_mult_out[33] ;
   wire \UUT/Mpath/the_mult/x_mult_out[34] ;
   wire \UUT/Mpath/the_mult/x_mult_out[35] ;
   wire \UUT/Mpath/the_mult/x_mult_out[36] ;
   wire \UUT/Mpath/the_mult/x_mult_out[37] ;
   wire \UUT/Mpath/the_mult/x_mult_out[38] ;
   wire \UUT/Mpath/the_mult/x_mult_out[39] ;
   wire \UUT/Mpath/the_mult/x_mult_out[40] ;
   wire \UUT/Mpath/the_mult/x_mult_out[41] ;
   wire \UUT/Mpath/the_mult/x_mult_out[42] ;
   wire \UUT/Mpath/the_mult/x_mult_out[43] ;
   wire \UUT/Mpath/the_mult/x_mult_out[44] ;
   wire \UUT/Mpath/the_mult/x_mult_out[45] ;
   wire \UUT/Mpath/the_mult/x_mult_out[46] ;
   wire \UUT/Mpath/the_mult/x_mult_out[47] ;
   wire \UUT/Mpath/the_mult/x_mult_out[48] ;
   wire \UUT/Mpath/the_mult/x_mult_out[49] ;
   wire \UUT/Mpath/the_mult/x_mult_out[50] ;
   wire \UUT/Mpath/the_mult/x_mult_out[51] ;
   wire \UUT/Mpath/the_mult/x_mult_out[52] ;
   wire \UUT/Mpath/the_mult/x_mult_out[53] ;
   wire \UUT/Mpath/the_mult/x_mult_out[54] ;
   wire \UUT/Mpath/the_mult/x_mult_out[55] ;
   wire \UUT/Mpath/the_mult/x_mult_out[56] ;
   wire \UUT/Mpath/the_mult/x_mult_out[57] ;
   wire \UUT/Mpath/the_mult/x_mult_out[58] ;
   wire \UUT/Mpath/the_mult/x_mult_out[59] ;
   wire \UUT/Mpath/the_mult/x_mult_out[60] ;
   wire \UUT/Mpath/the_mult/x_mult_out[61] ;
   wire \UUT/Mpath/the_mult/x_mult_out[62] ;
   wire \UUT/Mpath/the_mult/x_mult_out[63] ;
   wire \UUT/Mpath/the_mult/x_mul_command[0] ;
   wire \UUT/Mpath/the_mult/x_mul_command[1] ;
   wire \UUT/Mpath/the_mult/x_mul_command[2] ;
   wire \UUT/Mpath/the_mult/x_mul_command[3] ;
   wire \UUT/Mpath/the_mult/x_mul_command[4] ;
   wire \UUT/Mpath/the_mult/x_mul_command[5] ;
   wire \UUT/Mpath/the_mult/x_operand1[0] ;
   wire \UUT/Mpath/the_mult/x_operand1[1] ;
   wire \UUT/Mpath/the_mult/x_operand1[2] ;
   wire \UUT/Mpath/the_mult/x_operand1[3] ;
   wire \UUT/Mpath/the_mult/x_operand1[4] ;
   wire \UUT/Mpath/the_mult/x_operand1[5] ;
   wire \UUT/Mpath/the_mult/x_operand1[6] ;
   wire \UUT/Mpath/the_mult/x_operand1[7] ;
   wire \UUT/Mpath/the_mult/x_operand1[8] ;
   wire \UUT/Mpath/the_mult/x_operand1[9] ;
   wire \UUT/Mpath/the_mult/x_operand1[10] ;
   wire \UUT/Mpath/the_mult/x_operand1[11] ;
   wire \UUT/Mpath/the_mult/x_operand1[12] ;
   wire \UUT/Mpath/the_mult/x_operand1[13] ;
   wire \UUT/Mpath/the_mult/x_operand1[14] ;
   wire \UUT/Mpath/the_mult/x_operand1[15] ;
   wire \UUT/Mpath/the_mult/x_operand1[16] ;
   wire \UUT/Mpath/the_mult/x_operand1[17] ;
   wire \UUT/Mpath/the_mult/x_operand1[18] ;
   wire \UUT/Mpath/the_mult/x_operand1[19] ;
   wire \UUT/Mpath/the_mult/x_operand1[20] ;
   wire \UUT/Mpath/the_mult/x_operand1[21] ;
   wire \UUT/Mpath/the_mult/x_operand1[22] ;
   wire \UUT/Mpath/the_mult/x_operand1[23] ;
   wire \UUT/Mpath/the_mult/x_operand1[24] ;
   wire \UUT/Mpath/the_mult/x_operand1[25] ;
   wire \UUT/Mpath/the_mult/x_operand1[26] ;
   wire \UUT/Mpath/the_mult/x_operand1[27] ;
   wire \UUT/Mpath/the_mult/x_operand1[28] ;
   wire \UUT/Mpath/the_mult/x_operand1[29] ;
   wire \UUT/Mpath/the_mult/x_operand1[30] ;
   wire \UUT/Mpath/the_mult/x_operand1[31] ;
   wire \UUT/Mpath/the_memhandle/N242 ;
   wire \UUT/Mpath/the_memhandle/N241 ;
   wire \UUT/Mpath/the_memhandle/N240 ;
   wire \UUT/Mpath/the_memhandle/N239 ;
   wire \UUT/Mpath/the_memhandle/N238 ;
   wire \UUT/Mpath/the_memhandle/N237 ;
   wire \UUT/Mpath/the_memhandle/N236 ;
   wire \UUT/Mpath/the_memhandle/N235 ;
   wire \UUT/Mpath/the_memhandle/N234 ;
   wire \UUT/Mpath/the_memhandle/N120 ;
   wire \UUT/Mpath/the_memhandle/N86 ;
   wire \UUT/Mpath/the_memhandle/N76 ;
   wire \UUT/Mpath/the_memhandle/N72 ;
   wire \UUT/Mpath/the_memhandle/N39 ;
   wire \UUT/Mpath/the_memhandle/N37 ;
   wire \UUT/Mpath/the_memhandle/N36 ;
   wire \UUT/Mpath/the_memhandle/N34 ;
   wire \UUT/Mpath/the_memhandle/smdr_out[8] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[9] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[10] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[11] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[12] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[13] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[14] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[15] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[16] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[17] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[18] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[19] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[20] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[21] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[22] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[23] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[24] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[25] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[26] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[27] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[28] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[29] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[30] ;
   wire \UUT/Mpath/the_memhandle/smdr_out[31] ;
   wire \localbus/N338 ;
   wire \localbus/N335 ;
   wire \localbus/N329 ;
   wire \localbus/N322 ;
   wire \localbus/N321 ;
   wire \localbus/N320 ;
   wire \localbus/N319 ;
   wire \localbus/N318 ;
   wire \localbus/N293 ;
   wire \localbus/N258 ;
   wire \localbus/N257 ;
   wire \localbus/N256 ;
   wire \localbus/N252 ;
   wire \localbus/N251 ;
   wire \localbus/N250 ;
   wire \localbus/N229 ;
   wire \localbus/N227 ;
   wire \localbus/N225 ;
   wire \localbus/N219 ;
   wire \localbus/N218 ;
   wire \localbus/N214 ;
   wire \localbus/N95 ;
   wire \localbus/N93 ;
   wire \localbus/c2_op[OP][1] ;
   wire \localbus/c2_op[SLAVE][0] ;
   wire \localbus/c2_op[SLAVE][1] ;
   wire \localbus/c2_op[SLAVE][2] ;
   wire \localbus/c2_op[MASTER] ;
   wire \localbus/N90 ;
   wire \localbus/N89 ;
   wire \localbus/N86 ;
   wire \localbus/N85 ;
   wire \localbus/N62 ;
   wire \localbus/N61 ;
   wire \localbus/N60 ;
   wire \localbus/N57 ;
   wire \localbus/N56 ;
   wire \localbus/N55 ;
   wire \localbus/N51 ;
   wire \localbus/c1_addr_outbus[13] ;
   wire \localbus/c1_addr_outbus[14] ;
   wire \localbus/c1_addr_outbus[15] ;
   wire \localbus/c1_addr_outbus[16] ;
   wire \localbus/c1_addr_outbus[17] ;
   wire \localbus/c1_addr_outbus[18] ;
   wire \localbus/c1_addr_outbus[19] ;
   wire \localbus/c1_addr_outbus[20] ;
   wire \localbus/c1_addr_outbus[21] ;
   wire \localbus/c1_addr_outbus[22] ;
   wire \localbus/c1_addr_outbus[23] ;
   wire \localbus/c1_addr_outbus[24] ;
   wire \localbus/c1_addr_outbus[25] ;
   wire \localbus/c1_addr_outbus[26] ;
   wire \localbus/c1_addr_outbus[27] ;
   wire \localbus/c1_addr_outbus[28] ;
   wire \localbus/c1_addr_outbus[29] ;
   wire \localbus/c1_addr_outbus[30] ;
   wire \localbus/N50 ;
   wire \localbus/N46 ;
   wire \localbus/c1_op[OP][0] ;
   wire \localbus/c1_op[OP][1] ;
   wire \localbus/c1_op[SLAVE][0] ;
   wire \localbus/c1_op[MASTER] ;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1011;
   wire n1012;
   wire n1014;
   wire n1015;
   wire n1017;
   wire n1018;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1178;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2594;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2639;
   wire n2642;
   wire n2645;
   wire n2648;
   wire n2651;
   wire n2654;
   wire n2657;
   wire n2660;
   wire n2663;
   wire n2666;
   wire n2668;
   wire n2671;
   wire n2677;
   wire n2679;
   wire n2682;
   wire n2685;
   wire n2688;
   wire n2691;
   wire n2694;
   wire n2698;
   wire n2725;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2732;
   wire n2735;
   wire n2737;
   wire n2739;
   wire n2741;
   wire n2748;
   wire n2750;
   wire n2752;
   wire n2754;
   wire n2756;
   wire n2781;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3711;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3773;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3804;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire n3844;
   wire n3845;
   wire n3846;
   wire n3847;
   wire n3848;
   wire n3849;
   wire n3850;
   wire n3851;
   wire n3852;
   wire n3853;
   wire n3854;
   wire n3855;
   wire n3856;
   wire n3857;
   wire n3858;
   wire n3859;
   wire n3860;
   wire n3861;
   wire n3862;
   wire n3863;
   wire n3864;
   wire n3865;
   wire n3866;
   wire n3867;
   wire n3868;
   wire n3869;
   wire n3870;
   wire n3871;
   wire n3872;
   wire n3873;
   wire n3874;
   wire n3875;
   wire n3876;
   wire n3877;
   wire n3878;
   wire n3879;
   wire n3880;
   wire n3881;
   wire n3882;
   wire n3883;
   wire n3884;
   wire n3885;
   wire n3886;
   wire n3887;
   wire n3888;
   wire n3889;
   wire n3890;
   wire n3891;
   wire n3892;
   wire n3893;
   wire n3894;
   wire n3895;
   wire n3896;
   wire n3897;
   wire n3898;
   wire n3899;
   wire n3900;
   wire n3901;
   wire n3902;
   wire n3903;
   wire n3904;
   wire n3905;
   wire n3906;
   wire n3907;
   wire n3908;
   wire n3909;
   wire n3910;
   wire n3911;
   wire n3912;
   wire n3913;
   wire n3914;
   wire n3915;
   wire n3916;
   wire n3917;
   wire n3918;
   wire n3919;
   wire n3920;
   wire n3921;
   wire n3922;
   wire n3923;
   wire n3924;
   wire n3925;
   wire n3926;
   wire n3927;
   wire n3928;
   wire n3929;
   wire n3930;
   wire n3931;
   wire n3932;
   wire n3933;
   wire n3934;
   wire n3935;
   wire n3936;
   wire n3937;
   wire n3938;
   wire n3939;
   wire n3940;
   wire n3941;
   wire n3942;
   wire n3943;
   wire n3944;
   wire n3945;
   wire n3946;
   wire n3947;
   wire n3948;
   wire n3949;
   wire n3950;
   wire n3951;
   wire n3952;
   wire n3953;
   wire n3954;
   wire n3955;
   wire n3956;
   wire n3957;
   wire n3958;
   wire n3959;
   wire n3960;
   wire n3961;
   wire n3962;
   wire n3963;
   wire n3964;
   wire n3965;
   wire n3966;
   wire n3967;
   wire n3968;
   wire n3969;
   wire n3970;
   wire n3971;
   wire n3972;
   wire n3973;
   wire n3974;
   wire n3975;
   wire n3976;
   wire n3977;
   wire n3978;
   wire n3979;
   wire n3980;
   wire n3981;
   wire n3982;
   wire n3983;
   wire n3984;
   wire n3985;
   wire n3986;
   wire n3987;
   wire n3988;
   wire n3989;
   wire n3990;
   wire n3991;
   wire n3992;
   wire n3993;
   wire n3994;
   wire n3995;
   wire n3996;
   wire n3997;
   wire n3998;
   wire n3999;
   wire n4000;
   wire n4001;
   wire n4002;
   wire n4003;
   wire n4004;
   wire n4005;
   wire n4006;
   wire n4007;
   wire n4008;
   wire n4009;
   wire n4010;
   wire n4011;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4016;
   wire n4017;
   wire n4018;
   wire n4019;
   wire n4020;
   wire n4021;
   wire n4022;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4026;
   wire n4027;
   wire n4028;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire n4042;
   wire n4043;
   wire n4044;
   wire n4045;
   wire n4046;
   wire n4047;
   wire n4048;
   wire n4049;
   wire n4050;
   wire n4051;
   wire n4052;
   wire n4053;
   wire n4054;
   wire n4055;
   wire n4056;
   wire n4057;
   wire n4058;
   wire n4059;
   wire n4060;
   wire n4063;
   wire n4064;
   wire n4065;
   wire n4066;
   wire n4067;
   wire n4068;
   wire n4069;
   wire n4070;
   wire n4071;
   wire n4072;
   wire n4073;
   wire n4074;
   wire n4075;
   wire n4076;
   wire n4077;
   wire n4078;
   wire n4079;
   wire n4080;
   wire n4081;
   wire n4082;
   wire n4083;
   wire n4084;
   wire n4085;
   wire n4086;
   wire n4087;
   wire n4088;
   wire n4089;
   wire n4090;
   wire n4091;
   wire n4092;
   wire n4093;
   wire n4094;
   wire n4095;
   wire n4096;
   wire n4097;
   wire n4098;
   wire n4099;
   wire n4100;
   wire n4101;
   wire n4102;
   wire n4103;
   wire n4104;
   wire n4105;
   wire n4106;
   wire n4107;
   wire n4108;
   wire n4109;
   wire n4110;
   wire n4111;
   wire n4112;
   wire n4113;
   wire n4114;
   wire n4115;
   wire n4116;
   wire n4117;
   wire n4118;
   wire n4119;
   wire n4120;
   wire n4121;
   wire n4122;
   wire n4123;
   wire n4124;
   wire n4125;
   wire n4126;
   wire n4127;
   wire n4128;
   wire n4129;
   wire n4130;
   wire n4131;
   wire n4132;
   wire n4133;
   wire n4134;
   wire n4135;
   wire n4136;
   wire n4137;
   wire n4138;
   wire n4139;
   wire n4140;
   wire n4141;
   wire n4142;
   wire n4143;
   wire n4144;
   wire n4145;
   wire n4146;
   wire n4147;
   wire n4148;
   wire n4149;
   wire n4150;
   wire n4151;
   wire n4152;
   wire n4153;
   wire n4154;
   wire n4155;
   wire n4156;
   wire n4157;
   wire n4158;
   wire n4159;
   wire n4160;
   wire n4161;
   wire n4162;
   wire n4163;
   wire n4164;
   wire n4165;
   wire n4166;
   wire n4167;
   wire n4168;
   wire n4169;
   wire n4170;
   wire n4171;
   wire n4172;
   wire n4173;
   wire n4174;
   wire n4175;
   wire n4176;
   wire n4177;
   wire n4178;
   wire n4179;
   wire n4180;
   wire n4181;
   wire n4182;
   wire n4183;
   wire n4184;
   wire n4185;
   wire n4186;
   wire n4187;
   wire n4188;
   wire n4189;
   wire n4190;
   wire n4191;
   wire n4192;
   wire n4193;
   wire n4194;
   wire n4195;
   wire n4196;
   wire n4197;
   wire n4198;
   wire n4199;
   wire n4200;
   wire n4201;
   wire n4202;
   wire n4203;
   wire n4204;
   wire n4205;
   wire n4206;
   wire n4207;
   wire n4208;
   wire n4209;
   wire n4210;
   wire n4211;
   wire n4212;
   wire n4213;
   wire n4214;
   wire n4215;
   wire n4216;
   wire n4217;
   wire n4218;
   wire n4219;
   wire n4220;
   wire n4221;
   wire n4222;
   wire n4223;
   wire n4224;
   wire n4225;
   wire n4226;
   wire n4227;
   wire n4228;
   wire n4229;
   wire n4230;
   wire n4231;
   wire n4232;
   wire n4233;
   wire n4234;
   wire n4235;
   wire n4236;
   wire n4237;
   wire n4238;
   wire n4239;
   wire n4240;
   wire n4241;
   wire n4242;
   wire n4243;
   wire n4244;
   wire n4245;
   wire n4246;
   wire n4247;
   wire n4248;
   wire n4249;
   wire n4250;
   wire n4251;
   wire n4252;
   wire n4253;
   wire n4254;
   wire n4255;
   wire n4256;
   wire n4257;
   wire n4258;
   wire n4259;
   wire n4260;
   wire n4261;
   wire n4262;
   wire n4263;
   wire n4264;
   wire n4265;
   wire n4266;
   wire n4267;
   wire n4268;
   wire n4269;
   wire n4270;
   wire n4271;
   wire n4272;
   wire n4273;
   wire n4274;
   wire n4275;
   wire n4276;
   wire n4277;
   wire n4278;
   wire n4279;
   wire n4280;
   wire n4281;
   wire n4282;
   wire n4283;
   wire n4284;
   wire n4285;
   wire n4286;
   wire n4287;
   wire n4288;
   wire n4289;
   wire n4290;
   wire n4291;
   wire n4292;
   wire n4293;
   wire n4294;
   wire n4295;
   wire n4296;
   wire n4297;
   wire n4298;
   wire n4299;
   wire n4300;
   wire n4301;
   wire n4302;
   wire n4303;
   wire n4304;
   wire n4305;
   wire n4306;
   wire n4307;
   wire n4308;
   wire n4309;
   wire n4310;
   wire n4311;
   wire n4312;
   wire n4313;
   wire n4314;
   wire n4315;
   wire n4316;
   wire n4317;
   wire n4318;
   wire n4319;
   wire n4320;
   wire n4321;
   wire n4322;
   wire n4324;
   wire n4325;
   wire n4327;
   wire n4328;
   wire n4329;
   wire n4330;
   wire n4331;
   wire n4332;
   wire n4333;
   wire n4334;
   wire n4335;
   wire n4337;
   wire n4339;
   wire n4340;
   wire n4343;
   wire n4344;
   wire n4345;
   wire n4346;
   wire n4347;
   wire n4348;
   wire n4349;
   wire n4350;
   wire n4352;
   wire n4353;
   wire n4354;
   wire n4355;
   wire n4356;
   wire n4357;
   wire n4358;
   wire n4359;
   wire n4360;
   wire n4361;
   wire n4362;
   wire n4363;
   wire n4364;
   wire n4365;
   wire n4366;
   wire n4367;
   wire n4368;
   wire n4369;
   wire n4370;
   wire n4371;
   wire n4372;
   wire n4373;
   wire n4374;
   wire n4375;
   wire n4376;
   wire n4377;
   wire n4378;
   wire n4379;
   wire n4380;
   wire n4381;
   wire n4382;
   wire n4383;
   wire n4384;
   wire n4385;
   wire n4386;
   wire n4387;
   wire n4388;
   wire n4389;
   wire n4390;
   wire n4391;
   wire n4392;
   wire n4393;
   wire n4394;
   wire n4395;
   wire n4396;
   wire n4397;
   wire n4398;
   wire n4399;
   wire n4400;
   wire n4401;
   wire n4402;
   wire n4403;
   wire n4404;
   wire n4405;
   wire n4406;
   wire n4407;
   wire n4408;
   wire n4409;
   wire n4411;
   wire n4412;
   wire n4413;
   wire n4414;
   wire n4415;
   wire n4416;
   wire n4417;
   wire n4418;
   wire n4419;
   wire n4420;
   wire n4421;
   wire n4422;
   wire n4423;
   wire n4424;
   wire n4425;
   wire n4426;
   wire n4427;
   wire n4428;
   wire n4429;
   wire n4430;
   wire n4431;
   wire n4432;
   wire n4433;
   wire n4434;
   wire n4435;
   wire n4436;
   wire n4437;
   wire n4438;
   wire n4439;
   wire n4440;
   wire n4441;
   wire n4442;
   wire n4443;
   wire n4444;
   wire n4445;
   wire n4446;
   wire n4447;
   wire n4448;
   wire n4449;
   wire n4450;
   wire n4451;
   wire n4452;
   wire n4453;
   wire n4454;
   wire n4455;
   wire n4456;
   wire n4457;
   wire n4458;
   wire n4459;
   wire n4460;
   wire n4461;
   wire n4462;
   wire n4463;
   wire n4464;
   wire n4465;
   wire n4466;
   wire n4467;
   wire n4468;
   wire n4469;
   wire n4470;
   wire n4471;
   wire n4472;
   wire n4473;
   wire n4474;
   wire n4475;
   wire n4476;
   wire n4477;
   wire n4478;
   wire n4479;
   wire n4480;
   wire n4481;
   wire n4482;
   wire n4483;
   wire n4484;
   wire n4485;
   wire n4486;
   wire n4487;
   wire n4488;
   wire n4489;
   wire n4490;
   wire n4491;
   wire n4492;
   wire n4493;
   wire n4494;
   wire n4495;
   wire n4496;
   wire n4497;
   wire n4498;
   wire n4499;
   wire n4500;
   wire n4501;
   wire n4502;
   wire n4503;
   wire n4504;
   wire n4505;
   wire n4506;
   wire n4507;
   wire n4508;
   wire n4509;
   wire n4510;
   wire n4511;
   wire n4512;
   wire n4513;
   wire n4514;
   wire n4515;
   wire n4516;
   wire n4517;
   wire n4518;
   wire n4519;
   wire n4520;
   wire n4521;
   wire n4522;
   wire n4523;
   wire n4524;
   wire n4525;
   wire n4526;
   wire n4527;
   wire n4528;
   wire n4529;
   wire n4530;
   wire n4531;
   wire n4532;
   wire n4533;
   wire n4534;
   wire n4535;
   wire n4536;
   wire n4537;
   wire n4538;
   wire n4539;
   wire n4540;
   wire n4541;
   wire n4542;
   wire n4543;
   wire n4544;
   wire n4545;
   wire n4546;
   wire n4547;
   wire n4548;
   wire n4549;
   wire n4550;
   wire n4551;
   wire n4552;
   wire n4553;
   wire n4554;
   wire n4555;
   wire n4556;
   wire n4557;
   wire n4558;
   wire n4559;
   wire n4560;
   wire n4561;
   wire n4562;
   wire n4563;
   wire n4564;
   wire n4565;
   wire n4566;
   wire n4567;
   wire n4568;
   wire n4569;
   wire n4570;
   wire n4571;
   wire n4572;
   wire n4573;
   wire n4574;
   wire n4575;
   wire n4576;
   wire n4577;
   wire n4578;
   wire n4579;
   wire n4580;
   wire n4581;
   wire n4582;
   wire n4583;
   wire n4584;
   wire n4585;
   wire n4586;
   wire n4587;
   wire n4588;
   wire n4589;
   wire n4590;
   wire n4591;
   wire n4592;
   wire n4593;
   wire n4594;
   wire n4595;
   wire n4596;
   wire n4597;
   wire n4598;
   wire n4599;
   wire n4600;
   wire n4601;
   wire n4602;
   wire n4603;
   wire n4604;
   wire n4605;
   wire n4606;
   wire n4607;
   wire n4608;
   wire n4609;
   wire n4610;
   wire n4611;
   wire n4612;
   wire n4613;
   wire n4614;
   wire n4615;
   wire n4616;
   wire n4617;
   wire n4618;
   wire n4619;
   wire n4620;
   wire n4621;
   wire n4622;
   wire n4623;
   wire n4624;
   wire n4625;
   wire n4626;
   wire n4627;
   wire n4628;
   wire n4629;
   wire n4630;
   wire n4631;
   wire n4632;
   wire n4633;
   wire n4634;
   wire n4635;
   wire n4636;
   wire n4637;
   wire n4638;
   wire n4639;
   wire n4640;
   wire n4641;
   wire n4642;
   wire n4643;
   wire n4644;
   wire n4645;
   wire n4646;
   wire n4647;
   wire n4648;
   wire n4649;
   wire n4650;
   wire n4651;
   wire n4652;
   wire n4653;
   wire n4654;
   wire n4655;
   wire n4656;
   wire n4657;
   wire n4658;
   wire n4659;
   wire n4660;
   wire n4661;
   wire n4662;
   wire n4663;
   wire n4664;
   wire n4665;
   wire n4666;
   wire n4667;
   wire n4668;
   wire n4669;
   wire n4670;
   wire n4671;
   wire n4672;
   wire n4673;
   wire n4674;
   wire n4675;
   wire n4676;
   wire n4677;
   wire n4678;
   wire n4679;
   wire n4680;
   wire n4681;
   wire n4682;
   wire n4683;
   wire n4684;
   wire n4685;
   wire n4686;
   wire n4687;
   wire n4688;
   wire n4689;
   wire n4690;
   wire n4691;
   wire n4692;
   wire n4693;
   wire n4694;
   wire n4695;
   wire n4696;
   wire n4697;
   wire n4698;
   wire n4699;
   wire n4700;
   wire n4701;
   wire n4702;
   wire n4703;
   wire n4704;
   wire n4705;
   wire n4706;
   wire n4707;
   wire n4708;
   wire n4709;
   wire n4710;
   wire n4711;
   wire n4712;
   wire n4713;
   wire n4714;
   wire n4715;
   wire n4716;
   wire n4717;
   wire n4718;
   wire n4719;
   wire n4720;
   wire n4721;
   wire n4722;
   wire n4723;
   wire n4724;
   wire n4725;
   wire n4726;
   wire n4727;
   wire n4728;
   wire n4729;
   wire n4730;
   wire n4731;
   wire n4732;
   wire n4733;
   wire n4734;
   wire n4735;
   wire n4736;
   wire n4737;
   wire n4738;
   wire n4739;
   wire n4740;
   wire n4741;
   wire n4742;
   wire n4743;
   wire n4744;
   wire n4745;
   wire n4746;
   wire n4747;
   wire n4748;
   wire n4749;
   wire n4750;
   wire n4751;
   wire n4752;
   wire n4753;
   wire n4754;
   wire n4755;
   wire n4756;
   wire n4757;
   wire n4758;
   wire n4759;
   wire n4760;
   wire n4761;
   wire n4762;
   wire n4763;
   wire n4764;
   wire n4765;
   wire n4766;
   wire n4767;
   wire n4768;
   wire n4769;
   wire n4770;
   wire n4771;
   wire n4772;
   wire n4773;
   wire n4774;
   wire n4775;
   wire n4776;
   wire n4777;
   wire n4778;
   wire n4779;
   wire n4780;
   wire n4781;
   wire n4782;
   wire n4783;
   wire n4784;
   wire n4785;
   wire n4786;
   wire n4787;
   wire n4788;
   wire n4789;
   wire n4790;
   wire n4791;
   wire n4792;
   wire n4793;
   wire n4794;
   wire n4795;
   wire n4796;
   wire n4797;
   wire n4798;
   wire n4799;
   wire n4800;
   wire n4801;
   wire n4802;
   wire n4803;
   wire n4804;
   wire n4805;
   wire n4806;
   wire n4807;
   wire n4808;
   wire n4809;
   wire n4810;
   wire n4811;
   wire n4812;
   wire n4813;
   wire n4814;
   wire n4815;
   wire n4816;
   wire n4817;
   wire n4818;
   wire n4819;
   wire n4820;
   wire n4821;
   wire n4822;
   wire n4823;
   wire n4824;
   wire n4825;
   wire n4826;
   wire n4827;
   wire n4828;
   wire n4829;
   wire n4830;
   wire n4831;
   wire n4832;
   wire n4833;
   wire n4834;
   wire n4835;
   wire n4836;
   wire n4837;
   wire n4838;
   wire n4839;
   wire n4840;
   wire n4841;
   wire n4842;
   wire n4843;
   wire n4844;
   wire n4845;
   wire n4846;
   wire n4847;
   wire n4848;
   wire n4849;
   wire n4850;
   wire n4851;
   wire n4852;
   wire n4853;
   wire n4854;
   wire n4855;
   wire n4856;
   wire n4857;
   wire n4858;
   wire n4859;
   wire n4860;
   wire n4861;
   wire n4862;
   wire n4863;
   wire n4864;
   wire n4865;
   wire n4866;
   wire n4867;
   wire n4868;
   wire n4869;
   wire n4870;
   wire n4871;
   wire n4872;
   wire n4873;
   wire n4874;
   wire n4875;
   wire n4876;
   wire n4877;
   wire n4878;
   wire n4879;
   wire n4880;
   wire n4881;
   wire n4882;
   wire n4883;
   wire n4884;
   wire n4885;
   wire n4886;
   wire n4887;
   wire n4888;
   wire n4889;
   wire n4890;
   wire n4891;
   wire n4892;
   wire n4893;
   wire n4894;
   wire n4895;
   wire n4896;
   wire n4897;
   wire n4898;
   wire n4899;
   wire n4900;
   wire n4901;
   wire n4902;
   wire n4903;
   wire n4904;
   wire n4905;
   wire n4906;
   wire n4907;
   wire n4908;
   wire n4909;
   wire n4910;
   wire n4911;
   wire n4912;
   wire n4913;
   wire n4914;
   wire n4915;
   wire n4916;
   wire n4917;
   wire n4918;
   wire n4919;
   wire n4920;
   wire n4921;
   wire n4922;
   wire n4923;
   wire n4924;
   wire n4925;
   wire n4926;
   wire n4927;
   wire n4928;
   wire n4929;
   wire n4930;
   wire n4931;
   wire n4932;
   wire n4933;
   wire n4934;
   wire n4935;
   wire n4936;
   wire n4937;
   wire n4938;
   wire n4939;
   wire n4940;
   wire n4941;
   wire n4942;
   wire n4943;
   wire n4944;
   wire n4945;
   wire n4946;
   wire n4947;
   wire n4948;
   wire n4949;
   wire n4950;
   wire n4951;
   wire n4952;
   wire n4953;
   wire n4954;
   wire n4955;
   wire n4956;
   wire n4957;
   wire n4958;
   wire n4959;
   wire n4960;
   wire n4961;
   wire n4962;
   wire n4963;
   wire n4964;
   wire n4965;
   wire n4966;
   wire n4967;
   wire n4968;
   wire n4969;
   wire n4970;
   wire n4971;
   wire n4972;
   wire n4973;
   wire n4974;
   wire n4975;
   wire n4976;
   wire n4977;
   wire n4978;
   wire n4979;
   wire n4980;
   wire n4981;
   wire n4982;
   wire n4983;
   wire n4984;
   wire n4985;
   wire n4986;
   wire n4987;
   wire n4988;
   wire n4989;
   wire n4990;
   wire n4991;
   wire n4992;
   wire n4993;
   wire n4994;
   wire n4995;
   wire n4996;
   wire n4997;
   wire n4998;
   wire n4999;
   wire n5000;
   wire n5001;
   wire n5002;
   wire n5003;
   wire n5004;
   wire n5005;
   wire n5006;
   wire n5007;
   wire n5008;
   wire n5009;
   wire n5010;
   wire n5011;
   wire n5012;
   wire n5013;
   wire n5014;
   wire n5015;
   wire n5016;
   wire n5017;
   wire n5018;
   wire n5019;
   wire n5020;
   wire n5021;
   wire n5022;
   wire n5023;
   wire n5024;
   wire n5025;
   wire n5026;
   wire n5027;
   wire n5028;
   wire n5029;
   wire n5030;
   wire n5031;
   wire n5032;
   wire n5033;
   wire n5034;
   wire n5035;
   wire n5036;
   wire n5037;
   wire n5038;
   wire n5039;
   wire n5040;
   wire n5041;
   wire n5042;
   wire n5043;
   wire n5044;
   wire n5045;
   wire n5046;
   wire n5047;
   wire n5048;
   wire n5049;
   wire n5050;
   wire n5051;
   wire n5052;
   wire n5053;
   wire n5054;
   wire n5055;
   wire n5056;
   wire n5057;
   wire n5058;
   wire n5059;
   wire n5060;
   wire n5061;
   wire n5062;
   wire n5063;
   wire n5064;
   wire n5065;
   wire n5066;
   wire n5067;
   wire n5068;
   wire n5069;
   wire n5070;
   wire n5071;
   wire n5072;
   wire n5073;
   wire n5074;
   wire n5075;
   wire n5076;
   wire n5077;
   wire n5078;
   wire n5079;
   wire n5080;
   wire n5081;
   wire n5082;
   wire n5083;
   wire n5084;
   wire n5085;
   wire n5086;
   wire n5087;
   wire n5088;
   wire n5089;
   wire n5090;
   wire n5091;
   wire n5092;
   wire n5093;
   wire n5094;
   wire n5095;
   wire n5096;
   wire n5097;
   wire n5098;
   wire n5099;
   wire n5100;
   wire n5101;
   wire n5102;
   wire n5103;
   wire n5104;
   wire n5105;
   wire n5106;
   wire n5107;
   wire n5108;
   wire n5109;
   wire n5110;
   wire n5111;
   wire n5112;
   wire n5113;
   wire n5114;
   wire n5115;
   wire n5116;
   wire n5117;
   wire n5118;
   wire n5119;
   wire n5120;
   wire n5121;
   wire n5122;
   wire n5123;
   wire n5124;
   wire n5125;
   wire n5126;
   wire n5127;
   wire n5128;
   wire n5129;
   wire n5130;
   wire n5131;
   wire n5132;
   wire n5133;
   wire n5134;
   wire n5135;
   wire n5136;
   wire n5137;
   wire n5138;
   wire n5139;
   wire n5140;
   wire n5141;
   wire n5142;
   wire n5143;
   wire n5144;
   wire n5145;
   wire n5146;
   wire n5147;
   wire n5148;
   wire n5149;
   wire n5150;
   wire n5151;
   wire n5152;
   wire n5153;
   wire n5154;
   wire n5155;
   wire n5156;
   wire n5157;
   wire n5158;
   wire n5159;
   wire n5160;
   wire n5161;
   wire n5162;
   wire n5163;
   wire n5164;
   wire n5165;
   wire n5166;
   wire n5167;
   wire n5168;
   wire n5169;
   wire n5170;
   wire n5171;
   wire n5172;
   wire n5173;
   wire n5174;
   wire n5175;
   wire n5176;
   wire n5177;
   wire n5178;
   wire n5179;
   wire n5180;
   wire n5181;
   wire n5182;
   wire n5183;
   wire n5184;
   wire n5185;
   wire n5186;
   wire n5187;
   wire n5188;
   wire n5189;
   wire n5190;
   wire n5191;
   wire n5192;
   wire n5193;
   wire n5194;
   wire n5195;
   wire n5196;
   wire n5197;
   wire n5198;
   wire n5199;
   wire n5200;
   wire n5201;
   wire n5202;
   wire n5203;
   wire n5204;
   wire n5205;
   wire n5206;
   wire n5207;
   wire n5208;
   wire n5209;
   wire n5210;
   wire n5211;
   wire n5212;
   wire n5213;
   wire n5214;
   wire n5215;
   wire n5216;
   wire n5217;
   wire n5218;
   wire n5219;
   wire n5220;
   wire n5221;
   wire n5222;
   wire n5223;
   wire n5224;
   wire n5225;
   wire n5226;
   wire n5227;
   wire n5228;
   wire n5229;
   wire n5230;
   wire n5231;
   wire n5232;
   wire n5233;
   wire n5234;
   wire n5235;
   wire n5236;
   wire n5237;
   wire n5238;
   wire n5239;
   wire n5240;
   wire n5241;
   wire n5242;
   wire n5243;
   wire n5244;
   wire n5245;
   wire n5246;
   wire n5247;
   wire n5248;
   wire n5249;
   wire n5250;
   wire n5251;
   wire n5252;
   wire n5253;
   wire n5254;
   wire n5255;
   wire n5256;
   wire n5257;
   wire n5258;
   wire n5259;
   wire n5260;
   wire n5261;
   wire n5262;
   wire n5263;
   wire n5264;
   wire n5265;
   wire n5266;
   wire n5267;
   wire n5268;
   wire n5269;
   wire n5270;
   wire n5271;
   wire n5272;
   wire n5273;
   wire n5274;
   wire n5275;
   wire n5276;
   wire n5277;
   wire n5278;
   wire n5279;
   wire n5280;
   wire n5281;
   wire n5282;
   wire n5283;
   wire n5284;
   wire n5285;
   wire n5286;
   wire n5287;
   wire n5288;
   wire n5289;
   wire n5290;
   wire n5291;
   wire n5292;
   wire n5293;
   wire n5294;
   wire n5295;
   wire n5296;
   wire n5297;
   wire n5298;
   wire n5299;
   wire n5300;
   wire n5301;
   wire n5302;
   wire n5303;
   wire n5304;
   wire n5305;
   wire n5306;
   wire n5307;
   wire n5308;
   wire n5309;
   wire n5310;
   wire n5311;
   wire n5312;
   wire n5313;
   wire n5314;
   wire n5315;
   wire n5316;
   wire n5317;
   wire n5318;
   wire n5319;
   wire n5320;
   wire n5321;
   wire n5322;
   wire n5323;
   wire n5324;
   wire n5325;
   wire n5326;
   wire n5327;
   wire n5328;
   wire n5329;
   wire n5330;
   wire n5331;
   wire n5332;
   wire n5333;
   wire n5334;
   wire n5335;
   wire n5336;
   wire n5337;
   wire n5338;
   wire n5339;
   wire n5340;
   wire n5341;
   wire n5342;
   wire n5343;
   wire n5344;
   wire n5345;
   wire n5346;
   wire n5347;
   wire n5348;
   wire n5349;
   wire n5350;
   wire n5351;
   wire n5352;
   wire n5353;
   wire n5354;
   wire n5355;
   wire n5356;
   wire n5357;
   wire n5358;
   wire n5359;
   wire n5360;
   wire n5361;
   wire n5362;
   wire n5363;
   wire n5364;
   wire n5365;
   wire n5366;
   wire n5367;
   wire n5368;
   wire n5369;
   wire n5370;
   wire n5371;
   wire n5372;
   wire n5373;
   wire n5374;
   wire n5375;
   wire n5376;
   wire n5377;
   wire n5378;
   wire n5379;
   wire n5380;
   wire n5381;
   wire n5382;
   wire n5383;
   wire n5384;
   wire n5385;
   wire n5386;
   wire n5387;
   wire n5388;
   wire n5389;
   wire n5390;
   wire n5391;
   wire n5392;
   wire n5393;
   wire n5394;
   wire n5395;
   wire n5396;
   wire n5397;
   wire n5398;
   wire n5399;
   wire n5400;
   wire n5401;
   wire n5402;
   wire n5403;
   wire n5404;
   wire n5405;
   wire n5406;
   wire n5407;
   wire n5408;
   wire n5409;
   wire n5410;
   wire n5411;
   wire n5412;
   wire n5413;
   wire n5414;
   wire n5415;
   wire n5416;
   wire n5417;
   wire n5418;
   wire n5419;
   wire n5420;
   wire n5421;
   wire n5422;
   wire n5423;
   wire n5424;
   wire n5425;
   wire n5426;
   wire n5427;
   wire n5428;
   wire n5429;
   wire n5430;
   wire n5431;
   wire n5432;
   wire n5433;
   wire n5434;
   wire n5435;
   wire n5436;
   wire n5437;
   wire n5438;
   wire n5439;
   wire n5440;
   wire n5441;
   wire n5442;
   wire n5443;
   wire n5444;
   wire n5445;
   wire n5446;
   wire n5447;
   wire n5448;
   wire n5449;
   wire n5450;
   wire n5451;
   wire n5452;
   wire n5454;
   wire n5455;
   wire n5456;
   wire n5457;
   wire n5458;
   wire n5459;
   wire n5460;
   wire n5461;
   wire n5462;
   wire n5463;
   wire n5464;
   wire n5465;
   wire n5466;
   wire n5467;
   wire n5468;
   wire n5469;
   wire n5470;
   wire n5471;
   wire n5472;
   wire n5473;
   wire n5474;
   wire n5475;
   wire n5476;
   wire n5477;
   wire n5478;
   wire n5479;
   wire n5480;
   wire n5481;
   wire n5482;
   wire n5483;
   wire n5484;
   wire n5485;
   wire n5486;
   wire n5487;
   wire n5488;
   wire n5489;
   wire n5490;
   wire n5491;
   wire n5492;
   wire n5493;
   wire n5494;
   wire n5495;
   wire n5496;
   wire n5497;
   wire n5498;
   wire n5499;
   wire n5500;
   wire n5501;
   wire n5502;
   wire n5503;
   wire n5504;
   wire n5505;
   wire n5506;
   wire n5507;
   wire n5508;
   wire n5509;
   wire n5510;
   wire n5511;
   wire n5512;
   wire n5513;
   wire n5514;
   wire n5515;
   wire n5516;
   wire n5517;
   wire n5518;
   wire n5519;
   wire n5520;
   wire n5521;
   wire n5522;
   wire n5523;
   wire n5524;
   wire n5525;
   wire n5526;
   wire n5527;
   wire n5528;
   wire n5529;
   wire n5530;
   wire n5531;
   wire n5532;
   wire n5533;
   wire n5534;
   wire n5535;
   wire n5536;
   wire n5537;
   wire n5538;
   wire n5539;
   wire n5540;
   wire n5541;
   wire n5542;
   wire n5543;
   wire n5544;
   wire n5545;
   wire n5546;
   wire n5547;
   wire n5548;
   wire n5549;
   wire n5551;
   wire n5552;
   wire n5553;
   wire n5554;
   wire n5555;
   wire n5557;
   wire n5558;
   wire n5559;
   wire n5560;
   wire n5561;
   wire n5562;
   wire n5563;
   wire n5564;
   wire n5565;
   wire n5566;
   wire n5567;
   wire n5568;
   wire n5569;
   wire n5570;
   wire n5571;
   wire n5572;
   wire n5573;
   wire n5574;
   wire n5575;
   wire n5576;
   wire n5577;
   wire n5578;
   wire n5579;
   wire n5580;
   wire n5581;
   wire n5582;
   wire n5583;
   wire n5584;
   wire n5585;
   wire n5586;
   wire n5587;
   wire n5588;
   wire n5589;
   wire n5590;
   wire n5591;
   wire n5592;
   wire n5593;
   wire n5594;
   wire n5595;
   wire n5596;
   wire n5597;
   wire n5598;
   wire n5599;
   wire n5600;
   wire n5601;
   wire n5602;
   wire n5603;
   wire n5604;
   wire n5605;
   wire n5606;
   wire n5607;
   wire n5608;
   wire n5609;
   wire n5610;
   wire n5611;
   wire n5612;
   wire n5613;
   wire n5614;
   wire n5615;
   wire n5616;
   wire n5617;
   wire n5618;
   wire n5619;
   wire n5620;
   wire n5621;
   wire n5622;
   wire n5623;
   wire n5624;
   wire n5625;
   wire n5626;
   wire n5627;
   wire n5628;
   wire n5629;
   wire n5630;
   wire n5631;
   wire n5632;
   wire n5633;
   wire n5634;
   wire n5635;
   wire n5636;
   wire n5637;
   wire n5638;
   wire n5639;
   wire n5640;
   wire n5641;
   wire n5642;
   wire n5643;
   wire n5644;
   wire n5645;
   wire n5646;
   wire n5647;
   wire n5648;
   wire n5649;
   wire n5650;
   wire n5651;
   wire n5652;
   wire n5653;
   wire n5654;
   wire n5655;
   wire n5656;
   wire n5657;
   wire n5658;
   wire n5659;
   wire n5660;
   wire n5661;
   wire n5662;
   wire n5663;
   wire n5664;
   wire n5665;
   wire n5666;
   wire n5667;
   wire n5668;
   wire n5669;
   wire n5670;
   wire n5671;
   wire n5672;
   wire n5673;
   wire n5674;
   wire n5675;
   wire n5676;
   wire n5677;
   wire n5678;
   wire n5679;
   wire n5680;
   wire n5681;
   wire n5682;
   wire n5683;
   wire n5684;
   wire n5685;
   wire n5686;
   wire n5687;
   wire n5688;
   wire n5689;
   wire n5690;
   wire n5691;
   wire n5692;
   wire n5693;
   wire n5694;
   wire n5695;
   wire n5696;
   wire n5697;
   wire n5698;
   wire n5699;
   wire n5700;
   wire n5701;
   wire n5702;
   wire n5703;
   wire n5704;
   wire n5705;
   wire n5706;
   wire n5707;
   wire n5708;
   wire n5709;
   wire n5710;
   wire n5711;
   wire n5712;
   wire n5713;
   wire n5715;
   wire n5716;
   wire n5717;
   wire n5718;
   wire n5719;
   wire n5720;
   wire n5721;
   wire n5722;
   wire n5723;
   wire n5724;
   wire n5725;
   wire n5726;
   wire n5727;
   wire n5728;
   wire n5729;
   wire n5730;
   wire n5731;
   wire n5732;
   wire n5733;
   wire n5734;
   wire n5735;
   wire n5736;
   wire n5737;
   wire n5738;
   wire n5739;
   wire n5740;
   wire n5741;
   wire n5742;
   wire n5743;
   wire n5744;
   wire n5745;
   wire n5746;
   wire n5747;
   wire n5749;
   wire n5750;
   wire n5751;
   wire n5752;
   wire n5753;
   wire n5754;
   wire n5755;
   wire n5756;
   wire n5757;
   wire n5759;
   wire n5760;
   wire n5761;
   wire n5762;
   wire n5763;
   wire n5764;
   wire n5765;
   wire n5766;
   wire n5767;
   wire n5768;
   wire n5769;
   wire n5771;
   wire n5772;
   wire n5773;
   wire n5774;
   wire n5775;
   wire n5776;
   wire n5778;
   wire n5779;
   wire n5780;
   wire n5781;
   wire n5782;
   wire n5783;
   wire n5784;
   wire n5785;
   wire n5786;
   wire n5788;
   wire n5789;
   wire n5790;
   wire n5791;
   wire n5792;
   wire n5793;
   wire n5794;
   wire n5795;
   wire n5796;
   wire n5797;
   wire n5798;
   wire n5799;
   wire n5801;
   wire n5802;
   wire n5803;
   wire n5804;
   wire n5805;
   wire n5806;
   wire n5807;
   wire n5808;
   wire n5809;
   wire n5810;
   wire n5811;
   wire n5812;
   wire n5814;
   wire n5815;
   wire n5816;
   wire n5817;
   wire n5818;
   wire n5819;
   wire n5820;
   wire n5821;
   wire n5822;
   wire n5823;
   wire n5824;
   wire n5825;
   wire n5826;
   wire n5827;
   wire n5828;
   wire n5829;
   wire n5830;
   wire n5831;
   wire n5832;
   wire n5833;
   wire n5834;
   wire n5835;
   wire n5836;
   wire n5837;
   wire n5838;
   wire n5840;
   wire n5841;
   wire n5842;
   wire n5843;
   wire n5844;
   wire n5845;
   wire n5846;
   wire n5847;
   wire n5848;
   wire n5849;
   wire n5850;
   wire n5851;
   wire n5852;
   wire n5853;
   wire n5854;
   wire n5855;
   wire n5856;
   wire n5857;
   wire n5858;
   wire n5859;
   wire n5860;
   wire n5861;
   wire n5862;
   wire n5863;
   wire n5864;
   wire n5865;
   wire n5866;
   wire n5867;
   wire n5868;
   wire n5869;
   wire n5870;
   wire n5871;
   wire n5872;
   wire n5873;
   wire n5874;
   wire n5875;
   wire n5876;
   wire n5877;
   wire n5878;
   wire n5879;
   wire n5880;
   wire n5881;
   wire n5882;
   wire n5883;
   wire n5884;
   wire n5885;
   wire n5886;
   wire n5887;
   wire n5888;
   wire n5889;
   wire n5890;
   wire n5891;
   wire n5892;
   wire n5893;
   wire n5894;
   wire n5895;
   wire n5896;
   wire n5897;
   wire n5898;
   wire n5899;
   wire n5900;
   wire n5901;
   wire n5902;
   wire n5903;
   wire n5904;
   wire n5905;
   wire n5906;
   wire n5907;
   wire n5908;
   wire n5909;
   wire n5910;
   wire n5911;
   wire n5912;
   wire n5913;
   wire n5914;
   wire n5915;
   wire n5916;
   wire n5917;
   wire n5918;
   wire n5919;
   wire n5920;
   wire n5921;
   wire n5922;
   wire n5923;
   wire n5924;
   wire n5925;
   wire n5926;
   wire n5927;
   wire n5928;
   wire n5929;
   wire n5930;
   wire n5931;
   wire n5932;
   wire n5933;
   wire n5934;
   wire n5935;
   wire n5936;
   wire n5937;
   wire n5938;
   wire n5939;
   wire n5940;
   wire n5941;
   wire n5942;
   wire n5943;
   wire n5944;
   wire n5945;
   wire n5946;
   wire n5947;
   wire n5948;
   wire n5949;
   wire n5950;
   wire n5951;
   wire n5952;
   wire n5953;
   wire n5954;
   wire n5955;
   wire n5956;
   wire n5957;
   wire n5958;
   wire n5959;
   wire n5960;
   wire n5961;
   wire n5962;
   wire n5963;
   wire n5964;
   wire n5965;
   wire n5966;
   wire n5967;
   wire n5968;
   wire n5969;
   wire n5970;
   wire n5971;
   wire n5972;
   wire n5973;
   wire n5974;
   wire n5975;
   wire n5976;
   wire n5977;
   wire n5978;
   wire n5979;
   wire n5980;
   wire n5981;
   wire n5982;
   wire n5983;
   wire n5984;
   wire n5985;
   wire n5986;
   wire n5987;
   wire n5988;
   wire n5989;
   wire n5990;
   wire n5991;
   wire n5992;
   wire n5993;
   wire n5994;
   wire n5995;
   wire n5996;
   wire n5997;
   wire n5998;
   wire n5999;
   wire n6000;
   wire n6001;
   wire n6002;
   wire n6003;
   wire n6004;
   wire n6005;
   wire n6006;
   wire n6007;
   wire n6008;
   wire n6009;
   wire n6010;
   wire n6011;
   wire n6012;
   wire n6013;
   wire n6014;
   wire n6015;
   wire n6016;
   wire n6017;
   wire n6018;
   wire n6019;
   wire n6020;
   wire n6021;
   wire n6022;
   wire n6023;
   wire n6024;
   wire n6025;
   wire n6026;
   wire n6027;
   wire n6028;
   wire n6029;
   wire n6030;
   wire n6031;
   wire n6032;
   wire n6033;
   wire n6034;
   wire n6035;
   wire n6036;
   wire n6037;
   wire n6038;
   wire n6039;
   wire n6040;
   wire n6041;
   wire n6042;
   wire n6043;
   wire n6044;
   wire n6045;
   wire n6046;
   wire n6048;
   wire n6050;
   wire n6051;
   wire n6052;
   wire n6053;
   wire n6054;
   wire n6055;
   wire n6056;
   wire n6057;
   wire n6058;
   wire n6059;
   wire n6060;
   wire n6061;
   wire n6062;
   wire n6063;
   wire n6064;
   wire n6065;
   wire n6066;
   wire n6067;
   wire n6068;
   wire n6069;
   wire n6070;
   wire n6073;
   wire n6074;
   wire n6075;
   wire n6076;
   wire n6077;
   wire n6078;
   wire n6079;
   wire n6080;
   wire n6081;
   wire n6082;
   wire n6083;
   wire n6084;
   wire n6085;
   wire n6086;
   wire n6087;
   wire n6088;
   wire n6089;
   wire n6090;
   wire n6091;
   wire n6092;
   wire n6093;
   wire n6094;
   wire n6095;
   wire n6096;
   wire n6097;
   wire n6098;
   wire n6099;
   wire n6100;
   wire n6101;
   wire n6102;
   wire n6103;
   wire n6104;
   wire n6105;
   wire n6106;
   wire n6107;
   wire n6108;
   wire n6109;
   wire n6110;
   wire n6111;
   wire n6112;
   wire n6113;
   wire n6114;
   wire n6115;
   wire n6116;
   wire n6117;
   wire n6118;
   wire n6119;
   wire n6120;
   wire n6121;
   wire n6122;
   wire n6123;
   wire n6124;
   wire n6126;
   wire n6127;
   wire n6128;
   wire n6129;
   wire n6130;
   wire n6131;
   wire n6132;
   wire n6133;
   wire n6134;
   wire n6135;
   wire n6136;
   wire n6137;
   wire n6138;
   wire n6139;
   wire n6140;
   wire n6141;
   wire n6142;
   wire n6143;
   wire n6144;
   wire n6145;
   wire n6146;
   wire n6147;
   wire n6148;
   wire n6149;
   wire n6150;
   wire n6151;
   wire n6152;
   wire n6153;
   wire n6154;
   wire n6155;
   wire n6156;
   wire n6157;
   wire n6158;
   wire n6159;
   wire n6160;
   wire n6161;
   wire n6162;
   wire n6163;
   wire n6164;
   wire n6165;
   wire n6166;
   wire n6167;
   wire n6168;
   wire n6169;
   wire n6170;
   wire n6172;
   wire n6173;
   wire n6174;
   wire n6175;
   wire n6176;
   wire n6177;
   wire n6178;
   wire n6179;
   wire n6180;
   wire n6181;
   wire n6182;
   wire n6183;
   wire n6184;
   wire n6185;
   wire n6186;
   wire n6187;
   wire n6188;
   wire n6189;
   wire n6190;
   wire n6191;
   wire n6192;
   wire n6193;
   wire n6194;
   wire n6195;
   wire n6197;
   wire n6198;
   wire n6199;
   wire n6200;
   wire n6201;
   wire n6202;
   wire n6203;
   wire n6204;
   wire n6205;
   wire n6206;
   wire n6207;
   wire n6208;
   wire n6209;
   wire n6210;
   wire n6211;
   wire n6212;
   wire n6213;
   wire n6214;
   wire n6215;
   wire n6216;
   wire n6217;
   wire n6218;
   wire n6219;
   wire n6220;
   wire n6221;
   wire n6222;
   wire n6223;
   wire n6224;
   wire n6225;
   wire n6226;
   wire n6227;
   wire n6228;
   wire n6229;
   wire n6230;
   wire n6231;
   wire n6232;
   wire n6233;
   wire n6234;
   wire n6235;
   wire n6236;
   wire n6237;
   wire n6238;
   wire n6239;
   wire n6240;
   wire n6241;
   wire n6242;
   wire n6243;
   wire n6244;
   wire n6245;
   wire n6246;
   wire n6247;
   wire n6248;
   wire n6249;
   wire n6250;
   wire n6251;
   wire n6252;
   wire n6253;
   wire n6254;
   wire n6255;
   wire n6256;
   wire n6257;
   wire n6258;
   wire n6259;
   wire n6260;
   wire n6261;
   wire n6262;
   wire n6263;
   wire n6264;
   wire n6265;
   wire n6266;
   wire n6267;
   wire n6268;
   wire n6269;
   wire n6270;
   wire n6271;
   wire n6272;
   wire n6273;
   wire n6274;
   wire n6275;
   wire n6276;
   wire n6277;
   wire n6278;
   wire n6279;
   wire n6280;
   wire n6281;
   wire n6282;
   wire n6283;
   wire n6284;
   wire n6285;
   wire n6286;
   wire n6287;
   wire n6288;
   wire n6289;
   wire n6291;
   wire n6292;
   wire n6293;
   wire n6294;
   wire n6296;
   wire n6297;
   wire n6298;
   wire n6299;
   wire n6300;
   wire n6301;
   wire n6302;
   wire n6303;
   wire n6304;
   wire n6305;
   wire n6306;
   wire n6307;
   wire n6308;
   wire n6309;
   wire n6310;
   wire n6311;
   wire n6312;
   wire n6313;
   wire n6314;
   wire n6315;
   wire n6316;
   wire n6317;
   wire n6318;
   wire n6319;
   wire n6320;
   wire n6321;
   wire n6322;
   wire n6323;
   wire n6324;
   wire n6325;
   wire n6326;
   wire n6327;
   wire n6328;
   wire n6329;
   wire n6330;
   wire n6331;
   wire n6332;
   wire n6333;
   wire n6334;
   wire n6335;
   wire n6336;
   wire n6337;
   wire n6338;
   wire n6339;
   wire n6340;
   wire n6341;
   wire n6342;
   wire n6343;
   wire n6344;
   wire n6345;
   wire n6347;
   wire n6348;
   wire n6349;
   wire n6350;
   wire n6351;
   wire n6352;
   wire n6353;
   wire n6354;
   wire n6355;
   wire n6356;
   wire net54953;
   wire net54895;
   wire net54893;
   wire net54891;
   wire net54889;
   wire net54887;
   wire net54885;
   wire net54883;
   wire net54881;
   wire net54879;
   wire net54877;
   wire net54875;
   wire net54873;
   wire net54871;
   wire net54869;
   wire net54867;
   wire net54865;
   wire net54863;
   wire net54861;
   wire net54859;
   wire net54857;
   wire net54855;
   wire net54853;
   wire net54851;
   wire net54849;
   wire net54847;
   wire net54845;
   wire net54843;
   wire net56414;
   wire net87679;
   wire n6369;
   wire n6370;
   wire n6371;
   wire n6373;
   wire n6374;
   wire n6375;
   wire n6376;
   wire n6380;
   wire n6381;
   wire n6382;
   wire n6383;
   wire n6384;
   wire n6385;
   wire n6386;
   wire n6387;
   wire n6388;
   wire n6389;
   wire n6390;
   wire n6391;
   wire n6392;
   wire n6393;
   wire n6394;
   wire n6395;
   wire n6396;
   wire n6397;
   wire n6398;
   wire n6399;
   wire n6400;
   wire n6401;
   wire n6402;
   wire n6403;
   wire n6404;
   wire n6405;
   wire n6406;
   wire n6407;
   wire n6408;
   wire n6410;
   wire n6411;
   wire n6412;
   wire n6413;
   wire n6414;
   wire n6415;
   wire n6416;
   wire n6417;
   wire n6418;
   wire n6419;
   wire n6420;
   wire n6421;
   wire n6422;
   wire n6423;
   wire n6424;
   wire n6425;
   wire n6426;
   wire n6428;
   wire n6429;
   wire n6430;
   wire n6431;
   wire n6432;
   wire n6433;
   wire n6434;
   wire n6435;
   wire n6436;
   wire n6437;
   wire n6438;
   wire n6439;
   wire n6440;
   wire n6443;
   wire n6444;
   wire n6445;
   wire n6447;
   wire n6449;
   wire n6451;
   wire n6454;
   wire n6455;
   wire n6456;
   wire n6457;
   wire n6458;
   wire n6459;
   wire n6460;
   wire n6461;
   wire n6462;
   wire n6463;
   wire n6465;
   wire n6466;
   wire n6467;
   wire n6468;
   wire n6469;
   wire n6470;
   wire n6471;
   wire n6472;
   wire n6473;
   wire n6474;
   wire n6476;
   wire n6477;
   wire n6478;
   wire n6479;
   wire n6480;
   wire n6481;
   wire n6482;
   wire n6483;
   wire n6484;
   wire n6487;
   wire n6488;
   wire n6489;
   wire n6490;
   wire n6491;
   wire n6492;
   wire n6493;
   wire n6494;
   wire n6495;
   wire n6496;
   wire n6497;
   wire n6498;
   wire n6499;
   wire n6500;
   wire n6501;
   wire n6502;
   wire n6504;
   wire n6505;
   wire n6506;
   wire n6507;
   wire n6508;
   wire n6509;
   wire n6510;
   wire n6511;
   wire n6512;
   wire n6513;
   wire n6514;
   wire n6515;
   wire n6516;
   wire n6519;
   wire n6520;
   wire n6521;
   wire n6522;
   wire n6523;
   wire n6524;
   wire n6526;
   wire n6527;
   wire n6528;
   wire n6529;
   wire n6530;
   wire n6531;
   wire n6532;
   wire n6533;
   wire n6534;
   wire n6535;
   wire n6536;
   wire n6537;
   wire n6538;
   wire n6543;
   wire n6544;
   wire n6545;
   wire n6546;
   wire n6547;
   wire n6548;
   wire n6549;
   wire n6550;
   wire n6551;
   wire n6552;
   wire n6553;
   wire n6554;
   wire n6555;
   wire n6556;
   wire n6558;
   wire n6559;
   wire n6560;
   wire n6561;
   wire n6562;
   wire n6563;
   wire n6564;
   wire n6565;
   wire n6566;
   wire n6567;
   wire n6568;
   wire n6569;
   wire n6570;
   wire n6571;
   wire n6572;
   wire n6573;
   wire n6575;
   wire n6576;
   wire n6577;
   wire n6578;
   wire n6579;
   wire n6580;
   wire n6581;
   wire n6582;
   wire n6583;
   wire n6584;
   wire n6585;
   wire n6586;
   wire n6587;
   wire n6589;
   wire n6590;
   wire n6591;
   wire n6592;
   wire n6593;
   wire n6594;
   wire n6595;
   wire n6596;
   wire n6597;
   wire n6598;
   wire n6599;
   wire n6600;
   wire n6601;
   wire n6602;
   wire n6603;
   wire n6604;
   wire n6605;
   wire n6606;
   wire n6607;
   wire n6608;
   wire n6609;
   wire n6610;
   wire n6611;
   wire n6612;
   wire n6613;
   wire n6614;
   wire n6615;
   wire n6616;
   wire n6617;
   wire n6618;
   wire n6619;
   wire n6621;
   wire n6623;
   wire n6624;
   wire n6626;
   wire n6627;
   wire n6628;
   wire n6629;
   wire n6630;
   wire n6631;
   wire n6632;
   wire n6633;
   wire n6634;
   wire n6635;
   wire n6636;
   wire n6637;
   wire n6640;
   wire n6641;
   wire n6642;
   wire n6644;
   wire n6647;
   wire n6648;
   wire n6649;
   wire n6650;
   wire n6651;
   wire n6652;
   wire n6653;
   wire n6654;
   wire n6655;
   wire n6657;
   wire n6660;
   wire n6661;
   wire n6662;
   wire n6663;
   wire n6664;
   wire n6665;
   wire n6666;
   wire n6667;
   wire n6668;
   wire n6669;
   wire n6670;
   wire n6671;
   wire n6672;
   wire n6673;
   wire n6676;
   wire n6677;
   wire n6680;
   wire n6681;
   wire n6682;
   wire n6684;
   wire n6685;
   wire n6686;
   wire n6687;
   wire n6688;
   wire n6689;
   wire n6690;
   wire n6691;
   wire n6692;
   wire n6693;
   wire n6694;
   wire n6695;
   wire n6696;
   wire n6697;
   wire n6699;
   wire n6700;
   wire n6703;
   wire n6704;
   wire n6705;
   wire n6707;
   wire n6708;
   wire n6709;
   wire n6711;
   wire n6712;
   wire n6714;
   wire n6717;
   wire n6718;
   wire n6719;
   wire n6720;
   wire n6721;
   wire n6723;
   wire n6724;
   wire n6725;
   wire n6726;
   wire n6727;
   wire n6728;
   wire n6729;
   wire n6730;
   wire n6731;
   wire n6732;
   wire n6733;
   wire n6734;
   wire n6735;
   wire n6736;
   wire n6737;
   wire n6740;
   wire n6741;
   wire n6742;
   wire n6744;
   wire n6745;
   wire n6746;
   wire n6747;
   wire n6748;
   wire n6749;
   wire n6750;
   wire n6751;
   wire n6752;
   wire n6754;
   wire n6756;
   wire n6757;
   wire n6759;
   wire n6760;
   wire n6761;
   wire n6763;
   wire n6764;
   wire n6765;
   wire n6767;
   wire n6769;
   wire n6771;
   wire n6772;
   wire n6774;
   wire n6775;
   wire n6776;
   wire n6777;
   wire n6779;
   wire n6781;
   wire n6785;
   wire n6786;
   wire n6787;
   wire n6788;
   wire n6789;
   wire n6790;
   wire n6792;
   wire n6794;
   wire n6796;
   wire n6797;
   wire n6799;
   wire n6801;
   wire n6802;
   wire n6803;
   wire n6804;
   wire n6805;
   wire n6809;
   wire n6813;
   wire n6814;
   wire n6815;
   wire n6816;
   wire n6819;
   wire n6822;
   wire n6824;
   wire n6825;
   wire n6826;
   wire n6829;
   wire n6830;
   wire n6831;
   wire n6832;
   wire n6833;
   wire n6834;
   wire n6836;
   wire n6838;
   wire n6843;
   wire n6844;
   wire n6845;
   wire n6846;
   wire n6848;
   wire n6849;
   wire n6850;
   wire n6851;
   wire n6852;
   wire n6854;
   wire n6855;
   wire n6856;
   wire n6858;
   wire n6859;
   wire n6860;
   wire n6861;
   wire n6862;
   wire n6863;
   wire n6864;
   wire n6865;
   wire n6866;
   wire n6868;
   wire n6870;
   wire n6872;
   wire n6875;
   wire n6876;
   wire n6877;
   wire n6880;
   wire n6881;
   wire n6882;
   wire n6883;
   wire n6885;
   wire n6887;
   wire n6888;
   wire n6889;
   wire n6890;
   wire n6893;
   wire n6894;
   wire n6902;
   wire n6903;
   wire n6904;
   wire n6905;
   wire n6906;
   wire n6907;
   wire n6908;
   wire n6909;
   wire n6910;
   wire n6911;
   wire n6912;
   wire n6913;
   wire n6914;
   wire n6915;
   wire n6916;
   wire n6917;
   wire n6918;
   wire n6919;
   wire n6920;
   wire n6921;
   wire n6922;
   wire n6923;
   wire n6924;
   wire n6925;
   wire n6926;
   wire n6927;
   wire n6928;
   wire n6929;
   wire n6930;
   wire n6931;
   wire n6932;
   wire n6933;
   wire n6934;
   wire n6935;
   wire n6936;
   wire n6937;
   wire n6938;
   wire n6939;
   wire [31:0] I_DATA_INBUS;
   wire [31:0] D_ADDR_OUTBUS;
   wire [31:0] D_DATA_OUTBUS;
   wire [12:2] dram_addr_outbus;
   wire [31:0] dram_data_inbus;
   wire [31:0] dram_data_outbus;
   wire [31:0] d_select;
   wire [5:0] \UUT/d_mul_command ;
   wire [2:0] \UUT/exe_outsel ;
   wire [2:0] \UUT/shift_op ;
   wire [23:0] \UUT/jar_in ;
   wire [31:0] \UUT/branch_regb ;
   wire [31:0] \UUT/branch_rega ;
   wire [4:0] \UUT/rd_addr ;
   wire [4:0] \UUT/rs2_addr ;
   wire [4:0] \UUT/rs1_addr ;
   wire [31:0] \UUT/daddr_out ;
   wire [5:0] \UUT/Mcontrol/x_mul_command ;
   wire [31:0] \UUT/Mcontrol/d_instr ;
   wire [31:0] \UUT/Mcontrol/d_sampled_finstr ;
   wire [23:0] \UUT/Mcontrol/f_currpc ;
   wire [23:0] \UUT/Mcontrol/Nextpc_decoding/Bta ;
   wire [1:0] \UUT/Mpath/mem_baddr ;
   wire [31:0] \UUT/Mpath/the_shift/sh_sll ;
   wire [31:0] \UUT/Mpath/the_shift/sh_srl ;
   wire [31:0] \UUT/Mpath/the_shift/sh_sra ;
   wire [31:0] \UUT/Mpath/the_shift/sh_ror ;
   wire [31:0] \UUT/Mpath/the_shift/sh_rol ;
   wire [63:0] \UUT/Mpath/the_mult/Mad_out ;
   wire [31:0] \UUT/Mpath/the_mult/x_operand2 ;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;

   assign BUS_BUSY = 1'b1 ;
   assign \UUT/Mcontrol/int_reset  = reset ;

   BUF_X8 FE_OFCC208_FE_OFN7_n312 (.Z(FE_OFCN208_FE_OFN7_n312), 
	.A(FE_OFN7_n312));
   BUF_X4 FE_OFCC207_n316 (.Z(FE_OFCN207_n316), 
	.A(n316));
   BUF_X16 FE_OFCC206_FE_OFN186_n546 (.Z(FE_OFCN206_FE_OFN186_n546), 
	.A(FE_OFN186_n546));
   BUF_X8 FE_OFCC205_FE_OFN104_UUT_Mpath_out_regA_0_ (.Z(FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_), 
	.A(FE_OFN104_UUT_Mpath_out_regA_0_));
   BUF_X8 FE_OFCC204_FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_ (.Z(FE_OFCN204_FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_));
   BUF_X8 FE_OFCC203_FE_OFN160_UUT_Mpath_out_regB_4_ (.Z(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_), 
	.A(FE_OFN160_UUT_Mpath_out_regB_4_));
   BUF_X16 FE_OFCC202_FE_OFN164_UUT_Mpath_out_regB_3_ (.Z(FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_), 
	.A(FE_OFN164_UUT_Mpath_out_regB_3_));
   BUF_X16 FE_OFCC201_FE_OFN176_UUT_Mpath_out_regB_1_ (.Z(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.A(FE_OFN176_UUT_Mpath_out_regB_1_));
   BUF_X8 FE_OFCC200_FE_OFN175_UUT_Mpath_out_regB_1_ (.Z(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_), 
	.A(FE_OFN175_UUT_Mpath_out_regB_1_));
   BUF_X4 FE_OFCC199_UUT_rs1_addr_3_ (.Z(FE_OFCN199_UUT_rs1_addr_3_), 
	.A(\UUT/rs1_addr [3]));
   BUF_X8 FE_OFCC198_UUT_Mpath_out_regA_2_ (.Z(FE_OFCN198_UUT_Mpath_out_regA_2_), 
	.A(\UUT/Mpath/out_regA[2] ));
   CLKBUF_X1 FE_OFC197_n741 (.Z(FE_OFN197_n741), 
	.A(n741));
   CLKBUF_X1 FE_OFC196_n764 (.Z(FE_OFN196_n764), 
	.A(n764));
   CLKBUF_X1 FE_OFC195_n5438 (.Z(FE_OFN195_n5438), 
	.A(n5438));
   CLKBUF_X1 FE_OFC194_n5429 (.Z(FE_OFN194_n5429), 
	.A(n5429));
   CLKBUF_X1 FE_OFC193_n5522 (.Z(FE_OFN193_n5522), 
	.A(n5522));
   CLKBUF_X1 FE_OFC192_n208 (.Z(FE_OFN192_n208), 
	.A(n208));
   CLKBUF_X1 FE_OFC191_n5435 (.Z(FE_OFN191_n5435), 
	.A(n5435));
   CLKBUF_X1 FE_OFC190_n5447 (.Z(FE_OFN190_n5447), 
	.A(n5447));
   CLKBUF_X1 FE_OFC189_n5459 (.Z(FE_OFN189_n5459), 
	.A(n5459));
   CLKBUF_X1 FE_OFC188_n5492 (.Z(FE_OFN188_n5492), 
	.A(n5492));
   CLKBUF_X1 FE_OFC187_UUT_branch_rega_1_ (.Z(FE_OFN187_UUT_branch_rega_1_), 
	.A(\UUT/branch_rega [1]));
   CLKBUF_X2 FE_OFC186_n546 (.Z(FE_OFN186_n546), 
	.A(n546));
   BUF_X4 FE_OFC185_UUT_Mpath_out_regB_0_ (.Z(FE_OFN185_UUT_Mpath_out_regB_0_), 
	.A(FE_OFN182_UUT_Mpath_out_regB_0_));
   CLKBUF_X1 FE_OFC184_UUT_Mpath_out_regB_0_ (.Z(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.A(FE_OFN182_UUT_Mpath_out_regB_0_));
   BUF_X4 FE_OFC182_UUT_Mpath_out_regB_0_ (.Z(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.A(\UUT/Mpath/out_regB[0] ));
   BUF_X1 FE_OFC177_UUT_Mpath_the_mult_x_operand1_31_ (.Z(FE_OFN177_UUT_Mpath_the_mult_x_operand1_31_), 
	.A(\UUT/Mpath/the_mult/x_operand1[31] ));
   CLKBUF_X3 FE_OFC176_UUT_Mpath_out_regB_1_ (.Z(FE_OFN176_UUT_Mpath_out_regB_1_), 
	.A(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_));
   CLKBUF_X3 FE_OFC175_UUT_Mpath_out_regB_1_ (.Z(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.A(\UUT/Mpath/out_regB[1] ));
   CLKBUF_X2 FE_OFC173_UUT_Mpath_the_mult_x_operand1_23_ (.Z(FE_OFN173_UUT_Mpath_the_mult_x_operand1_23_), 
	.A(\UUT/Mpath/the_mult/x_operand1[23] ));
   BUF_X1 FE_OFC171_UUT_Mpath_the_mult_x_operand1_1_ (.Z(FE_OFN171_UUT_Mpath_the_mult_x_operand1_1_), 
	.A(\UUT/Mpath/the_mult/x_operand1[1] ));
   CLKBUF_X2 FE_OFC170_UUT_Mpath_the_mult_x_operand2_1_ (.Z(FE_OFN170_UUT_Mpath_the_mult_x_operand2_1_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [1]));
   CLKBUF_X3 FE_OFC169_UUT_Mpath_out_regB_2_ (.Z(FE_OFN169_UUT_Mpath_out_regB_2_), 
	.A(FE_OFN168_UUT_Mpath_out_regB_2_));
   BUF_X4 FE_OFC168_UUT_Mpath_out_regB_2_ (.Z(FE_OFN168_UUT_Mpath_out_regB_2_), 
	.A(\UUT/Mpath/out_regB[2] ));
   CLKBUF_X2 FE_OFC167_UUT_Mpath_the_mult_x_operand2_2_ (.Z(FE_OFN167_UUT_Mpath_the_mult_x_operand2_2_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [2]));
   BUF_X2 FE_OFC165_UUT_Mpath_the_mult_x_operand1_3_ (.Z(FE_OFN165_UUT_Mpath_the_mult_x_operand1_3_), 
	.A(\UUT/Mpath/the_mult/x_operand1[3] ));
   CLKBUF_X3 FE_OFC164_UUT_Mpath_out_regB_3_ (.Z(FE_OFN164_UUT_Mpath_out_regB_3_), 
	.A(FE_OFN163_UUT_Mpath_out_regB_3_));
   CLKBUF_X3 FE_OFC163_UUT_Mpath_out_regB_3_ (.Z(FE_OFN163_UUT_Mpath_out_regB_3_), 
	.A(FE_OFN162_UUT_Mpath_out_regB_3_));
   CLKBUF_X3 FE_OFC162_UUT_Mpath_out_regB_3_ (.Z(FE_OFN162_UUT_Mpath_out_regB_3_), 
	.A(\UUT/Mpath/out_regB[3] ));
   CLKBUF_X3 FE_OFC160_UUT_Mpath_out_regB_4_ (.Z(FE_OFN160_UUT_Mpath_out_regB_4_), 
	.A(FE_OFN159_UUT_Mpath_out_regB_4_));
   BUF_X4 FE_OFC159_UUT_Mpath_out_regB_4_ (.Z(FE_OFN159_UUT_Mpath_out_regB_4_), 
	.A(\UUT/Mpath/out_regB[4] ));
   BUF_X1 FE_OFC156_UUT_Mpath_the_mult_x_operand1_5_ (.Z(FE_OFN156_UUT_Mpath_the_mult_x_operand1_5_), 
	.A(\UUT/Mpath/the_mult/x_operand1[5] ));
   BUF_X1 FE_OFC152_UUT_Mpath_the_mult_x_operand1_7_ (.Z(FE_OFN152_UUT_Mpath_the_mult_x_operand1_7_), 
	.A(\UUT/Mpath/the_mult/x_operand1[7] ));
   BUF_X1 FE_OFC149_UUT_Mpath_the_mult_x_operand1_9_ (.Z(FE_OFN149_UUT_Mpath_the_mult_x_operand1_9_), 
	.A(\UUT/Mpath/the_mult/x_operand1[9] ));
   BUF_X1 FE_OFC146_UUT_Mpath_the_mult_x_operand1_11_ (.Z(FE_OFN146_UUT_Mpath_the_mult_x_operand1_11_), 
	.A(\UUT/Mpath/the_mult/x_operand1[11] ));
   BUF_X1 FE_OFC142_UUT_Mpath_the_mult_x_operand1_13_ (.Z(FE_OFN142_UUT_Mpath_the_mult_x_operand1_13_), 
	.A(\UUT/Mpath/the_mult/x_operand1[13] ));
   CLKBUF_X2 FE_OFC140_UUT_Mpath_the_mult_x_operand2_14_ (.Z(FE_OFN140_UUT_Mpath_the_mult_x_operand2_14_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [14]));
   BUF_X1 FE_OFC138_UUT_Mpath_the_mult_x_operand1_15_ (.Z(FE_OFN138_UUT_Mpath_the_mult_x_operand1_15_), 
	.A(\UUT/Mpath/the_mult/x_operand1[15] ));
   CLKBUF_X2 FE_OFC137_UUT_Mpath_the_mult_x_operand2_15_ (.Z(FE_OFN137_UUT_Mpath_the_mult_x_operand2_15_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [15]));
   CLKBUF_X2 FE_OFC136_UUT_Mpath_the_mult_x_operand2_16_ (.Z(FE_OFN136_UUT_Mpath_the_mult_x_operand2_16_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [16]));
   BUF_X2 FE_OFC134_UUT_Mpath_the_mult_x_operand1_17_ (.Z(FE_OFN134_UUT_Mpath_the_mult_x_operand1_17_), 
	.A(\UUT/Mpath/the_mult/x_operand1[17] ));
   CLKBUF_X2 FE_OFC133_UUT_Mpath_the_mult_x_operand2_17_ (.Z(FE_OFN133_UUT_Mpath_the_mult_x_operand2_17_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [17]));
   BUF_X2 FE_OFC130_UUT_Mpath_the_mult_x_operand1_19_ (.Z(FE_OFN130_UUT_Mpath_the_mult_x_operand1_19_), 
	.A(\UUT/Mpath/the_mult/x_operand1[19] ));
   CLKBUF_X2 FE_OFC129_UUT_Mpath_the_mult_x_operand2_19_ (.Z(FE_OFN129_UUT_Mpath_the_mult_x_operand2_19_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [19]));
   BUF_X1 FE_OFC126_UUT_Mpath_the_mult_x_operand1_21_ (.Z(FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_), 
	.A(\UUT/Mpath/the_mult/x_operand1[21] ));
   BUF_X2 FE_OFC121_UUT_Mpath_the_mult_x_operand1_25_ (.Z(FE_OFN121_UUT_Mpath_the_mult_x_operand1_25_), 
	.A(\UUT/Mpath/the_mult/x_operand1[25] ));
   CLKBUF_X2 FE_OFC120_UUT_Mpath_the_mult_x_operand2_25_ (.Z(FE_OFN120_UUT_Mpath_the_mult_x_operand2_25_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [25]));
   BUF_X2 FE_OFC117_UUT_Mpath_the_mult_x_operand1_27_ (.Z(FE_OFN117_UUT_Mpath_the_mult_x_operand1_27_), 
	.A(\UUT/Mpath/the_mult/x_operand1[27] ));
   BUF_X2 FE_OFC113_UUT_Mpath_the_mult_x_operand1_29_ (.Z(FE_OFN113_UUT_Mpath_the_mult_x_operand1_29_), 
	.A(\UUT/Mpath/the_mult/x_operand1[29] ));
   BUF_X2 FE_OFC105_UUT_Mpath_the_mult_x_operand2_0_ (.Z(FE_OFN105_UUT_Mpath_the_mult_x_operand2_0_), 
	.A(\UUT/Mpath/the_mult/x_operand2 [0]));
   CLKBUF_X1 FE_OFC104_UUT_Mpath_out_regA_0_ (.Z(FE_OFN104_UUT_Mpath_out_regA_0_), 
	.A(\UUT/Mpath/out_regA[0] ));
   CLKBUF_X1 FE_OFC103_UUT_Mcontrol_Nextpc_decoding_N255 (.Z(FE_OFN103_UUT_Mcontrol_Nextpc_decoding_N255), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N255 ));
   CLKBUF_X1 FE_OFC102_n117 (.Z(FE_OFN102_n117), 
	.A(n117));
   CLKBUF_X1 FE_OFC101_n292 (.Z(FE_OFN101_n292), 
	.A(n292));
   CLKBUF_X1 FE_OFC100_n327 (.Z(FE_OFN100_n327), 
	.A(n327));
   CLKBUF_X1 FE_OFC99_n348 (.Z(FE_OFN99_n348), 
	.A(n348));
   CLKBUF_X1 FE_OFC98_UUT_rs1_addr_1_ (.Z(FE_OFN98_UUT_rs1_addr_1_), 
	.A(\UUT/rs1_addr [1]));
   CLKBUF_X2 FE_OFC97_n5529 (.Z(FE_OFN97_n5529), 
	.A(n5529));
   CLKBUF_X2 FE_OFC96_n5530 (.Z(FE_OFN96_n5530), 
	.A(n5530));
   CLKBUF_X1 FE_OFC95_n2409 (.Z(FE_OFN95_n2409), 
	.A(n2409));
   CLKBUF_X1 FE_OFC94_n2455 (.Z(FE_OFN94_n2455), 
	.A(n2455));
   CLKBUF_X1 FE_OFC93_n1878 (.Z(FE_OFN93_n1878), 
	.A(n1878));
   CLKBUF_X2 FE_OFC92_n5780 (.Z(FE_OFN92_n5780), 
	.A(n5780));
   CLKBUF_X2 FE_OFC91_n285 (.Z(FE_OFN91_n285), 
	.A(n285));
   CLKBUF_X2 FE_OFC90_n325 (.Z(FE_OFN90_n325), 
	.A(n325));
   CLKBUF_X2 FE_OFC89_n290 (.Z(FE_OFN89_n290), 
	.A(n290));
   CLKBUF_X2 FE_OFC88_n6201 (.Z(FE_OFN88_n6201), 
	.A(n6201));
   CLKBUF_X2 FE_OFC87_n1211 (.Z(FE_OFN87_n1211), 
	.A(n1211));
   CLKBUF_X2 FE_OFC86_n1214 (.Z(FE_OFN86_n1214), 
	.A(n1214));
   CLKBUF_X1 FE_OFC85_n2173 (.Z(FE_OFN85_n2173), 
	.A(n2173));
   CLKBUF_X1 FE_OFC84_n1498 (.Z(FE_OFN84_n1498), 
	.A(n1498));
   CLKBUF_X1 FE_OFC83_n2340 (.Z(FE_OFN83_n2340), 
	.A(n2340));
   CLKBUF_X1 FE_OFC82_n1718 (.Z(FE_OFN82_n1718), 
	.A(n1718));
   CLKBUF_X1 FE_OFC80_n2581 (.Z(FE_OFN80_n2581), 
	.A(n2581));
   CLKBUF_X1 FE_OFC79_n1778 (.Z(FE_OFN79_n1778), 
	.A(n1778));
   CLKBUF_X1 FE_OFC77_n2547 (.Z(FE_OFN77_n2547), 
	.A(n2547));
   CLKBUF_X1 FE_OFC76_n1798 (.Z(FE_OFN76_n1798), 
	.A(n1798));
   CLKBUF_X1 FE_OFC74_n2525 (.Z(FE_OFN74_n2525), 
	.A(n2525));
   CLKBUF_X1 FE_OFC73_n1818 (.Z(FE_OFN73_n1818), 
	.A(n1818));
   CLKBUF_X1 FE_OFC71_n2501 (.Z(FE_OFN71_n2501), 
	.A(n2501));
   CLKBUF_X1 FE_OFC69_n2478 (.Z(FE_OFN69_n2478), 
	.A(n2478));
   CLKBUF_X1 FE_OFC68_n1858 (.Z(FE_OFN68_n1858), 
	.A(n1858));
   CLKBUF_X1 FE_OFC63_n2386 (.Z(FE_OFN63_n2386), 
	.A(n2386));
   CLKBUF_X1 FE_OFC62_n1318 (.Z(FE_OFN62_n1318), 
	.A(n1318));
   CLKBUF_X1 FE_OFC60_n2363 (.Z(FE_OFN60_n2363), 
	.A(n2363));
   CLKBUF_X1 FE_OFC59_n1338 (.Z(FE_OFN59_n1338), 
	.A(n1338));
   CLKBUF_X1 FE_OFC57_n2313 (.Z(FE_OFN57_n2313), 
	.A(n2313));
   CLKBUF_X1 FE_OFC56_n1358 (.Z(FE_OFN56_n1358), 
	.A(n1358));
   CLKBUF_X1 FE_OFC54_n2293 (.Z(FE_OFN54_n2293), 
	.A(n2293));
   CLKBUF_X1 FE_OFC53_n1378 (.Z(FE_OFN53_n1378), 
	.A(n1378));
   CLKBUF_X1 FE_OFC50_n2253 (.Z(FE_OFN50_n2253), 
	.A(n2253));
   CLKBUF_X1 FE_OFC49_n1418 (.Z(FE_OFN49_n1418), 
	.A(n1418));
   CLKBUF_X1 FE_OFC30_n5450 (.Z(FE_OFN30_n5450), 
	.A(n5450));
   CLKBUF_X1 FE_OFC26_n180 (.Z(FE_OFN26_n180), 
	.A(n180));
   CLKBUF_X1 FE_OFC25_n859 (.Z(FE_OFN25_n859), 
	.A(n859));
   CLKBUF_X1 FE_OFC24_n128 (.Z(FE_OFN24_n128), 
	.A(n128));
   CLKBUF_X1 FE_OFC23_n152 (.Z(FE_OFN23_n152), 
	.A(n152));
   CLKBUF_X1 FE_OFC22_n164 (.Z(FE_OFN22_n164), 
	.A(n164));
   CLKBUF_X1 FE_OFC21_n193 (.Z(FE_OFN21_n193), 
	.A(n193));
   CLKBUF_X1 FE_OFC18_n5441 (.Z(FE_OFN18_n5441), 
	.A(n5441));
   CLKBUF_X1 FE_OFC17_n5444 (.Z(FE_OFN17_n5444), 
	.A(n5444));
   CLKBUF_X1 FE_OFC13_n953 (.Z(FE_OFN13_n953), 
	.A(n953));
   CLKBUF_X3 FE_OFC12_net54953 (.Z(FE_OFN12_net54953), 
	.A(FE_OFN11_net54953));
   CLKBUF_X3 FE_OFC11_net54953 (.Z(FE_OFN11_net54953), 
	.A(net54953));
   CLKBUF_X3 FE_OFC10_net54953 (.Z(FE_OFN10_net54953), 
	.A(net54953));
   CLKBUF_X1 FE_OFC9_n986 (.Z(FE_OFN9_n986), 
	.A(n986));
   CLKBUF_X3 FE_OFC8_n73 (.Z(FE_OFN8_n73), 
	.A(n73));
   CLKBUF_X1 FE_OFC7_n312 (.Z(FE_OFN7_n312), 
	.A(n312));
   CLKBUF_X1 FE_OFC6_n314 (.Z(FE_OFN6_n314), 
	.A(n314));
   CLKBUF_X2 FE_OFC5_n318 (.Z(FE_OFN5_n318), 
	.A(n318));
   CLKBUF_X1 FE_OFC4_n319 (.Z(FE_OFN4_n319), 
	.A(n319));
   CLKBUF_X1 FE_OFC3_n202 (.Z(FE_OFN3_n202), 
	.A(n202));
   CLKBUF_X1 FE_OFC1_n189 (.Z(FE_OFN1_n189), 
	.A(n189));
   CLKBUF_X1 FE_OFC0_n173 (.Z(FE_OFN0_n173), 
	.A(n173));
   SRAM DMem (.address(dram_addr_outbus), 
	.bit_wen(dram_data_outbus), 
	.data_in({ d_select[31],
		d_select[31],
		d_select[31],
		d_select[31],
		d_select[31],
		d_select[31],
		d_select[31],
		d_select[31],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[23],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[9],
		d_select[7],
		d_select[7],
		d_select[7],
		d_select[7],
		d_select[7],
		d_select[7],
		d_select[7],
		d_select[7] }), 
	.data_out(dram_data_inbus), 
	.clk(CLK), 
	.rdn(dram_mr), 
	.wrn(dram_mw));
   SRAM IMem (.address({ n6686,
		n6487,
		\UUT/Mcontrol/Program_counter/N24 ,
		\UUT/Mcontrol/Program_counter/N22 ,
		FE_UNCONNECTED_1,
		n6649,
		n6654,
		n6848,
		n6855,
		n6647,
		FE_UNCONNECTED_0 }), 
	.bit_wen({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.data_in({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.data_out(I_DATA_INBUS), 
	.clk(CLK), 
	.rdn(iram_rd), 
	.wrn(1'b1));
   OR2_X1 \localbus/C745  (.ZN(\localbus/N214 ), 
	.A2(\localbus/N227 ), 
	.A1(\localbus/c1_op[SLAVE][0] ));
   INV_X1 \localbus/I_2  (.ZN(\localbus/N218 ), 
	.A(\localbus/N214 ));
   OR2_X2 \localbus/C756  (.ZN(\localbus/N225 ), 
	.A2(\localbus/N227 ), 
	.A1(n6637));
   INV_X1 \localbus/I_7  (.ZN(\localbus/N229 ), 
	.A(\localbus/N225 ));
   INV_X1 \localbus/I_16  (.ZN(\localbus/N250 ), 
	.A(\localbus/c1_op[OP][0] ));
   OR2_X1 \localbus/C790  (.ZN(\localbus/N251 ), 
	.A2(\localbus/c1_op[OP][1] ), 
	.A1(\localbus/N250 ));
   INV_X1 \localbus/I_17  (.ZN(\localbus/N252 ), 
	.A(\localbus/N251 ));
   INV_X1 \localbus/I_19  (.ZN(\localbus/N256 ), 
	.A(\localbus/c1_op[OP][1] ));
   OR2_X1 \localbus/C796  (.ZN(\localbus/N257 ), 
	.A2(\localbus/N256 ), 
	.A1(\localbus/c1_op[OP][0] ));
   INV_X1 \localbus/I_20  (.ZN(\localbus/N258 ), 
	.A(\localbus/N257 ));
   OR2_X1 \localbus/C881  (.ZN(\localbus/N318 ), 
	.A2(\localbus/c2_op[SLAVE][2] ), 
	.A1(\localbus/c2_op[SLAVE][1] ));
   OR2_X1 \localbus/C882  (.ZN(\localbus/N319 ), 
	.A2(\localbus/N318 ), 
	.A1(\localbus/N219 ));
   INV_X1 \localbus/I_46  (.ZN(\localbus/N320 ), 
	.A(\localbus/N319 ));
   OR2_X1 \localbus/C885  (.ZN(\localbus/N321 ), 
	.A2(\localbus/c2_op[OP][1] ), 
	.A1(\localbus/N293 ));
   INV_X1 \localbus/I_47  (.ZN(\localbus/N322 ), 
	.A(\localbus/N321 ));
   OR2_X1 \localbus/C895  (.ZN(\localbus/N329 ), 
	.A2(\localbus/N318 ), 
	.A1(\localbus/c2_op[SLAVE][0] ));
   INV_X1 \localbus/I_52  (.ZN(\localbus/N335 ), 
	.A(\localbus/N329 ));
   OR2_X1 \localbus/C906  (.ZN(\localbus/N338 ), 
	.A2(\localbus/c1_op[OP][1] ), 
	.A1(\localbus/c1_op[OP][0] ));
   INV_X1 \localbus/I_55  (.ZN(\localbus/c1_op[OP][0] ), 
	.A(dmem_read));
   INV_X1 \localbus/I_56  (.ZN(\localbus/N46 ), 
	.A(dmem_write));
   AND2_X1 \localbus/C959  (.ZN(\localbus/N51 ), 
	.A2(\localbus/N258 ), 
	.A1(\localbus/N50 ));
   AND2_X1 \localbus/C964  (.ZN(\localbus/N57 ), 
	.A2(\localbus/N56 ), 
	.A1(\localbus/N55 ));
   AND2_X1 \localbus/C967  (.ZN(\localbus/N62 ), 
	.A2(\localbus/N61 ), 
	.A1(\localbus/N60 ));
   AND2_X1 \localbus/C983  (.ZN(\localbus/N85 ), 
	.A2(\localbus/N218 ), 
	.A1(\localbus/N252 ));
   AND2_X1 \localbus/C984  (.ZN(\localbus/N86 ), 
	.A2(\localbus/N229 ), 
	.A1(\localbus/N252 ));
   AND2_X1 \localbus/C987  (.ZN(\localbus/N89 ), 
	.A2(\localbus/N218 ), 
	.A1(\localbus/N258 ));
   AND2_X1 \localbus/C988  (.ZN(\localbus/N90 ), 
	.A2(\localbus/N229 ), 
	.A1(\localbus/N258 ));
   AND2_X1 \localbus/C993  (.ZN(\localbus/N95 ), 
	.A2(\localbus/N322 ), 
	.A1(\localbus/N320 ));
   INV_X1 \UUT/Mpath/the_memhandle/I_0  (.ZN(\UUT/Mpath/the_memhandle/N234 ), 
	.A(dmem_isbyte));
   INV_X1 \UUT/Mpath/the_memhandle/I_3  (.ZN(\UUT/Mpath/the_memhandle/N237 ), 
	.A(dmem_ishalf));
   AND2_X1 \UUT/Mpath/the_memhandle/C342  (.ZN(\UUT/Mpath/the_memhandle/N34 ), 
	.A2(\UUT/Mpath/the_memhandle/N236 ), 
	.A1(\UUT/Mpath/the_memhandle/N235 ));
   AND2_X1 \UUT/Mpath/the_memhandle/C344  (.ZN(\UUT/Mpath/the_memhandle/N36 ), 
	.A2(\UUT/Mpath/the_memhandle/N240 ), 
	.A1(\UUT/Mpath/the_memhandle/N239 ));
   INV_X1 \UUT/Mpath/the_memhandle/I_8  (.ZN(\UUT/Mpath/the_memhandle/N37 ), 
	.A(\UUT/Mpath/the_memhandle/N241 ));
   OR2_X1 \UUT/Mpath/the_memhandle/C348  (.ZN(\UUT/Mpath/the_memhandle/N241 ), 
	.A2(\UUT/Mpath/the_memhandle/N240 ), 
	.A1(\UUT/Mpath/mem_baddr [1]));
   OR2_X1 \UUT/Mpath/the_memhandle/C351  (.ZN(\UUT/Mpath/the_memhandle/N242 ), 
	.A2(\UUT/Mpath/mem_baddr [0]), 
	.A1(\UUT/Mpath/the_memhandle/N239 ));
   AND2_X1 \UUT/Mpath/the_memhandle/C353  (.ZN(\UUT/Mpath/the_memhandle/N39 ), 
	.A2(\UUT/Mpath/mem_baddr [0]), 
	.A1(\UUT/Mpath/mem_baddr [1]));
   AND2_X1 \UUT/Mpath/the_memhandle/C354  (.ZN(\UUT/Mpath/the_memhandle/N72 ), 
	.A2(\UUT/Mpath/the_memhandle/N236 ), 
	.A1(\UUT/m_mem_command[SIGN] ));
   INV_X1 \UUT/Mpath/the_memhandle/I_12  (.ZN(\UUT/Mpath/the_memhandle/N76 ), 
	.A(\UUT/Mpath/the_memhandle/N242 ));
   AND2_X1 \UUT/Mpath/the_memhandle/C366  (.ZN(\UUT/Mpath/the_memhandle/N86 ), 
	.A2(\UUT/Mpath/the_memhandle/N238 ), 
	.A1(\UUT/Mpath/the_memhandle/N235 ));
   AND2_X1 \UUT/Mpath/the_memhandle/C369  (.ZN(\UUT/Mpath/the_memhandle/N120 ), 
	.A2(\UUT/Mpath/the_memhandle/N238 ), 
	.A1(\UUT/m_mem_command[SIGN] ));
   OR2_X1 \UUT/Mpath/the_mult/C331  (.ZN(\UUT/Mpath/the_mult/N194 ), 
	.A2(\UUT/Mpath/the_mult/x_mul_command[5] ), 
	.A1(\UUT/Mpath/the_mult/x_mul_command[4] ));
   OR2_X1 \UUT/Mpath/the_mult/C332  (.ZN(\UUT/Mpath/the_mult/N195 ), 
	.A2(\UUT/Mpath/the_mult/N194 ), 
	.A1(\UUT/Mpath/the_mult/N192 ));
   OR2_X1 \UUT/Mpath/the_mult/C333  (.ZN(\UUT/Mpath/the_mult/N196 ), 
	.A2(\UUT/Mpath/the_mult/N195 ), 
	.A1(\UUT/Mpath/the_mult/x_mul_command[2] ));
   OR2_X1 \UUT/Mpath/the_mult/C334  (.ZN(\UUT/Mpath/the_mult/N197 ), 
	.A2(\UUT/Mpath/the_mult/N196 ), 
	.A1(\UUT/Mpath/the_mult/x_mul_command[1] ));
   OR2_X1 \UUT/Mpath/the_mult/C335  (.ZN(\UUT/Mpath/the_mult/N198 ), 
	.A2(\UUT/Mpath/the_mult/N197 ), 
	.A1(\UUT/Mpath/the_mult/N193 ));
   INV_X1 \UUT/Mpath/the_mult/I_8  (.ZN(\UUT/Mpath/the_mult/N220 ), 
	.A(\UUT/d_mul_command [3]));
   INV_X1 \UUT/Mpath/the_mult/I_9  (.ZN(\UUT/Mpath/the_mult/N221 ), 
	.A(\UUT/d_mul_command [2]));
   INV_X1 \UUT/Mpath/the_mult/I_10  (.ZN(\UUT/Mpath/the_mult/N222 ), 
	.A(\UUT/d_mul_command [1]));
   INV_X1 \UUT/Mpath/the_mult/I_11  (.ZN(\UUT/Mpath/the_mult/N223 ), 
	.A(\UUT/d_mul_command [0]));
   OR2_X1 \UUT/Mpath/the_mult/C370  (.ZN(\UUT/Mpath/the_mult/N224 ), 
	.A2(\UUT/d_mul_command [5]), 
	.A1(\UUT/d_mul_command [4]));
   OR2_X1 \UUT/Mpath/the_mult/C371  (.ZN(\UUT/Mpath/the_mult/N225 ), 
	.A2(\UUT/Mpath/the_mult/N224 ), 
	.A1(\UUT/Mpath/the_mult/N220 ));
   OR2_X1 \UUT/Mpath/the_mult/C372  (.ZN(\UUT/Mpath/the_mult/N226 ), 
	.A2(\UUT/Mpath/the_mult/N225 ), 
	.A1(\UUT/Mpath/the_mult/N221 ));
   OR2_X1 \UUT/Mpath/the_mult/C373  (.ZN(\UUT/Mpath/the_mult/N227 ), 
	.A2(\UUT/Mpath/the_mult/N226 ), 
	.A1(\UUT/Mpath/the_mult/N222 ));
   OR2_X1 \UUT/Mpath/the_mult/C404  (.ZN(\UUT/Mpath/the_mult/N251 ), 
	.A2(\UUT/Mpath/the_mult/m_mul_command[5] ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[4] ));
   OR2_X1 \UUT/Mpath/the_mult/C405  (.ZN(\UUT/Mpath/the_mult/N252 ), 
	.A2(\UUT/Mpath/the_mult/N251 ), 
	.A1(\UUT/Mpath/the_mult/N229 ));
   OR2_X1 \UUT/Mpath/the_mult/C406  (.ZN(\UUT/Mpath/the_mult/N253 ), 
	.A2(\UUT/Mpath/the_mult/N252 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[2] ));
   OR2_X1 \UUT/Mpath/the_mult/C407  (.ZN(\UUT/Mpath/the_mult/N254 ), 
	.A2(\UUT/Mpath/the_mult/N253 ), 
	.A1(\UUT/Mpath/the_mult/N230 ));
   OR2_X1 \UUT/Mpath/the_mult/C408  (.ZN(\UUT/Mpath/the_mult/N255 ), 
	.A2(\UUT/Mpath/the_mult/N254 ), 
	.A1(\UUT/Mpath/the_mult/N231 ));
   OR2_X1 \UUT/Mpath/the_mult/C411  (.ZN(\UUT/Mpath/the_mult/N258 ), 
	.A2(\UUT/Mpath/the_mult/N251 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[3] ));
   OR2_X1 \UUT/Mpath/the_mult/C412  (.ZN(\UUT/Mpath/the_mult/N259 ), 
	.A2(\UUT/Mpath/the_mult/N258 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[2] ));
   OR2_X1 \UUT/Mpath/the_mult/C413  (.ZN(\UUT/Mpath/the_mult/N260 ), 
	.A2(\UUT/Mpath/the_mult/N259 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[1] ));
   OR2_X1 \UUT/Mpath/the_mult/C414  (.ZN(\UUT/Mpath/the_mult/N261 ), 
	.A2(\UUT/Mpath/the_mult/N260 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[0] ));
   INV_X1 \UUT/Mpath/the_mult/I_21  (.ZN(\UUT/Mpath/the_mult/N262 ), 
	.A(\UUT/Mpath/the_mult/N261 ));
   OR2_X1 \UUT/Mpath/the_mult/C421  (.ZN(\UUT/Mpath/the_mult/N267 ), 
	.A2(\UUT/Mpath/the_mult/N260 ), 
	.A1(\UUT/Mpath/the_mult/N231 ));
   INV_X1 \UUT/Mpath/the_mult/I_22  (.ZN(\UUT/Mpath/the_mult/N268 ), 
	.A(\UUT/Mpath/the_mult/N267 ));
   OR2_X1 \UUT/Mpath/the_mult/C426  (.ZN(\UUT/Mpath/the_mult/N271 ), 
	.A2(\UUT/Mpath/the_mult/N258 ), 
	.A1(\UUT/Mpath/the_mult/N244 ));
   OR2_X1 \UUT/Mpath/the_mult/C427  (.ZN(\UUT/Mpath/the_mult/N272 ), 
	.A2(\UUT/Mpath/the_mult/N271 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[1] ));
   OR2_X1 \UUT/Mpath/the_mult/C428  (.ZN(\UUT/Mpath/the_mult/N273 ), 
	.A2(\UUT/Mpath/the_mult/N272 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[0] ));
   INV_X1 \UUT/Mpath/the_mult/I_23  (.ZN(\UUT/Mpath/the_mult/N274 ), 
	.A(\UUT/Mpath/the_mult/N273 ));
   OR2_X1 \UUT/Mpath/the_mult/C436  (.ZN(\UUT/Mpath/the_mult/N279 ), 
	.A2(\UUT/Mpath/the_mult/N272 ), 
	.A1(\UUT/Mpath/the_mult/N231 ));
   INV_X1 \UUT/Mpath/the_mult/I_24  (.ZN(\UUT/Mpath/the_mult/N280 ), 
	.A(\UUT/Mpath/the_mult/N279 ));
   OR2_X1 \UUT/Mpath/the_mult/C444  (.ZN(\UUT/Mpath/the_mult/N285 ), 
	.A2(\UUT/Mpath/the_mult/N254 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[0] ));
   OR2_X1 \UUT/Mpath/the_mult/C496  (.ZN(\UUT/Mpath/the_mult/N311 ), 
	.A2(\UUT/Mpath/the_mult/N268 ), 
	.A1(\UUT/Mpath/the_mult/N262 ));
   OR2_X1 \UUT/Mpath/the_mult/C499  (.ZN(\UUT/Mpath/the_mult/N312 ), 
	.A2(\UUT/Mpath/the_mult/N280 ), 
	.A1(\UUT/Mpath/the_mult/N274 ));
   OR2_X1 \UUT/Mpath/the_shift/C151  (.ZN(\UUT/Mpath/the_shift/N106 ), 
	.A2(\UUT/Mpath/the_shift/N104 ), 
	.A1(\UUT/shift_op [1]));
   OR2_X1 \UUT/Mpath/the_shift/C152  (.ZN(\UUT/Mpath/the_shift/N107 ), 
	.A2(\UUT/Mpath/the_shift/N106 ), 
	.A1(\UUT/Mpath/the_shift/N105 ));
   INV_X1 \UUT/Mpath/the_shift/I_2  (.ZN(\UUT/Mpath/the_shift/N108 ), 
	.A(\UUT/Mpath/the_shift/N107 ));
   OR2_X1 \UUT/Mpath/the_shift/C156  (.ZN(\UUT/Mpath/the_shift/N110 ), 
	.A2(\UUT/Mpath/the_shift/N106 ), 
	.A1(\UUT/shift_op [0]));
   INV_X1 \UUT/Mpath/the_shift/I_3  (.ZN(\UUT/Mpath/the_shift/N111 ), 
	.A(\UUT/Mpath/the_shift/N110 ));
   OR2_X1 \UUT/Mpath/the_shift/C159  (.ZN(\UUT/Mpath/the_shift/N113 ), 
	.A2(\UUT/shift_op [2]), 
	.A1(\UUT/Mpath/the_shift/N112 ));
   OR2_X1 \UUT/Mpath/the_shift/C160  (.ZN(\UUT/Mpath/the_shift/N114 ), 
	.A2(\UUT/Mpath/the_shift/N113 ), 
	.A1(\UUT/shift_op [0]));
   INV_X1 \UUT/Mpath/the_shift/I_5  (.ZN(\UUT/Mpath/the_shift/N115 ), 
	.A(\UUT/Mpath/the_shift/N114 ));
   OR2_X1 \UUT/Mpath/the_shift/C163  (.ZN(\UUT/Mpath/the_shift/N116 ), 
	.A2(\UUT/shift_op [2]), 
	.A1(\UUT/shift_op [1]));
   OR2_X1 \UUT/Mpath/the_shift/C164  (.ZN(\UUT/Mpath/the_shift/N117 ), 
	.A2(\UUT/Mpath/the_shift/N116 ), 
	.A1(\UUT/Mpath/the_shift/N105 ));
   INV_X2 \UUT/Mpath/the_shift/I_6  (.ZN(\UUT/Mpath/the_shift/N118 ), 
	.A(\UUT/Mpath/the_shift/N117 ));
   OR2_X1 \UUT/Mpath/the_alu/C476  (.ZN(\UUT/Mpath/the_alu/N469 ), 
	.A2(\UUT/Mpath/the_alu/N466 ), 
	.A1(\UUT/Mpath/the_alu/N453 ));
   OR2_X1 \UUT/Mpath/the_alu/C477  (.ZN(\UUT/Mpath/the_alu/N470 ), 
	.A2(\UUT/Mpath/the_alu/N469 ), 
	.A1(\UUT/Alu_command[OP][3] ));
   OR2_X1 \UUT/Mpath/the_alu/C478  (.ZN(\UUT/Mpath/the_alu/N471 ), 
	.A2(\UUT/Mpath/the_alu/N470 ), 
	.A1(\UUT/Alu_command[OP][2] ));
   OR2_X1 \UUT/Mpath/the_alu/C479  (.ZN(\UUT/Mpath/the_alu/N472 ), 
	.A2(\UUT/Mpath/the_alu/N471 ), 
	.A1(\UUT/Mpath/the_alu/N467 ));
   OR2_X1 \UUT/Mpath/the_alu/C480  (.ZN(\UUT/Mpath/the_alu/N473 ), 
	.A2(\UUT/Mpath/the_alu/N472 ), 
	.A1(\UUT/Mpath/the_alu/N468 ));
   INV_X1 \UUT/Mpath/the_alu/I_9  (.ZN(\UUT/Mpath/the_alu/N474 ), 
	.A(\UUT/Mpath/the_alu/N473 ));
   OR2_X1 \UUT/Mpath/the_alu/C489  (.ZN(\UUT/Mpath/the_alu/N479 ), 
	.A2(\UUT/Mpath/the_alu/N472 ), 
	.A1(\UUT/Alu_command[OP][0] ));
   INV_X1 \UUT/Mpath/the_alu/I_10  (.ZN(\UUT/Mpath/the_alu/N480 ), 
	.A(\UUT/Mpath/the_alu/N479 ));
   OR2_X1 \UUT/Mpath/the_alu/C497  (.ZN(\UUT/Mpath/the_alu/N484 ), 
	.A2(\UUT/Mpath/the_alu/N471 ), 
	.A1(\UUT/Alu_command[OP][1] ));
   OR2_X1 \UUT/Mpath/the_alu/C498  (.ZN(\UUT/Mpath/the_alu/N485 ), 
	.A2(\UUT/Mpath/the_alu/N484 ), 
	.A1(\UUT/Mpath/the_alu/N468 ));
   INV_X1 \UUT/Mpath/the_alu/I_11  (.ZN(\UUT/Mpath/the_alu/N486 ), 
	.A(\UUT/Mpath/the_alu/N485 ));
   OR2_X1 \UUT/Mpath/the_alu/C506  (.ZN(\UUT/Mpath/the_alu/N491 ), 
	.A2(\UUT/Mpath/the_alu/N484 ), 
	.A1(\UUT/Alu_command[OP][0] ));
   OR2_X1 \UUT/Mpath/the_alu/C510  (.ZN(\UUT/Mpath/the_alu/N493 ), 
	.A2(\UUT/Mpath/the_alu/N466 ), 
	.A1(\UUT/Alu_command[OP][4] ));
   OR2_X1 \UUT/Mpath/the_alu/C511  (.ZN(\UUT/Mpath/the_alu/N494 ), 
	.A2(\UUT/Mpath/the_alu/N493 ), 
	.A1(\UUT/Alu_command[OP][3] ));
   OR2_X1 \UUT/Mpath/the_alu/C512  (.ZN(\UUT/Mpath/the_alu/N495 ), 
	.A2(\UUT/Mpath/the_alu/N494 ), 
	.A1(\UUT/Alu_command[OP][2] ));
   OR2_X1 \UUT/Mpath/the_alu/C513  (.ZN(\UUT/Mpath/the_alu/N496 ), 
	.A2(\UUT/Mpath/the_alu/N495 ), 
	.A1(\UUT/Alu_command[OP][1] ));
   OR2_X1 \UUT/Mpath/the_alu/C514  (.ZN(\UUT/Mpath/the_alu/N497 ), 
	.A2(\UUT/Mpath/the_alu/N496 ), 
	.A1(\UUT/Mpath/the_alu/N468 ));
   INV_X1 \UUT/Mpath/the_alu/I_13  (.ZN(\UUT/Mpath/the_alu/N498 ), 
	.A(\UUT/Mpath/the_alu/N497 ));
   OR2_X1 \UUT/Mpath/the_alu/C521  (.ZN(\UUT/Mpath/the_alu/N503 ), 
	.A2(\UUT/Mpath/the_alu/N496 ), 
	.A1(\UUT/Alu_command[OP][0] ));
   OR2_X1 \UUT/Mpath/the_alu/C524  (.ZN(\UUT/Mpath/the_alu/N505 ), 
	.A2(\UUT/Alu_command[OP][5] ), 
	.A1(\UUT/Mpath/the_alu/N453 ));
   OR2_X1 \UUT/Mpath/the_alu/C525  (.ZN(\UUT/Mpath/the_alu/N506 ), 
	.A2(\UUT/Mpath/the_alu/N505 ), 
	.A1(\UUT/Alu_command[OP][3] ));
   OR2_X1 \UUT/Mpath/the_alu/C526  (.ZN(\UUT/Mpath/the_alu/N507 ), 
	.A2(\UUT/Mpath/the_alu/N506 ), 
	.A1(\UUT/Alu_command[OP][2] ));
   OR2_X1 \UUT/Mpath/the_alu/C527  (.ZN(\UUT/Mpath/the_alu/N508 ), 
	.A2(\UUT/Mpath/the_alu/N507 ), 
	.A1(\UUT/Alu_command[OP][1] ));
   OR2_X1 \UUT/Mpath/the_alu/C528  (.ZN(\UUT/Mpath/the_alu/N509 ), 
	.A2(\UUT/Mpath/the_alu/N508 ), 
	.A1(\UUT/Alu_command[OP][0] ));
   OR2_X1 \UUT/Mpath/the_alu/C536  (.ZN(\UUT/Mpath/the_alu/N515 ), 
	.A2(\UUT/Mpath/the_alu/N508 ), 
	.A1(\UUT/Mpath/the_alu/N468 ));
   OR2_X1 \UUT/Mpath/the_alu/C538  (.ZN(\UUT/Mpath/the_alu/N517 ), 
	.A2(\UUT/Alu_command[OP][5] ), 
	.A1(\UUT/Alu_command[OP][4] ));
   OR2_X1 \UUT/Mpath/the_alu/C539  (.ZN(\UUT/Mpath/the_alu/N518 ), 
	.A2(\UUT/Mpath/the_alu/N517 ), 
	.A1(\UUT/Alu_command[OP][3] ));
   OR2_X1 \UUT/Mpath/the_alu/C540  (.ZN(\UUT/Mpath/the_alu/N519 ), 
	.A2(\UUT/Mpath/the_alu/N518 ), 
	.A1(\UUT/Alu_command[OP][2] ));
   OR2_X1 \UUT/Mpath/the_alu/C541  (.ZN(\UUT/Mpath/the_alu/N520 ), 
	.A2(\UUT/Mpath/the_alu/N519 ), 
	.A1(\UUT/Alu_command[OP][1] ));
   AND2_X1 \UUT/Mpath/the_alu/C575  (.ZN(\UUT/Mpath/the_alu/N94 ), 
	.A2(\UUT/Mpath/out_regB[31] ), 
	.A1(\UUT/Mpath/out_regA[31] ));
   OR2_X1 \UUT/Mpath/the_alu/C608  (.ZN(\UUT/Mpath/the_alu/N126 ), 
	.A2(\UUT/Mpath/out_regB[31] ), 
	.A1(\UUT/Mpath/out_regA[31] ));
   XOR2_X1 \UUT/Mpath/the_alu/C641  (.Z(\UUT/Mpath/the_alu/N158 ), 
	.B(\UUT/Mpath/out_regB[31] ), 
	.A(\UUT/Mpath/out_regA[31] ));
   XOR2_X1 \UUT/Mpath/the_alu/C642  (.Z(\UUT/Mpath/the_alu/N159 ), 
	.B(\UUT/Mpath/out_regB[30] ), 
	.A(\UUT/Mpath/out_regA[30] ));
   XOR2_X1 \UUT/Mpath/the_alu/C643  (.Z(\UUT/Mpath/the_alu/N160 ), 
	.B(\UUT/Mpath/out_regB[29] ), 
	.A(\UUT/Mpath/out_regA[29] ));
   XOR2_X1 \UUT/Mpath/the_alu/C644  (.Z(\UUT/Mpath/the_alu/N161 ), 
	.B(\UUT/Mpath/out_regB[28] ), 
	.A(\UUT/Mpath/out_regA[28] ));
   XOR2_X1 \UUT/Mpath/the_alu/C645  (.Z(\UUT/Mpath/the_alu/N162 ), 
	.B(\UUT/Mpath/out_regB[27] ), 
	.A(\UUT/Mpath/out_regA[27] ));
   XOR2_X1 \UUT/Mpath/the_alu/C646  (.Z(\UUT/Mpath/the_alu/N163 ), 
	.B(\UUT/Mpath/out_regB[26] ), 
	.A(\UUT/Mpath/out_regA[26] ));
   XOR2_X1 \UUT/Mpath/the_alu/C647  (.Z(\UUT/Mpath/the_alu/N164 ), 
	.B(\UUT/Mpath/out_regB[25] ), 
	.A(\UUT/Mpath/out_regA[25] ));
   XOR2_X1 \UUT/Mpath/the_alu/C648  (.Z(\UUT/Mpath/the_alu/N165 ), 
	.B(\UUT/Mpath/out_regB[24] ), 
	.A(\UUT/Mpath/out_regA[24] ));
   XOR2_X1 \UUT/Mpath/the_alu/C649  (.Z(\UUT/Mpath/the_alu/N166 ), 
	.B(\UUT/Mpath/out_regB[23] ), 
	.A(\UUT/Mpath/out_regA[23] ));
   XOR2_X1 \UUT/Mpath/the_alu/C650  (.Z(\UUT/Mpath/the_alu/N167 ), 
	.B(\UUT/Mpath/out_regB[22] ), 
	.A(\UUT/Mpath/out_regA[22] ));
   XOR2_X1 \UUT/Mpath/the_alu/C651  (.Z(\UUT/Mpath/the_alu/N168 ), 
	.B(\UUT/Mpath/out_regB[21] ), 
	.A(\UUT/Mpath/out_regA[21] ));
   XOR2_X1 \UUT/Mpath/the_alu/C652  (.Z(\UUT/Mpath/the_alu/N169 ), 
	.B(\UUT/Mpath/out_regB[20] ), 
	.A(\UUT/Mpath/out_regA[20] ));
   XOR2_X1 \UUT/Mpath/the_alu/C653  (.Z(\UUT/Mpath/the_alu/N170 ), 
	.B(\UUT/Mpath/out_regB[19] ), 
	.A(\UUT/Mpath/out_regA[19] ));
   XOR2_X1 \UUT/Mpath/the_alu/C654  (.Z(\UUT/Mpath/the_alu/N171 ), 
	.B(\UUT/Mpath/out_regB[18] ), 
	.A(\UUT/Mpath/out_regA[18] ));
   XOR2_X1 \UUT/Mpath/the_alu/C655  (.Z(\UUT/Mpath/the_alu/N172 ), 
	.B(\UUT/Mpath/out_regB[17] ), 
	.A(\UUT/Mpath/out_regA[17] ));
   XOR2_X1 \UUT/Mpath/the_alu/C656  (.Z(\UUT/Mpath/the_alu/N173 ), 
	.B(\UUT/Mpath/out_regB[16] ), 
	.A(\UUT/Mpath/out_regA[16] ));
   XOR2_X1 \UUT/Mpath/the_alu/C657  (.Z(\UUT/Mpath/the_alu/N174 ), 
	.B(\UUT/Mpath/out_regB[15] ), 
	.A(\UUT/Mpath/out_regA[15] ));
   XOR2_X1 \UUT/Mpath/the_alu/C658  (.Z(\UUT/Mpath/the_alu/N175 ), 
	.B(\UUT/Mpath/out_regB[14] ), 
	.A(\UUT/Mpath/out_regA[14] ));
   XOR2_X1 \UUT/Mpath/the_alu/C659  (.Z(\UUT/Mpath/the_alu/N176 ), 
	.B(\UUT/Mpath/out_regB[13] ), 
	.A(\UUT/Mpath/out_regA[13] ));
   XOR2_X1 \UUT/Mpath/the_alu/C660  (.Z(\UUT/Mpath/the_alu/N177 ), 
	.B(\UUT/Mpath/out_regB[12] ), 
	.A(\UUT/Mpath/out_regA[12] ));
   XOR2_X1 \UUT/Mpath/the_alu/C661  (.Z(\UUT/Mpath/the_alu/N178 ), 
	.B(\UUT/Mpath/out_regB[11] ), 
	.A(\UUT/Mpath/out_regA[11] ));
   XOR2_X1 \UUT/Mpath/the_alu/C662  (.Z(\UUT/Mpath/the_alu/N179 ), 
	.B(\UUT/Mpath/out_regB[10] ), 
	.A(\UUT/Mpath/out_regA[10] ));
   XOR2_X1 \UUT/Mpath/the_alu/C663  (.Z(\UUT/Mpath/the_alu/N180 ), 
	.B(\UUT/Mpath/out_regB[9] ), 
	.A(\UUT/Mpath/out_regA[9] ));
   XOR2_X1 \UUT/Mpath/the_alu/C664  (.Z(\UUT/Mpath/the_alu/N181 ), 
	.B(\UUT/Mpath/out_regB[8] ), 
	.A(\UUT/Mpath/out_regA[8] ));
   XOR2_X1 \UUT/Mpath/the_alu/C665  (.Z(\UUT/Mpath/the_alu/N182 ), 
	.B(\UUT/Mpath/out_regB[7] ), 
	.A(\UUT/Mpath/out_regA[7] ));
   XOR2_X1 \UUT/Mpath/the_alu/C666  (.Z(\UUT/Mpath/the_alu/N183 ), 
	.B(\UUT/Mpath/out_regB[6] ), 
	.A(\UUT/Mpath/out_regA[6] ));
   XOR2_X1 \UUT/Mpath/the_alu/C667  (.Z(\UUT/Mpath/the_alu/N184 ), 
	.B(\UUT/Mpath/out_regB[5] ), 
	.A(\UUT/Mpath/out_regA[5] ));
   XOR2_X1 \UUT/Mpath/the_alu/C668  (.Z(\UUT/Mpath/the_alu/N185 ), 
	.B(\UUT/Mpath/out_regB[4] ), 
	.A(\UUT/Mpath/out_regA[4] ));
   XOR2_X1 \UUT/Mpath/the_alu/C669  (.Z(\UUT/Mpath/the_alu/N186 ), 
	.B(\UUT/Mpath/out_regB[3] ), 
	.A(\UUT/Mpath/out_regA[3] ));
   XOR2_X1 \UUT/Mpath/the_alu/C670  (.Z(\UUT/Mpath/the_alu/N187 ), 
	.B(FE_OFN168_UUT_Mpath_out_regB_2_), 
	.A(FE_OFCN198_UUT_Mpath_out_regA_2_));
   XOR2_X1 \UUT/Mpath/the_alu/C672  (.Z(\UUT/Mpath/the_alu/N189 ), 
	.B(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.A(FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_));
   AND2_X1 \UUT/Mpath/the_alu/C674  (.ZN(\UUT/Mpath/the_alu/N190 ), 
	.A2(\UUT/Mpath/the_alu/N22 ), 
	.A1(\UUT/Mpath/the_alu/N21 ));
   AND2_X1 \UUT/Mpath/the_alu/C675  (.ZN(\UUT/Mpath/the_alu/N191 ), 
	.A2(\UUT/Mpath/the_alu/N24 ), 
	.A1(\UUT/Mpath/the_alu/N23 ));
   AND2_X1 \UUT/Mpath/the_alu/C676  (.ZN(\UUT/Mpath/the_alu/N192 ), 
	.A2(\UUT/Mpath/the_alu/N26 ), 
	.A1(\UUT/Mpath/the_alu/N25 ));
   AND2_X1 \UUT/Mpath/the_alu/C677  (.ZN(\UUT/Mpath/the_alu/N193 ), 
	.A2(\UUT/Mpath/the_alu/N28 ), 
	.A1(\UUT/Mpath/the_alu/N27 ));
   AND2_X1 \UUT/Mpath/the_alu/C678  (.ZN(\UUT/Mpath/the_alu/N194 ), 
	.A2(\UUT/Mpath/the_alu/N30 ), 
	.A1(\UUT/Mpath/the_alu/N29 ));
   AND2_X1 \UUT/Mpath/the_alu/C679  (.ZN(\UUT/Mpath/the_alu/N195 ), 
	.A2(\UUT/Mpath/the_alu/N32 ), 
	.A1(\UUT/Mpath/the_alu/N31 ));
   AND2_X1 \UUT/Mpath/the_alu/C680  (.ZN(\UUT/Mpath/the_alu/N196 ), 
	.A2(\UUT/Mpath/the_alu/N34 ), 
	.A1(\UUT/Mpath/the_alu/N33 ));
   AND2_X1 \UUT/Mpath/the_alu/C681  (.ZN(\UUT/Mpath/the_alu/N197 ), 
	.A2(\UUT/Mpath/the_alu/N36 ), 
	.A1(\UUT/Mpath/the_alu/N35 ));
   AND2_X1 \UUT/Mpath/the_alu/C682  (.ZN(\UUT/Mpath/the_alu/N198 ), 
	.A2(\UUT/Mpath/the_alu/N38 ), 
	.A1(\UUT/Mpath/the_alu/N37 ));
   AND2_X1 \UUT/Mpath/the_alu/C683  (.ZN(\UUT/Mpath/the_alu/N199 ), 
	.A2(\UUT/Mpath/the_alu/N40 ), 
	.A1(\UUT/Mpath/the_alu/N39 ));
   AND2_X1 \UUT/Mpath/the_alu/C684  (.ZN(\UUT/Mpath/the_alu/N200 ), 
	.A2(\UUT/Mpath/the_alu/N42 ), 
	.A1(\UUT/Mpath/the_alu/N41 ));
   AND2_X1 \UUT/Mpath/the_alu/C685  (.ZN(\UUT/Mpath/the_alu/N201 ), 
	.A2(\UUT/Mpath/the_alu/N44 ), 
	.A1(\UUT/Mpath/the_alu/N43 ));
   AND2_X1 \UUT/Mpath/the_alu/C686  (.ZN(\UUT/Mpath/the_alu/N202 ), 
	.A2(\UUT/Mpath/the_alu/N46 ), 
	.A1(\UUT/Mpath/the_alu/N45 ));
   AND2_X1 \UUT/Mpath/the_alu/C687  (.ZN(\UUT/Mpath/the_alu/N203 ), 
	.A2(\UUT/Mpath/the_alu/N48 ), 
	.A1(\UUT/Mpath/the_alu/N47 ));
   AND2_X1 \UUT/Mpath/the_alu/C688  (.ZN(\UUT/Mpath/the_alu/N204 ), 
	.A2(\UUT/Mpath/the_alu/N50 ), 
	.A1(\UUT/Mpath/the_alu/N49 ));
   AND2_X1 \UUT/Mpath/the_alu/C689  (.ZN(\UUT/Mpath/the_alu/N205 ), 
	.A2(\UUT/Mpath/the_alu/N52 ), 
	.A1(\UUT/Mpath/the_alu/N51 ));
   AND2_X1 \UUT/Mpath/the_alu/C690  (.ZN(\UUT/Mpath/the_alu/N206 ), 
	.A2(\UUT/Mpath/the_alu/N54 ), 
	.A1(\UUT/Mpath/the_alu/N53 ));
   AND2_X1 \UUT/Mpath/the_alu/C691  (.ZN(\UUT/Mpath/the_alu/N207 ), 
	.A2(\UUT/Mpath/the_alu/N56 ), 
	.A1(\UUT/Mpath/the_alu/N55 ));
   AND2_X1 \UUT/Mpath/the_alu/C692  (.ZN(\UUT/Mpath/the_alu/N208 ), 
	.A2(\UUT/Mpath/the_alu/N58 ), 
	.A1(\UUT/Mpath/the_alu/N57 ));
   AND2_X1 \UUT/Mpath/the_alu/C693  (.ZN(\UUT/Mpath/the_alu/N209 ), 
	.A2(\UUT/Mpath/the_alu/N60 ), 
	.A1(\UUT/Mpath/the_alu/N59 ));
   AND2_X1 \UUT/Mpath/the_alu/C694  (.ZN(\UUT/Mpath/the_alu/N210 ), 
	.A2(\UUT/Mpath/the_alu/N62 ), 
	.A1(\UUT/Mpath/the_alu/N61 ));
   AND2_X1 \UUT/Mpath/the_alu/C695  (.ZN(\UUT/Mpath/the_alu/N211 ), 
	.A2(\UUT/Mpath/the_alu/N64 ), 
	.A1(\UUT/Mpath/the_alu/N63 ));
   AND2_X1 \UUT/Mpath/the_alu/C696  (.ZN(\UUT/Mpath/the_alu/N212 ), 
	.A2(\UUT/Mpath/the_alu/N66 ), 
	.A1(\UUT/Mpath/the_alu/N65 ));
   AND2_X1 \UUT/Mpath/the_alu/C697  (.ZN(\UUT/Mpath/the_alu/N213 ), 
	.A2(\UUT/Mpath/the_alu/N68 ), 
	.A1(\UUT/Mpath/the_alu/N67 ));
   AND2_X1 \UUT/Mpath/the_alu/C698  (.ZN(\UUT/Mpath/the_alu/N214 ), 
	.A2(\UUT/Mpath/the_alu/N70 ), 
	.A1(\UUT/Mpath/the_alu/N69 ));
   AND2_X1 \UUT/Mpath/the_alu/C699  (.ZN(\UUT/Mpath/the_alu/N215 ), 
	.A2(\UUT/Mpath/the_alu/N72 ), 
	.A1(\UUT/Mpath/the_alu/N71 ));
   AND2_X1 \UUT/Mpath/the_alu/C700  (.ZN(\UUT/Mpath/the_alu/N216 ), 
	.A2(\UUT/Mpath/the_alu/N74 ), 
	.A1(\UUT/Mpath/the_alu/N73 ));
   AND2_X1 \UUT/Mpath/the_alu/C701  (.ZN(\UUT/Mpath/the_alu/N217 ), 
	.A2(\UUT/Mpath/the_alu/N76 ), 
	.A1(\UUT/Mpath/the_alu/N75 ));
   AND2_X1 \UUT/Mpath/the_alu/C702  (.ZN(\UUT/Mpath/the_alu/N218 ), 
	.A2(\UUT/Mpath/the_alu/N78 ), 
	.A1(\UUT/Mpath/the_alu/N77 ));
   AND2_X1 \UUT/Mpath/the_alu/C703  (.ZN(\UUT/Mpath/the_alu/N219 ), 
	.A2(\UUT/Mpath/the_alu/N80 ), 
	.A1(\UUT/Mpath/the_alu/N79 ));
   AND2_X1 \UUT/Mpath/the_alu/C705  (.ZN(\UUT/Mpath/the_alu/N221 ), 
	.A2(\UUT/Mpath/the_alu/N84 ), 
	.A1(\UUT/Mpath/the_alu/N83 ));
   OR2_X1 \UUT/Mpath/C262  (.ZN(\UUT/Mpath/N113 ), 
	.A2(\UUT/Mpath/N111 ), 
	.A1(\UUT/exe_outsel [1]));
   OR2_X1 \UUT/Mpath/C263  (.ZN(\UUT/Mpath/N114 ), 
	.A2(\UUT/Mpath/N113 ), 
	.A1(\UUT/Mpath/N112 ));
   INV_X1 \UUT/Mpath/I_3  (.ZN(\UUT/Mpath/N115 ), 
	.A(\UUT/Mpath/N114 ));
   OR2_X1 \UUT/Mpath/C266  (.ZN(\UUT/Mpath/N117 ), 
	.A2(\UUT/exe_outsel [2]), 
	.A1(\UUT/Mpath/N116 ));
   OR2_X1 \UUT/Mpath/C267  (.ZN(\UUT/Mpath/N118 ), 
	.A2(\UUT/Mpath/N117 ), 
	.A1(\UUT/exe_outsel [0]));
   INV_X2 \UUT/Mpath/I_5  (.ZN(\UUT/Mpath/N119 ), 
	.A(\UUT/Mpath/N118 ));
   OR2_X1 \UUT/Mpath/C275  (.ZN(\UUT/Mpath/N124 ), 
	.A2(\UUT/exe_outsel [2]), 
	.A1(\UUT/exe_outsel [1]));
   OR2_X1 \UUT/Mpath/C276  (.ZN(\UUT/Mpath/N125 ), 
	.A2(\UUT/Mpath/N124 ), 
	.A1(\UUT/Mpath/N112 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_4  (.ZN(\UUT/Mcontrol/st_logic/N55 ), 
	.A(\UUT/byp_controlA[2] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C75  (.ZN(\UUT/Mcontrol/st_logic/N18 ), 
	.A2(\UUT/Mcontrol/st_logic/N55 ), 
	.A1(\UUT/byp_controlA[0] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_5  (.ZN(\UUT/Mcontrol/st_logic/N19 ), 
	.A(\UUT/Mcontrol/st_logic/N18 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_6  (.ZN(\UUT/Mcontrol/st_logic/N52 ), 
	.A(\UUT/byp_controlB[2] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C79  (.ZN(\UUT/Mcontrol/st_logic/N22 ), 
	.A2(\UUT/Mcontrol/st_logic/N52 ), 
	.A1(\UUT/byp_controlB[0] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_7  (.ZN(\UUT/Mcontrol/st_logic/N23 ), 
	.A(\UUT/Mcontrol/st_logic/N22 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_8  (.ZN(\UUT/Mcontrol/st_logic/N24 ), 
	.A(\UUT/m_mem_command[MR] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C85  (.ZN(\UUT/Mcontrol/st_logic/N28 ), 
	.A2(\UUT/Mcontrol/x_mul_command [5]), 
	.A1(\UUT/Mcontrol/x_mul_command [4]));
   OR2_X1 \UUT/Mcontrol/st_logic/C86  (.ZN(\UUT/Mcontrol/st_logic/N29 ), 
	.A2(\UUT/Mcontrol/st_logic/N28 ), 
	.A1(\UUT/Mcontrol/x_mul_command [3]));
   OR2_X1 \UUT/Mcontrol/st_logic/C87  (.ZN(\UUT/Mcontrol/st_logic/N30 ), 
	.A2(\UUT/Mcontrol/st_logic/N29 ), 
	.A1(\UUT/Mcontrol/st_logic/N26 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C88  (.ZN(\UUT/Mcontrol/st_logic/N31 ), 
	.A2(\UUT/Mcontrol/st_logic/N30 ), 
	.A1(\UUT/Mcontrol/st_logic/N27 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C89  (.ZN(\UUT/Mcontrol/st_logic/N32 ), 
	.A2(\UUT/Mcontrol/st_logic/N31 ), 
	.A1(\UUT/Mcontrol/x_mul_command [0]));
   INV_X1 \UUT/Mcontrol/st_logic/I_12  (.ZN(\UUT/Mcontrol/st_logic/N33 ), 
	.A(\UUT/Mcontrol/st_logic/N32 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C98  (.ZN(\UUT/Mcontrol/st_logic/N39 ), 
	.A2(\UUT/Mcontrol/st_logic/N31 ), 
	.A1(\UUT/Mcontrol/st_logic/N34 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_14  (.ZN(\UUT/Mcontrol/st_logic/N40 ), 
	.A(\UUT/Mcontrol/st_logic/N39 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C104  (.ZN(\UUT/Mcontrol/st_logic/N44 ), 
	.A2(\UUT/Mcontrol/st_logic/N52 ), 
	.A1(\UUT/Mcontrol/st_logic/N42 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_17  (.ZN(\UUT/Mcontrol/st_logic/N45 ), 
	.A(\UUT/Mcontrol/st_logic/N44 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C110  (.ZN(\UUT/Mcontrol/st_logic/N49 ), 
	.A2(\UUT/Mcontrol/st_logic/N55 ), 
	.A1(\UUT/Mcontrol/st_logic/N47 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_20  (.ZN(\UUT/Mcontrol/st_logic/N50 ), 
	.A(\UUT/Mcontrol/st_logic/N49 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_24  (.ZN(\UUT/Mcontrol/st_logic/N58 ), 
	.A(\UUT/Mcontrol/d_jump_type[2] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C126  (.ZN(\UUT/Mcontrol/st_logic/N61 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N262 ), 
	.A1(\UUT/Mcontrol/st_logic/N58 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C128  (.ZN(\UUT/Mcontrol/st_logic/N63 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N264 ), 
	.A1(\UUT/Mcontrol/d_jump_type[0] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_26  (.ZN(\UUT/Mcontrol/st_logic/N65 ), 
	.A(\UUT/Mcontrol/d_jump_type[0] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C136  (.ZN(\UUT/Mcontrol/st_logic/N70 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N264 ), 
	.A1(\UUT/Mcontrol/st_logic/N65 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_27  (.ZN(\UUT/Mcontrol/st_logic/N71 ), 
	.A(\UUT/Mcontrol/st_logic/N70 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C155  (.ZN(\UUT/Mcontrol/st_logic/N86 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N262 ), 
	.A1(\UUT/Mcontrol/d_jump_type[2] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C157  (.ZN(\UUT/Mcontrol/st_logic/N88 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N252 ), 
	.A1(\UUT/Mcontrol/d_jump_type[0] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_30  (.ZN(\UUT/Mcontrol/st_logic/N89 ), 
	.A(\UUT/Mcontrol/st_logic/N88 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C164  (.ZN(\UUT/Mcontrol/st_logic/N94 ), 
	.A2(\UUT/Mcontrol/st_logic/N86 ), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N224 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C165  (.ZN(\UUT/Mcontrol/st_logic/N95 ), 
	.A2(\UUT/Mcontrol/st_logic/N94 ), 
	.A1(\UUT/Mcontrol/st_logic/N65 ));
   INV_X1 \UUT/Mcontrol/st_logic/I_32  (.ZN(\UUT/Mcontrol/st_logic/N96 ), 
	.A(\UUT/Mcontrol/st_logic/N95 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C172  (.ZN(\UUT/Mcontrol/st_logic/N100 ), 
	.A2(\UUT/Mcontrol/st_logic/N61 ), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N224 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C173  (.ZN(\UUT/Mcontrol/st_logic/N101 ), 
	.A2(\UUT/Mcontrol/st_logic/N100 ), 
	.A1(\UUT/Mcontrol/d_jump_type[0] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_33  (.ZN(\UUT/Mcontrol/st_logic/N102 ), 
	.A(\UUT/Mcontrol/st_logic/N101 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C179  (.ZN(\UUT/Mcontrol/st_logic/N106 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N114 ), 
	.A1(\UUT/Mcontrol/d_jump_type[2] ));
   INV_X1 \UUT/Mcontrol/st_logic/I_35  (.ZN(\UUT/Mcontrol/st_logic/N109 ), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N125 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C193  (.ZN(\UUT/Mcontrol/st_logic/N2 ), 
	.A2(\UUT/Mcontrol/st_logic/N110 ), 
	.A1(\localbus/c1_op[OP][0] ));
   OR2_X1 \UUT/Mcontrol/st_logic/C194  (.ZN(\UUT/Mcontrol/st_logic/N110 ), 
	.A2(\UUT/Mcontrol/st_logic/N23 ), 
	.A1(\UUT/Mcontrol/st_logic/N19 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C195  (.ZN(\UUT/Mcontrol/st_logic/N3 ), 
	.A2(\UUT/Mcontrol/st_logic/N109 ), 
	.A1(\UUT/Mcontrol/st_logic/N114 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C196  (.ZN(\UUT/Mcontrol/st_logic/N114 ), 
	.A2(\UUT/Mcontrol/st_logic/N102 ), 
	.A1(\UUT/Mcontrol/st_logic/N113 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C197  (.ZN(\UUT/Mcontrol/st_logic/N113 ), 
	.A2(\UUT/Mcontrol/st_logic/N96 ), 
	.A1(\UUT/Mcontrol/st_logic/N112 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C198  (.ZN(\UUT/Mcontrol/st_logic/N112 ), 
	.A2(\UUT/Mcontrol/st_logic/N89 ), 
	.A1(\UUT/Mcontrol/st_logic/N111 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C199  (.ZN(\UUT/Mcontrol/st_logic/N111 ), 
	.A2(\UUT/Mcontrol/st_logic/N71 ), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N266 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C201  (.ZN(\UUT/Mcontrol/st_logic/N5 ), 
	.A2(\UUT/Mcontrol/st_logic/N116 ), 
	.A1(\UUT/Mcontrol/st_logic/N115 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C202  (.ZN(\UUT/Mcontrol/st_logic/N115 ), 
	.A2(\UUT/Mcontrol/st_logic/N111 ), 
	.A1(\UUT/Mcontrol/st_logic/N45 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C203  (.ZN(\UUT/Mcontrol/st_logic/N116 ), 
	.A2(\UUT/Mcontrol/st_logic/N3 ), 
	.A1(\UUT/Mcontrol/st_logic/N50 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C204  (.ZN(\UUT/Mcontrol/st_logic/N6 ), 
	.A2(\UUT/Mcontrol/st_logic/N5 ), 
	.A1(\UUT/Mcontrol/st_logic/N24 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C205  (.ZN(\UUT/Mcontrol/st_logic/N7 ), 
	.A2(\UUT/Mcontrol/st_logic/N118 ), 
	.A1(\UUT/Mcontrol/st_logic/N117 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C206  (.ZN(\UUT/Mcontrol/st_logic/N117 ), 
	.A2(\UUT/Mcontrol/st_logic/N111 ), 
	.A1(\UUT/Mcontrol/st_logic/N23 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C207  (.ZN(\UUT/Mcontrol/st_logic/N118 ), 
	.A2(\UUT/Mcontrol/st_logic/N3 ), 
	.A1(\UUT/Mcontrol/st_logic/N19 ));
   AND2_X1 \UUT/Mcontrol/st_logic/C208  (.ZN(\UUT/Mcontrol/st_logic/N8 ), 
	.A2(\UUT/Mcontrol/st_logic/N7 ), 
	.A1(\UUT/Mcontrol/st_logic/N119 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C209  (.ZN(\UUT/Mcontrol/st_logic/N119 ), 
	.A2(\UUT/Mcontrol/st_logic/N40 ), 
	.A1(\UUT/Mcontrol/st_logic/N33 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C211  (.ZN(\UUT/Mcontrol/st_logic/N10 ), 
	.A2(\UUT/Mcontrol/st_logic/N8 ), 
	.A1(\UUT/Mcontrol/st_logic/N120 ));
   OR2_X1 \UUT/Mcontrol/st_logic/C212  (.ZN(\UUT/Mcontrol/st_logic/N120 ), 
	.A2(\UUT/Mcontrol/st_logic/N6 ), 
	.A1(\UUT/Mcontrol/st_logic/N2 ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C19  (.ZN(\UUT/Mcontrol/bp_logicB/N5 ), 
	.A2(\UUT/Mcontrol/x_rd[4] ), 
	.A1(\UUT/Mcontrol/x_rd[3] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C20  (.ZN(\UUT/Mcontrol/bp_logicB/N6 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N5 ), 
	.A1(\UUT/Mcontrol/x_rd[2] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C21  (.ZN(\UUT/Mcontrol/bp_logicB/N7 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N6 ), 
	.A1(\UUT/Mcontrol/x_rd[1] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C22  (.ZN(\UUT/Mcontrol/bp_logicB/N8 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N7 ), 
	.A1(\UUT/Mcontrol/x_rd[0] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C26  (.ZN(\UUT/Mcontrol/bp_logicB/N10 ), 
	.A2(\UUT/Mcontrol/m_sampled_xrd[4] ), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[3] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C27  (.ZN(\UUT/Mcontrol/bp_logicB/N11 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N10 ), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[2] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C28  (.ZN(\UUT/Mcontrol/bp_logicB/N12 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N11 ), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[1] ));
   OR2_X1 \UUT/Mcontrol/bp_logicB/C29  (.ZN(\UUT/Mcontrol/bp_logicB/N13 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N12 ), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[0] ));
   INV_X1 \UUT/Mcontrol/bp_logicB/I_3  (.ZN(\UUT/Mcontrol/bp_logicB/N14 ), 
	.A(\UUT/m_we ));
   AND2_X1 \UUT/Mcontrol/bp_logicB/C36  (.ZN(\UUT/Mcontrol/bp_logicB/exec_main ), 
	.A2(\UUT/Mcontrol/bp_logicB/N9 ), 
	.A1(\UUT/Mcontrol/bp_logicB/N15 ));
   AND2_X1 \UUT/Mcontrol/bp_logicB/C37  (.ZN(\UUT/Mcontrol/bp_logicB/N15 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N8 ), 
	.A1(\UUT/Mcontrol/bp_logicB/N2 ));
   AND2_X1 \UUT/Mcontrol/bp_logicB/C38  (.ZN(\UUT/Mcontrol/bp_logicB/memory_main ), 
	.A2(\UUT/Mcontrol/bp_logicB/N14 ), 
	.A1(\UUT/Mcontrol/bp_logicB/N16 ));
   AND2_X1 \UUT/Mcontrol/bp_logicB/C39  (.ZN(\UUT/Mcontrol/bp_logicB/N16 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N13 ), 
	.A1(\UUT/Mcontrol/bp_logicB/N3 ));
   INV_X1 \UUT/Mcontrol/bp_logicA/I_1  (.ZN(\UUT/Mcontrol/bp_logicA/N9 ), 
	.A(\UUT/x_we ));
   AND2_X1 \UUT/Mcontrol/bp_logicA/C36  (.ZN(\UUT/Mcontrol/bp_logicA/exec_main ), 
	.A2(\UUT/Mcontrol/bp_logicA/N9 ), 
	.A1(\UUT/Mcontrol/bp_logicA/N15 ));
   AND2_X1 \UUT/Mcontrol/bp_logicA/C37  (.ZN(\UUT/Mcontrol/bp_logicA/N15 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N8 ), 
	.A1(\UUT/Mcontrol/bp_logicA/N2 ));
   AND2_X1 \UUT/Mcontrol/bp_logicA/C38  (.ZN(\UUT/Mcontrol/bp_logicA/memory_main ), 
	.A2(\UUT/Mcontrol/bp_logicB/N14 ), 
	.A1(\UUT/Mcontrol/bp_logicA/N16 ));
   AND2_X1 \UUT/Mcontrol/bp_logicA/C39  (.ZN(\UUT/Mcontrol/bp_logicA/N16 ), 
	.A2(\UUT/Mcontrol/bp_logicB/N13 ), 
	.A1(\UUT/Mcontrol/bp_logicA/N3 ));
   INV_X1 \UUT/Mcontrol/Nextpc_decoding/I_0  (.ZN(\UUT/Mcontrol/st_logic/N103 ), 
	.A(\UUT/Mcontrol/d_jump_type[3] ));
   OR2_X1 \UUT/Mcontrol/Nextpc_decoding/C335  (.ZN(\UUT/Mcontrol/Nextpc_decoding/N241 ), 
	.A2(\UUT/Mcontrol/st_logic/N94 ), 
	.A1(\UUT/Mcontrol/d_jump_type[0] ));
   INV_X1 \UUT/Mcontrol/Nextpc_decoding/I_14  (.ZN(\UUT/Mcontrol/Nextpc_decoding/N242 ), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N241 ));
   OR2_X1 \UUT/Mcontrol/Nextpc_decoding/C342  (.ZN(\UUT/Mcontrol/Nextpc_decoding/N247 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N252 ), 
	.A1(\UUT/Mcontrol/st_logic/N65 ));
   INV_X1 \UUT/Mcontrol/Nextpc_decoding/I_18  (.ZN(\UUT/Mcontrol/Nextpc_decoding/N266 ), 
	.A(\UUT/Mcontrol/st_logic/N63 ));
   AND2_X2 \UUT/Mcontrol/Nextpc_decoding/C397  (.ZN(\UUT/Mcontrol/Nextpc_decoding/N32 ), 
	.A2(n6860), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N222 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_0  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1875 ), 
	.A(\UUT/Mcontrol/d_instr [31]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_1  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1876 ), 
	.A(\UUT/Mcontrol/d_instr [30]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_2  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1877 ), 
	.A(\UUT/Mcontrol/d_sampled_finstr [29]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2052  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1879 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1889 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1877 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2053  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1880 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1879 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2054  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1881 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1880 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2055  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1882 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1881 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2058  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1883 ), 
	.A2(\UUT/Mcontrol/d_instr [5]), 
	.A1(\UUT/Mcontrol/d_instr [4]));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2059  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1884 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1883 ), 
	.A1(\UUT/Mcontrol/d_instr [3]));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2060  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1885 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1884 ), 
	.A1(\UUT/Mcontrol/d_instr [2]));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2061  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1886 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1885 ), 
	.A1(\UUT/Mcontrol/d_instr [1]));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2062  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1887 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1886 ), 
	.A1(\UUT/Mcontrol/d_instr [0]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_4  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1888 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1887 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_7  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1900 ), 
	.A(\UUT/Mcontrol/d_instr [4]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_8  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1901 ), 
	.A(\UUT/Mcontrol/d_instr [0]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2082  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1902 ), 
	.A2(\UUT/Mcontrol/d_instr [5]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1900 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2083  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1903 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1902 ), 
	.A1(\UUT/Mcontrol/d_instr [3]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2084  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1904 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1903 ), 
	.A1(\UUT/Mcontrol/d_instr [2]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2085  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1905 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1904 ), 
	.A1(\UUT/Mcontrol/d_instr [1]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2086  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1906 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1905 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1901 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_9  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1907 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1906 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2088  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1908 ), 
	.A2(\UUT/Mcontrol/d_instr [5]), 
	.A1(\UUT/Mcontrol/d_instr [4]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2089  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1909 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1908 ), 
	.A1(\UUT/Mcontrol/d_instr [3]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2090  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1910 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1909 ), 
	.A1(\UUT/Mcontrol/d_instr [2]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2091  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1911 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1910 ), 
	.A1(\UUT/Mcontrol/d_instr [1]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2092  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1912 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1911 ), 
	.A1(\UUT/Mcontrol/d_instr [0]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_10  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1913 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1912 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2094  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1914 ), 
	.A2(\UUT/Mcontrol/d_instr [7]), 
	.A1(\UUT/Mcontrol/d_instr [6]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_11  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1915 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1914 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_13  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1921 ), 
	.A(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2109  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1924 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1923 ), 
	.A1(\UUT/Mcontrol/d_instr [29]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2110  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1925 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1924 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2111  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1926 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1925 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2112  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1927 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1926 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_15  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1928 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1927 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2120  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1933 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1926 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_16  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1934 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1933 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2127  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1938 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1925 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2128  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1939 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1938 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_17  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1940 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1939 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2142  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1948 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1923 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1877 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2143  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1949 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1948 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2144  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1950 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1949 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2145  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1951 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1950 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_19  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1952 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1951 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2154  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1957 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1950 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_20  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1958 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1957 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2162  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1962 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1949 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2163  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1963 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1962 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2171  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1969 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1962 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2177  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1972 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2020 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1877 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2178  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1973 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1972 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2179  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1974 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1973 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2180  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1974 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2188  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1980 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1973 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2189  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1980 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2197  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1987 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1980 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   INV_X1 \UUT/Mcontrol/Operation_decoding32/I_26  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1989 ), 
	.A(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2204  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1991 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2020 ), 
	.A1(\UUT/Mcontrol/d_instr [29]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2205  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1992 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1991 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1989 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2206  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1993 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1992 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2207  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1994 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1993 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2224  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2005 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1992 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2249  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2022 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1991 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2250  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2023 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2022 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2258  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2029 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2022 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2259  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2030 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2029 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2270  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2039 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2086 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1877 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2271  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2040 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2039 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2272  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2041 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2040 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2279  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2045 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2086 ), 
	.A1(\UUT/Mcontrol/d_instr [29]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2280  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2046 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2045 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1989 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2281  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2047 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2046 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2290  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2047 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2297  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2059 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2046 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2298  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2060 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2059 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2305  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2066 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2059 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2311  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2070 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2045 ), 
	.A1(\UUT/Mcontrol/d_instr [28]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2312  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2071 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2070 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1921 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2326  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2083 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2070 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2327  (.ZN(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2083 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   AND2_X1 \UUT/Mcontrol/Operation_decoding32/C2606  (.ZN(\UUT/Mcontrol/Operation_decoding32/N62 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1915 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1913 ));
   OR2_X1 \UUT/Mcontrol/Operation_decoding32/C2608  (.ZN(\UUT/Mcontrol/Operation_decoding32/N1871 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1888 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1882 ));
   AND2_X1 \UUT/Mcontrol/C112  (.ZN(I_BUSY), 
	.A2(net54843), 
	.A1(n978));
   OR2_X1 \UUT/regfile/C1388  (.ZN(\UUT/regfile/N260 ), 
	.A2(\UUT/rs1_addr [4]), 
	.A1(FE_OFCN199_UUT_rs1_addr_3_));
   OR2_X1 \UUT/regfile/C1389  (.ZN(\UUT/regfile/N261 ), 
	.A2(\UUT/regfile/N260 ), 
	.A1(\UUT/rs1_addr [2]));
   OR2_X1 \UUT/regfile/C1390  (.ZN(\UUT/regfile/N262 ), 
	.A2(\UUT/regfile/N261 ), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   OR2_X1 \UUT/regfile/C1394  (.ZN(\UUT/regfile/N265 ), 
	.A2(\UUT/rs2_addr [4]), 
	.A1(\UUT/rs2_addr [3]));
   OR2_X1 \UUT/regfile/C1395  (.ZN(\UUT/regfile/N266 ), 
	.A2(\UUT/regfile/N265 ), 
	.A1(\UUT/rs2_addr [2]));
   OR2_X1 \UUT/regfile/C1396  (.ZN(\UUT/regfile/N267 ), 
	.A2(\UUT/regfile/N266 ), 
	.A1(\UUT/rs2_addr [1]));
   OR2_X1 \UUT/regfile/C1401  (.ZN(\UUT/regfile/N272 ), 
	.A2(\UUT/regfile/N358 ), 
	.A1(\UUT/rd_addr [3]));
   OR2_X1 \UUT/regfile/C1402  (.ZN(\UUT/regfile/N273 ), 
	.A2(\UUT/regfile/N272 ), 
	.A1(\UUT/rd_addr [2]));
   INV_X1 \UUT/regfile/I_7  (.ZN(\UUT/regfile/N290 ), 
	.A(\UUT/rd_addr [2]));
   OR2_X1 \UUT/regfile/C1424  (.ZN(\UUT/regfile/N293 ), 
	.A2(\UUT/regfile/N272 ), 
	.A1(\UUT/regfile/N290 ));
   INV_X1 \UUT/regfile/I_12  (.ZN(\UUT/regfile/N315 ), 
	.A(\UUT/rd_addr [3]));
   OR2_X1 \UUT/regfile/C1455  (.ZN(\UUT/regfile/N317 ), 
	.A2(\UUT/regfile/N358 ), 
	.A1(\UUT/regfile/N315 ));
   OR2_X1 \UUT/regfile/C1456  (.ZN(\UUT/regfile/N318 ), 
	.A2(\UUT/regfile/N317 ), 
	.A1(\UUT/rd_addr [2]));
   OR2_X1 \UUT/regfile/C1489  (.ZN(\UUT/regfile/N342 ), 
	.A2(\UUT/regfile/N317 ), 
	.A1(\UUT/regfile/N290 ));
   INV_X1 \UUT/regfile/I_21  (.ZN(\UUT/regfile/N455 ), 
	.A(\UUT/regfile/N358 ));
   OR2_X1 \UUT/regfile/C1523  (.ZN(\UUT/regfile/N366 ), 
	.A2(\UUT/regfile/N455 ), 
	.A1(\UUT/rd_addr [3]));
   OR2_X1 \UUT/regfile/C1524  (.ZN(\UUT/regfile/N367 ), 
	.A2(\UUT/regfile/N366 ), 
	.A1(\UUT/rd_addr [2]));
   OR2_X1 \UUT/regfile/C1557  (.ZN(\UUT/regfile/N391 ), 
	.A2(\UUT/regfile/N366 ), 
	.A1(\UUT/regfile/N290 ));
   OR2_X1 \UUT/regfile/C1592  (.ZN(\UUT/regfile/N414 ), 
	.A2(\UUT/regfile/N455 ), 
	.A1(\UUT/regfile/N315 ));
   OR2_X1 \UUT/regfile/C1593  (.ZN(\UUT/regfile/N415 ), 
	.A2(\UUT/regfile/N414 ), 
	.A1(\UUT/rd_addr [2]));
   OR2_X1 \UUT/regfile/C1630  (.ZN(\UUT/regfile/N439 ), 
	.A2(\UUT/regfile/N414 ), 
	.A1(\UUT/regfile/N290 ));
   OR2_X1 \UUT/C150  (.ZN(\UUT/N3 ), 
	.A2(\localbus/N46 ), 
	.A1(\localbus/c1_op[OP][0] ));
   AND2_X1 C271 (.ZN(N178), 
	.A2(\UUT/Mpath/the_memhandle/N234 ), 
	.A1(dmem_ishalf));
   AND2_X1 C270 (.ZN(N42), 
	.A2(N172), 
	.A1(N178));
   AND2_X1 C267 (.ZN(N43), 
	.A2(N171), 
	.A1(N178));
   AND2_X1 C264 (.ZN(N35), 
	.A2(N168), 
	.A1(N178));
   AND2_X1 C261 (.ZN(N31), 
	.A2(N165), 
	.A1(N178));
   AND2_X1 C259 (.ZN(N174), 
	.A2(dmem_isbyte), 
	.A1(\UUT/Mpath/the_memhandle/N237 ));
   AND2_X1 C258 (.ZN(N27), 
	.A2(D_ADDR_OUTBUS[1]), 
	.A1(N174));
   AND2_X1 C255 (.ZN(N22), 
	.A2(N169), 
	.A1(N174));
   INV_X1 I_19 (.ZN(iram_rd), 
	.A(I_BUSY));
   AND2_X1 C246 (.ZN(N172), 
	.A2(D_ADDR_OUTBUS[1]), 
	.A1(D_ADDR_OUTBUS[0]));
   INV_X1 I_18 (.ZN(N171), 
	.A(N170));
   OR2_X1 C244 (.ZN(N170), 
	.A2(N169), 
	.A1(D_ADDR_OUTBUS[0]));
   INV_X1 I_17 (.ZN(N169), 
	.A(D_ADDR_OUTBUS[1]));
   INV_X1 I_16 (.ZN(N168), 
	.A(N167));
   OR2_X1 C241 (.ZN(N167), 
	.A2(D_ADDR_OUTBUS[1]), 
	.A1(N166));
   INV_X1 I_15 (.ZN(N166), 
	.A(D_ADDR_OUTBUS[0]));
   INV_X1 I_14 (.ZN(N165), 
	.A(N164));
   OR2_X1 C238 (.ZN(N164), 
	.A2(D_ADDR_OUTBUS[1]), 
	.A1(D_ADDR_OUTBUS[0]));
   DFFS_X1 \localbus/c2_op_reg[MASTER]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\localbus/c2_op[MASTER] ), 
	.D(\localbus/c1_op[MASTER] ), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N84 ), 
	.Q(\UUT/Mpath/out_regB[0] ), 
	.D(n4335), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [31]), 
	.D(n4334), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/N111 ), 
	.Q(\UUT/exe_outsel [2]), 
	.D(n4333), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[0] ), 
	.D(n4332), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5677), 
	.D(n4331), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5709), 
	.Q(\UUT/Mpath/the_mult/acc_out[32] ), 
	.D(n4330), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5455), 
	.D(n4328), 
	.CK(CLK));
   DFFR_X1 \localbus/c2_op_reg[SLAVE][1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\localbus/c2_op[SLAVE][1] ), 
	.D(1'b0), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N64 ), 
	.Q(\UUT/Mpath/out_regB[10] ), 
	.D(n4325), 
	.CK(CLK));
   DFFR_X1 \localbus/c2_op_reg[SLAVE][0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\localbus/N219 ), 
	.Q(\localbus/c2_op[SLAVE][0] ), 
	.D(\localbus/c1_op[SLAVE][0] ), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N68 ), 
	.Q(\UUT/Mpath/out_regB[8] ), 
	.D(n4324), 
	.CK(CLK));
   DFFS_X1 \localbus/c2_op_reg[SLAVE][2]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\localbus/c2_op[SLAVE][2] ), 
	.D(\localbus/N227 ), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_memhandle/N240 ), 
	.Q(\UUT/Mpath/mem_baddr [0]), 
	.D(n4322), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5527), 
	.D(n4321), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[63]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[63] ), 
	.D(n4320), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[62]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[62] ), 
	.D(n4319), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[61]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[61] ), 
	.D(n4318), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[60]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[60] ), 
	.D(n4317), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[59]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[59] ), 
	.D(n4316), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[58]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[58] ), 
	.D(n4315), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[57]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[57] ), 
	.D(n4314), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[56]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[56] ), 
	.D(n4313), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[55]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[55] ), 
	.D(n4312), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[54]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[54] ), 
	.D(n4311), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[53]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[53] ), 
	.D(n4310), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[52]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[52] ), 
	.D(n4309), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[51]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[51] ), 
	.D(n4308), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[49]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[49] ), 
	.D(n4306), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[48]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[48] ), 
	.D(n4305), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[47]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[47] ), 
	.D(n4304), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[46]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[46] ), 
	.D(n4303), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[45]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[45] ), 
	.D(n4302), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[44]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[44] ), 
	.D(n4301), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[43]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[43] ), 
	.D(n4300), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[42]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[42] ), 
	.D(n4299), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[41]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[41] ), 
	.D(n4298), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[40]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[40] ), 
	.D(n4297), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[39]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[39] ), 
	.D(n4296), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[38]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[38] ), 
	.D(n4295), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[37]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[37] ), 
	.D(n4294), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[36]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[36] ), 
	.D(n4293), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[35]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[35] ), 
	.D(n4292), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[34]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[34] ), 
	.D(n4291), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[33]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[33] ), 
	.D(n4290), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[32]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[32] ), 
	.D(n4289), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[31] ), 
	.D(n4288), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[30] ), 
	.D(n4287), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[29] ), 
	.D(n4286), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[28] ), 
	.D(n4285), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[27] ), 
	.D(n4284), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[26] ), 
	.D(n4283), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[25] ), 
	.D(n4282), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[24] ), 
	.D(n4281), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[23] ), 
	.D(n4280), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[22] ), 
	.D(n4279), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[21] ), 
	.D(n4278), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[20] ), 
	.D(n4277), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[19] ), 
	.D(n4276), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[18] ), 
	.D(n4275), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[17] ), 
	.D(n4274), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[16] ), 
	.D(n4273), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[15] ), 
	.D(n4272), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[14] ), 
	.D(n4271), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[13] ), 
	.D(n4270), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[12] ), 
	.D(n4269), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[11] ), 
	.D(n4268), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[10] ), 
	.D(n4267), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[9] ), 
	.D(n4266), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[8] ), 
	.D(n4265), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[7] ), 
	.D(n4264), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[6] ), 
	.D(n4263), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[5] ), 
	.D(n4262), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[4] ), 
	.D(n4261), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[3] ), 
	.D(n4260), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[2] ), 
	.D(n4259), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[1] ), 
	.D(n4258), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[0] ), 
	.D(n4257), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[0]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mcontrol/st_logic/N34 ), 
	.Q(\UUT/Mcontrol/x_mul_command [0]), 
	.D(n4255), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [30]), 
	.D(n4254), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [29]), 
	.D(n4253), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2785), 
	.Q(\UUT/Mcontrol/d_instr [28]), 
	.D(n4252), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2784), 
	.Q(\UUT/Mcontrol/d_instr [27]), 
	.D(n4251), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2783), 
	.Q(\UUT/Mcontrol/d_instr [26]), 
	.D(n4250), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[SIGN]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), 
	.D(n4249), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MW]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2781), 
	.Q(\UUT/Mcontrol/x_sampled_dmem_command[MW] ), 
	.D(n4248), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MR]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_sampled_dmem_command[MR] ), 
	.D(n4247), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MH]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_sampled_dmem_command[MH] ), 
	.D(n4246), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mem_command_reg[MB]  (.SN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_sampled_dmem_command[MB] ), 
	.D(n4245), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [25]), 
	.D(n4244), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [24]), 
	.D(n4243), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [23]), 
	.D(n4242), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [22]), 
	.D(n4241), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [21]), 
	.D(n4240), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [20]), 
	.D(n4239), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [19]), 
	.D(n4238), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [18]), 
	.D(n4237), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [17]), 
	.D(n4236), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [16]), 
	.D(n4235), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [15]), 
	.D(n4234), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [14]), 
	.D(n4233), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [13]), 
	.D(n4232), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [12]), 
	.D(n4231), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [11]), 
	.D(n4230), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [10]), 
	.D(n4229), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [9]), 
	.D(n4228), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [8]), 
	.D(n4227), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [7]), 
	.D(n4226), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [6]), 
	.D(n4225), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [5]), 
	.D(n4224), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2756), 
	.Q(\UUT/Mcontrol/x_mul_command [5]), 
	.D(n4223), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[5] ), 
	.D(n4222), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2754), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[5] ), 
	.D(n4221), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [4]), 
	.D(n4220), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2752), 
	.Q(\UUT/Mcontrol/x_mul_command [4]), 
	.D(n4219), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[4] ), 
	.D(n4218), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2750), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[4] ), 
	.D(n4217), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [3]), 
	.D(n4216), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[3]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2748), 
	.Q(\UUT/Mcontrol/x_mul_command [3]), 
	.D(n4215), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N192 ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[3] ), 
	.D(n4214), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N229 ), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[3] ), 
	.D(n4213), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [2]), 
	.D(n4212), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[2]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mcontrol/st_logic/N26 ), 
	.D(n4211), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[2] ), 
	.D(n4210), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N244 ), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[2] ), 
	.D(n4209), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [1]), 
	.D(n4208), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_mul_command_reg[1]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mcontrol/st_logic/N27 ), 
	.D(n4207), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[1] ), 
	.D(n4206), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N230 ), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[1] ), 
	.D(n4205), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_fd/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/d_sampled_finstr [0]), 
	.D(n4204), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multop/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N193 ), 
	.Q(\UUT/Mpath/the_mult/x_mul_command[0] ), 
	.D(n4203), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_command_reg/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_mult/N231 ), 
	.Q(\UUT/Mpath/the_mult/m_mul_command[0] ), 
	.D(n4202), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_rd[4] ), 
	.D(n4201), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2741), 
	.Q(\UUT/Mcontrol/m_sampled_xrd[4] ), 
	.D(n4200), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_rd[3] ), 
	.D(n4199), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2739), 
	.Q(\UUT/Mcontrol/m_sampled_xrd[3] ), 
	.D(n4198), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_rd[2] ), 
	.D(n4197), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2737), 
	.Q(\UUT/Mcontrol/m_sampled_xrd[2] ), 
	.D(n4196), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_rd[1] ), 
	.D(n4195), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2735), 
	.Q(\UUT/Mcontrol/m_sampled_xrd[1] ), 
	.D(n4194), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_rd1_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/x_rd[0] ), 
	.D(n4193), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_xm/out_rd1_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mcontrol/m_sampled_xrd[0] ), 
	.D(n4192), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[10]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2732), 
	.Q(\UUT/Mcontrol/f_currpc [10]), 
	.D(n4191), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_dx/out_rf_we_reg  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mcontrol/bp_logicB/N9 ), 
	.Q(\UUT/x_we ), 
	.D(n4190), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_xm/out_rf_we_reg  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n5413), 
	.Q(\UUT/m_we ), 
	.D(n4189), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5676), 
	.Q(\UUT/Mpath/the_mult/acc_out[0] ), 
	.D(n4188), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5092), 
	.D(n4187), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5091), 
	.D(n4186), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5068), 
	.D(n4185), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5062), 
	.D(n4184), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4644), 
	.D(n4183), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4643), 
	.D(n4182), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4620), 
	.D(n4181), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4614), 
	.D(n4180), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4580), 
	.Q(\UUT/regfile/reg_out[5][0] ), 
	.D(n4179), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4579), 
	.Q(\UUT/regfile/reg_out[5][10] ), 
	.D(n4178), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4556), 
	.Q(\UUT/regfile/reg_out[5][31] ), 
	.D(n4177), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4550), 
	.Q(\UUT/regfile/reg_out[5][8] ), 
	.D(n4176), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4516), 
	.D(n4175), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4515), 
	.D(n4174), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4492), 
	.D(n4173), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4486), 
	.D(n4172), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4452), 
	.D(n4171), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4451), 
	.D(n4170), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4428), 
	.D(n4169), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4422), 
	.D(n4168), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5380), 
	.D(n4167), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5379), 
	.D(n4166), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5356), 
	.D(n4165), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5350), 
	.D(n4164), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5316), 
	.D(n4163), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5315), 
	.D(n4162), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5292), 
	.D(n4161), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5286), 
	.D(n4160), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5252), 
	.D(n4159), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5251), 
	.D(n4158), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5228), 
	.D(n4157), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5222), 
	.D(n4156), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5188), 
	.D(n4155), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5187), 
	.D(n4154), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5164), 
	.D(n4153), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5158), 
	.D(n4152), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5124), 
	.Q(\UUT/regfile/reg_out[19][0] ), 
	.D(n4151), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5123), 
	.Q(\UUT/regfile/reg_out[19][10] ), 
	.D(n4150), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5100), 
	.Q(\UUT/regfile/reg_out[19][31] ), 
	.D(n4149), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5094), 
	.Q(\UUT/regfile/reg_out[19][8] ), 
	.D(n4148), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5028), 
	.Q(\UUT/regfile/reg_out[21][0] ), 
	.D(n4147), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5027), 
	.Q(\UUT/regfile/reg_out[21][10] ), 
	.D(n4146), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5004), 
	.Q(\UUT/regfile/reg_out[21][31] ), 
	.D(n4145), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4998), 
	.Q(\UUT/regfile/reg_out[21][8] ), 
	.D(n4144), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4964), 
	.D(n4143), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4963), 
	.D(n4142), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4940), 
	.D(n4141), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4934), 
	.D(n4140), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4900), 
	.Q(\UUT/regfile/reg_out[25][0] ), 
	.D(n4139), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4899), 
	.Q(\UUT/regfile/reg_out[25][10] ), 
	.D(n4138), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4876), 
	.Q(\UUT/regfile/reg_out[25][31] ), 
	.D(n4137), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4870), 
	.Q(\UUT/regfile/reg_out[25][8] ), 
	.D(n4136), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4836), 
	.D(n4135), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4835), 
	.D(n4134), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4812), 
	.D(n4133), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4806), 
	.D(n4132), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4772), 
	.Q(\UUT/regfile/reg_out[29][0] ), 
	.D(n4131), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4771), 
	.Q(\UUT/regfile/reg_out[29][10] ), 
	.D(n4130), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4748), 
	.Q(\UUT/regfile/reg_out[29][31] ), 
	.D(n4129), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4742), 
	.Q(\UUT/regfile/reg_out[29][8] ), 
	.D(n4128), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4676), 
	.D(n4127), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4675), 
	.D(n4126), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4652), 
	.D(n4125), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4646), 
	.D(n4124), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4740), 
	.D(n4123), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4739), 
	.D(n4122), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4716), 
	.D(n4121), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4710), 
	.D(n4120), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4612), 
	.Q(\UUT/regfile/reg_out[4][0] ), 
	.D(n4119), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4611), 
	.Q(\UUT/regfile/reg_out[4][10] ), 
	.D(n4118), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4588), 
	.Q(\UUT/regfile/reg_out[4][31] ), 
	.D(n4117), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4582), 
	.Q(\UUT/regfile/reg_out[4][8] ), 
	.D(n4116), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4548), 
	.D(n4115), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4547), 
	.D(n4114), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4524), 
	.D(n4113), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4518), 
	.D(n4112), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4484), 
	.D(n4111), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4483), 
	.D(n4110), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4460), 
	.D(n4109), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4454), 
	.D(n4108), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5412), 
	.D(n4107), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5411), 
	.D(n4106), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5388), 
	.D(n4105), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5382), 
	.D(n4104), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5348), 
	.D(n4103), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5347), 
	.D(n4102), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5324), 
	.D(n4101), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5318), 
	.D(n4100), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5284), 
	.D(n4099), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5283), 
	.D(n4098), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5260), 
	.D(n4097), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5254), 
	.D(n4096), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5220), 
	.D(n4095), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5219), 
	.D(n4094), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5196), 
	.D(n4093), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5190), 
	.D(n4092), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5156), 
	.Q(\UUT/regfile/reg_out[18][0] ), 
	.D(n4091), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5155), 
	.Q(\UUT/regfile/reg_out[18][10] ), 
	.D(n4090), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5132), 
	.Q(\UUT/regfile/reg_out[18][31] ), 
	.D(n4089), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5126), 
	.Q(\UUT/regfile/reg_out[18][8] ), 
	.D(n4088), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5060), 
	.Q(\UUT/regfile/reg_out[20][0] ), 
	.D(n4087), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5059), 
	.Q(\UUT/regfile/reg_out[20][10] ), 
	.D(n4086), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5036), 
	.Q(\UUT/regfile/reg_out[20][31] ), 
	.D(n4085), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5030), 
	.Q(\UUT/regfile/reg_out[20][8] ), 
	.D(n4084), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4996), 
	.D(n4083), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4995), 
	.D(n4082), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4972), 
	.D(n4081), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4966), 
	.D(n4080), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4932), 
	.Q(\UUT/regfile/reg_out[24][0] ), 
	.D(n4079), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4931), 
	.Q(\UUT/regfile/reg_out[24][10] ), 
	.D(n4078), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4908), 
	.Q(\UUT/regfile/reg_out[24][31] ), 
	.D(n4077), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4902), 
	.Q(\UUT/regfile/reg_out[24][8] ), 
	.D(n4076), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4868), 
	.D(n4075), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4867), 
	.D(n4074), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4844), 
	.D(n4073), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4838), 
	.D(n4072), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4804), 
	.Q(\UUT/regfile/reg_out[28][0] ), 
	.D(n4071), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4803), 
	.Q(\UUT/regfile/reg_out[28][10] ), 
	.D(n4070), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4780), 
	.Q(\UUT/regfile/reg_out[28][31] ), 
	.D(n4069), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4774), 
	.Q(\UUT/regfile/reg_out[28][8] ), 
	.D(n4068), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4708), 
	.D(n4067), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4707), 
	.D(n4066), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4684), 
	.D(n4065), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4678), 
	.D(n4064), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[SIGN]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_memhandle/N235 ), 
	.Q(\UUT/m_mem_command[SIGN] ), 
	.D(n4063), 
	.CK(CLK));
   DFFR_X1 \localbus/c2_op_reg[OP][0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\localbus/N293 ), 
	.D(\localbus/c1_op[OP][0] ), 
	.CK(CLK));
   DFFR_X1 \localbus/c2_op_reg[OP][1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\localbus/c2_op[OP][1] ), 
	.D(\localbus/c1_op[OP][1] ), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MH]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_memhandle/N238 ), 
	.D(n4059), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MB]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_memhandle/N236 ), 
	.D(n4058), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[31] ), 
	.D(n4056), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5629), 
	.D(n4055), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5628), 
	.Q(\UUT/Mpath/the_mult/acc_out[31] ), 
	.D(n4054), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/N116 ), 
	.Q(\UUT/exe_outsel [1]), 
	.D(n4053), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_exe_outsel1_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/N112 ), 
	.Q(\UUT/exe_outsel [0]), 
	.D(n4052), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_shift/N104 ), 
	.Q(\UUT/shift_op [2]), 
	.D(n4051), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_shift/N112 ), 
	.Q(\UUT/shift_op [1]), 
	.D(n4050), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_shift_op1_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_shift/N105 ), 
	.Q(\UUT/shift_op [0]), 
	.D(n4049), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N466 ), 
	.Q(\UUT/Alu_command[OP][5] ), 
	.D(n4048), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N453 ), 
	.Q(\UUT/Alu_command[OP][4] ), 
	.D(n4047), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2730), 
	.Q(\UUT/Alu_command[OP][3] ), 
	.D(n4046), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2729), 
	.Q(\UUT/Alu_command[OP][2] ), 
	.D(n4045), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N467 ), 
	.Q(\UUT/Alu_command[OP][1] ), 
	.D(n4044), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/ir_dx/out_alu_command_reg[OP][0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N468 ), 
	.Q(\UUT/Alu_command[OP][0] ), 
	.D(n4043), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[9]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2728), 
	.Q(\UUT/Mcontrol/f_currpc [9]), 
	.D(n4042), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[23]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2727), 
	.Q(\UUT/Mcontrol/f_currpc [23]), 
	.D(n4041), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[0] ), 
	.D(n4040), 
	.CK(CLK));
   DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2725), 
	.Q(\UUT/Mcontrol/f_currpc [0]), 
	.D(n4039), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[1] ), 
	.D(n4038), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[2] ), 
	.D(n4037), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[3] ), 
	.D(n4036), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[4] ), 
	.D(n4035), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[5] ), 
	.D(n4034), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[6] ), 
	.D(n4033), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[7] ), 
	.D(n4032), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[8] ), 
	.D(n4031), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[9] ), 
	.D(n4030), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[10] ), 
	.D(n4029), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[11] ), 
	.D(n4028), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[12] ), 
	.D(n4027), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[13] ), 
	.D(n4026), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[14] ), 
	.D(n4025), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[15] ), 
	.D(n4024), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[16] ), 
	.D(n4023), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[17] ), 
	.D(n4022), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[18] ), 
	.D(n4021), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[19] ), 
	.D(n4020), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[20] ), 
	.D(n4019), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[21] ), 
	.D(n4018), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[22] ), 
	.D(n4017), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/JAR/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/out_jar[23] ), 
	.D(n4016), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5482), 
	.D(n4015), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5458), 
	.D(n4013), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4429), 
	.D(n4012), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4461), 
	.D(n4011), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4493), 
	.D(n4010), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4525), 
	.D(n4009), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4557), 
	.Q(\UUT/regfile/reg_out[5][30] ), 
	.D(n4008), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4589), 
	.Q(\UUT/regfile/reg_out[4][30] ), 
	.D(n4007), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4621), 
	.D(n4006), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4653), 
	.D(n4005), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4685), 
	.D(n4004), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4717), 
	.D(n4003), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4749), 
	.Q(\UUT/regfile/reg_out[29][30] ), 
	.D(n4002), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4781), 
	.Q(\UUT/regfile/reg_out[28][30] ), 
	.D(n4001), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4813), 
	.D(n4000), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4845), 
	.D(n3999), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4877), 
	.Q(\UUT/regfile/reg_out[25][30] ), 
	.D(n3998), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4909), 
	.Q(\UUT/regfile/reg_out[24][30] ), 
	.D(n3997), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4941), 
	.D(n3996), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4973), 
	.D(n3995), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5005), 
	.Q(\UUT/regfile/reg_out[21][30] ), 
	.D(n3994), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5037), 
	.Q(\UUT/regfile/reg_out[20][30] ), 
	.D(n3993), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5069), 
	.D(n3992), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5101), 
	.Q(\UUT/regfile/reg_out[19][30] ), 
	.D(n3991), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5133), 
	.Q(\UUT/regfile/reg_out[18][30] ), 
	.D(n3990), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5165), 
	.D(n3989), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5197), 
	.D(n3988), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5229), 
	.D(n3987), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5261), 
	.D(n3986), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5293), 
	.D(n3985), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5325), 
	.D(n3984), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5357), 
	.D(n3983), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5389), 
	.D(n3982), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[30] ), 
	.D(n3980), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5631), 
	.D(n3979), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5630), 
	.Q(\UUT/Mpath/the_mult/acc_out[30] ), 
	.D(n3978), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5686), 
	.Q(\UUT/Mpath/the_mult/acc_out[62] ), 
	.D(n3977), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N24 ), 
	.Q(\UUT/Mpath/out_regB[30] ), 
	.D(n3976), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5464), 
	.D(n3975), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4431), 
	.D(n3974), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4463), 
	.D(n3973), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4495), 
	.D(n3972), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4527), 
	.D(n3971), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4559), 
	.Q(\UUT/regfile/reg_out[5][29] ), 
	.D(n3970), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4591), 
	.Q(\UUT/regfile/reg_out[4][29] ), 
	.D(n3969), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4623), 
	.D(n3968), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4655), 
	.D(n3967), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4687), 
	.D(n3966), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4719), 
	.D(n3965), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4751), 
	.Q(\UUT/regfile/reg_out[29][29] ), 
	.D(n3964), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4783), 
	.Q(\UUT/regfile/reg_out[28][29] ), 
	.D(n3963), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4815), 
	.D(n3962), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4847), 
	.D(n3961), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4879), 
	.Q(\UUT/regfile/reg_out[25][29] ), 
	.D(n3960), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4911), 
	.Q(\UUT/regfile/reg_out[24][29] ), 
	.D(n3959), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4943), 
	.D(n3958), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4975), 
	.D(n3957), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5007), 
	.Q(\UUT/regfile/reg_out[21][29] ), 
	.D(n3956), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5039), 
	.Q(\UUT/regfile/reg_out[20][29] ), 
	.D(n3955), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5071), 
	.D(n3954), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5103), 
	.Q(\UUT/regfile/reg_out[19][29] ), 
	.D(n3953), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5135), 
	.Q(\UUT/regfile/reg_out[18][29] ), 
	.D(n3952), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5167), 
	.D(n3951), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5199), 
	.D(n3950), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5231), 
	.D(n3949), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5263), 
	.D(n3948), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5295), 
	.D(n3947), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5327), 
	.D(n3946), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5359), 
	.D(n3945), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5391), 
	.D(n3944), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5467), 
	.D(n3942), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4432), 
	.D(n3941), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4464), 
	.D(n3940), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4496), 
	.D(n3939), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4528), 
	.D(n3938), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4560), 
	.Q(\UUT/regfile/reg_out[5][28] ), 
	.D(n3937), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4592), 
	.Q(\UUT/regfile/reg_out[4][28] ), 
	.D(n3936), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4624), 
	.D(n3935), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4656), 
	.D(n3934), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4688), 
	.D(n3933), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4720), 
	.D(n3932), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4752), 
	.Q(\UUT/regfile/reg_out[29][28] ), 
	.D(n3931), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4784), 
	.Q(\UUT/regfile/reg_out[28][28] ), 
	.D(n3930), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4816), 
	.D(n3929), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4848), 
	.D(n3928), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4880), 
	.Q(\UUT/regfile/reg_out[25][28] ), 
	.D(n3927), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4912), 
	.Q(\UUT/regfile/reg_out[24][28] ), 
	.D(n3926), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4944), 
	.D(n3925), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4976), 
	.D(n3924), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5008), 
	.Q(\UUT/regfile/reg_out[21][28] ), 
	.D(n3923), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5040), 
	.Q(\UUT/regfile/reg_out[20][28] ), 
	.D(n3922), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5072), 
	.D(n3921), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5104), 
	.Q(\UUT/regfile/reg_out[19][28] ), 
	.D(n3920), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5136), 
	.Q(\UUT/regfile/reg_out[18][28] ), 
	.D(n3919), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5168), 
	.D(n3918), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5200), 
	.D(n3917), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5232), 
	.D(n3916), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5264), 
	.D(n3915), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5296), 
	.D(n3914), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5328), 
	.D(n3913), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5360), 
	.D(n3912), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5392), 
	.D(n3911), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5470), 
	.D(n3909), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4433), 
	.D(n3908), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4465), 
	.D(n3907), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4497), 
	.D(n3906), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4529), 
	.D(n3905), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4561), 
	.Q(\UUT/regfile/reg_out[5][27] ), 
	.D(n3904), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4593), 
	.Q(\UUT/regfile/reg_out[4][27] ), 
	.D(n3903), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4625), 
	.D(n3902), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4657), 
	.D(n3901), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4689), 
	.D(n3900), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4721), 
	.D(n3899), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4753), 
	.Q(\UUT/regfile/reg_out[29][27] ), 
	.D(n3898), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4785), 
	.Q(\UUT/regfile/reg_out[28][27] ), 
	.D(n3897), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4817), 
	.D(n3896), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4849), 
	.D(n3895), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4881), 
	.Q(\UUT/regfile/reg_out[25][27] ), 
	.D(n3894), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4913), 
	.Q(\UUT/regfile/reg_out[24][27] ), 
	.D(n3893), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4945), 
	.D(n3892), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4977), 
	.D(n3891), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5009), 
	.Q(\UUT/regfile/reg_out[21][27] ), 
	.D(n3890), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5041), 
	.Q(\UUT/regfile/reg_out[20][27] ), 
	.D(n3889), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5073), 
	.D(n3888), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5105), 
	.Q(\UUT/regfile/reg_out[19][27] ), 
	.D(n3887), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5137), 
	.Q(\UUT/regfile/reg_out[18][27] ), 
	.D(n3886), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5169), 
	.D(n3885), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5201), 
	.D(n3884), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5233), 
	.D(n3883), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5265), 
	.D(n3882), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5297), 
	.D(n3881), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5329), 
	.D(n3880), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5361), 
	.D(n3879), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5393), 
	.D(n3878), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5473), 
	.D(n3876), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4434), 
	.D(n3875), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4466), 
	.D(n3874), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4498), 
	.D(n3873), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4530), 
	.D(n3872), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4562), 
	.Q(\UUT/regfile/reg_out[5][26] ), 
	.D(n3871), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4594), 
	.Q(\UUT/regfile/reg_out[4][26] ), 
	.D(n3870), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4626), 
	.D(n3869), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4658), 
	.D(n3868), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4690), 
	.D(n3867), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4722), 
	.D(n3866), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4754), 
	.Q(\UUT/regfile/reg_out[29][26] ), 
	.D(n3865), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4786), 
	.Q(\UUT/regfile/reg_out[28][26] ), 
	.D(n3864), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4818), 
	.D(n3863), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4850), 
	.D(n3862), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4882), 
	.Q(\UUT/regfile/reg_out[25][26] ), 
	.D(n3861), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4914), 
	.Q(\UUT/regfile/reg_out[24][26] ), 
	.D(n3860), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4946), 
	.D(n3859), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4978), 
	.D(n3858), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5010), 
	.Q(\UUT/regfile/reg_out[21][26] ), 
	.D(n3857), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5042), 
	.Q(\UUT/regfile/reg_out[20][26] ), 
	.D(n3856), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5074), 
	.D(n3855), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5106), 
	.Q(\UUT/regfile/reg_out[19][26] ), 
	.D(n3854), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5138), 
	.Q(\UUT/regfile/reg_out[18][26] ), 
	.D(n3853), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5170), 
	.D(n3852), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5202), 
	.D(n3851), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5234), 
	.D(n3850), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5266), 
	.D(n3849), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5298), 
	.D(n3848), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5330), 
	.D(n3847), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5362), 
	.D(n3846), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5394), 
	.D(n3845), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5476), 
	.D(n3843), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4435), 
	.D(n3842), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4467), 
	.D(n3841), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4499), 
	.D(n3840), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4531), 
	.D(n3839), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4563), 
	.Q(\UUT/regfile/reg_out[5][25] ), 
	.D(n3838), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4595), 
	.Q(\UUT/regfile/reg_out[4][25] ), 
	.D(n3837), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4627), 
	.D(n3836), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4659), 
	.D(n3835), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4691), 
	.D(n3834), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4723), 
	.D(n3833), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4755), 
	.Q(\UUT/regfile/reg_out[29][25] ), 
	.D(n3832), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4787), 
	.Q(\UUT/regfile/reg_out[28][25] ), 
	.D(n3831), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4819), 
	.D(n3830), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4851), 
	.D(n3829), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4883), 
	.Q(\UUT/regfile/reg_out[25][25] ), 
	.D(n3828), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4915), 
	.Q(\UUT/regfile/reg_out[24][25] ), 
	.D(n3827), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4947), 
	.D(n3826), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4979), 
	.D(n3825), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5011), 
	.Q(\UUT/regfile/reg_out[21][25] ), 
	.D(n3824), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5043), 
	.Q(\UUT/regfile/reg_out[20][25] ), 
	.D(n3823), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5075), 
	.D(n3822), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5107), 
	.Q(\UUT/regfile/reg_out[19][25] ), 
	.D(n3821), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5139), 
	.Q(\UUT/regfile/reg_out[18][25] ), 
	.D(n3820), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5171), 
	.D(n3819), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5203), 
	.D(n3818), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5235), 
	.D(n3817), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5267), 
	.D(n3816), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5299), 
	.D(n3815), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5331), 
	.D(n3814), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5363), 
	.D(n3813), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5395), 
	.D(n3812), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5494), 
	.D(n3810), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N82 ), 
	.Q(\UUT/Mpath/out_regB[1] ), 
	.D(n3809), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regMaddr/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_memhandle/N239 ), 
	.Q(\UUT/Mpath/mem_baddr [1]), 
	.D(n3808), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4437), 
	.D(n3807), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4469), 
	.D(n3806), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4501), 
	.D(n3805), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4533), 
	.D(n3804), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4565), 
	.Q(\UUT/regfile/reg_out[5][23] ), 
	.D(n3803), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4597), 
	.Q(\UUT/regfile/reg_out[4][23] ), 
	.D(n3802), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4629), 
	.D(n3801), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4661), 
	.D(n3800), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4693), 
	.D(n3799), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4725), 
	.D(n3798), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4757), 
	.Q(\UUT/regfile/reg_out[29][23] ), 
	.D(n3797), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4789), 
	.Q(\UUT/regfile/reg_out[28][23] ), 
	.D(n3796), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4821), 
	.D(n3795), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4853), 
	.D(n3794), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4885), 
	.Q(\UUT/regfile/reg_out[25][23] ), 
	.D(n3793), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4917), 
	.Q(\UUT/regfile/reg_out[24][23] ), 
	.D(n3792), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4949), 
	.D(n3791), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4981), 
	.D(n3790), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5013), 
	.Q(\UUT/regfile/reg_out[21][23] ), 
	.D(n3789), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5045), 
	.Q(\UUT/regfile/reg_out[20][23] ), 
	.D(n3788), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5077), 
	.D(n3787), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5109), 
	.Q(\UUT/regfile/reg_out[19][23] ), 
	.D(n3786), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5141), 
	.Q(\UUT/regfile/reg_out[18][23] ), 
	.D(n3785), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5173), 
	.D(n3784), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5205), 
	.D(n3783), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5237), 
	.D(n3782), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5269), 
	.D(n3781), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5301), 
	.D(n3780), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5333), 
	.D(n3779), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5365), 
	.D(n3778), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5397), 
	.D(n3777), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[23] ), 
	.D(n3775), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5647), 
	.D(n3774), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5646), 
	.Q(\UUT/Mpath/the_mult/acc_out[23] ), 
	.D(n3773), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5694), 
	.Q(\UUT/Mpath/the_mult/acc_out[55] ), 
	.D(n3772), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4441), 
	.D(n3771), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4473), 
	.D(n3770), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4505), 
	.D(n3769), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4537), 
	.D(n3768), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4569), 
	.Q(\UUT/regfile/reg_out[5][1] ), 
	.D(n3767), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4601), 
	.Q(\UUT/regfile/reg_out[4][1] ), 
	.D(n3766), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4633), 
	.D(n3765), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4665), 
	.D(n3764), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4697), 
	.D(n3763), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4729), 
	.D(n3762), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4761), 
	.Q(\UUT/regfile/reg_out[29][1] ), 
	.D(n3761), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4793), 
	.Q(\UUT/regfile/reg_out[28][1] ), 
	.D(n3760), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4825), 
	.D(n3759), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4857), 
	.D(n3758), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4889), 
	.Q(\UUT/regfile/reg_out[25][1] ), 
	.D(n3757), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4921), 
	.Q(\UUT/regfile/reg_out[24][1] ), 
	.D(n3756), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4953), 
	.D(n3755), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4985), 
	.D(n3754), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5017), 
	.Q(\UUT/regfile/reg_out[21][1] ), 
	.D(n3753), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5049), 
	.Q(\UUT/regfile/reg_out[20][1] ), 
	.D(n3752), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5081), 
	.D(n3751), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5113), 
	.Q(\UUT/regfile/reg_out[19][1] ), 
	.D(n3750), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5145), 
	.Q(\UUT/regfile/reg_out[18][1] ), 
	.D(n3749), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5177), 
	.D(n3748), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5209), 
	.D(n3747), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5241), 
	.D(n3746), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5273), 
	.D(n3745), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5305), 
	.D(n3744), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5337), 
	.D(n3743), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5369), 
	.D(n3742), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5401), 
	.D(n3741), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[1] ), 
	.D(n3739), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5655), 
	.D(n3738), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5654), 
	.Q(\UUT/Mpath/the_mult/acc_out[1] ), 
	.D(n3737), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5698), 
	.Q(\UUT/Mpath/the_mult/acc_out[33] ), 
	.D(n3736), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [1]), 
	.D(n3734), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5461), 
	.D(n3733), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4430), 
	.D(n3732), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4462), 
	.D(n3731), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4494), 
	.D(n3730), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4526), 
	.D(n3729), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4558), 
	.Q(\UUT/regfile/reg_out[5][2] ), 
	.D(n3728), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4590), 
	.Q(\UUT/regfile/reg_out[4][2] ), 
	.D(n3727), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4622), 
	.D(n3726), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4654), 
	.D(n3725), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4686), 
	.D(n3724), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4718), 
	.D(n3723), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4750), 
	.Q(\UUT/regfile/reg_out[29][2] ), 
	.D(n3722), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4782), 
	.Q(\UUT/regfile/reg_out[28][2] ), 
	.D(n3721), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4814), 
	.D(n3720), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4846), 
	.D(n3719), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4878), 
	.Q(\UUT/regfile/reg_out[25][2] ), 
	.D(n3718), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4910), 
	.Q(\UUT/regfile/reg_out[24][2] ), 
	.D(n3717), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4942), 
	.D(n3716), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4974), 
	.D(n3715), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5006), 
	.Q(\UUT/regfile/reg_out[21][2] ), 
	.D(n3714), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5038), 
	.Q(\UUT/regfile/reg_out[20][2] ), 
	.D(n3713), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5070), 
	.D(n3712), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5102), 
	.Q(\UUT/regfile/reg_out[19][2] ), 
	.D(n3711), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5134), 
	.Q(\UUT/regfile/reg_out[18][2] ), 
	.D(n3710), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5166), 
	.D(n3709), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5198), 
	.D(n3708), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5230), 
	.D(n3707), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5262), 
	.D(n3706), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5294), 
	.D(n3705), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5326), 
	.D(n3704), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5358), 
	.D(n3703), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5390), 
	.D(n3702), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[2] ), 
	.D(n3700), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5633), 
	.D(n3699), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5632), 
	.Q(\UUT/Mpath/the_mult/acc_out[2] ), 
	.D(n3698), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5687), 
	.Q(\UUT/Mpath/the_mult/acc_out[34] ), 
	.D(n3697), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N80 ), 
	.Q(\UUT/Mpath/out_regB[2] ), 
	.D(n3696), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [2]), 
	.D(n3695), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[2]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2694), 
	.Q(\UUT/Mcontrol/f_currpc [2]), 
	.D(n3694), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5452), 
	.D(n3693), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4427), 
	.D(n3692), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4459), 
	.D(n3691), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4491), 
	.D(n3690), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4523), 
	.D(n3689), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4555), 
	.Q(\UUT/regfile/reg_out[5][3] ), 
	.D(n3688), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4587), 
	.Q(\UUT/regfile/reg_out[4][3] ), 
	.D(n3687), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4619), 
	.D(n3686), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4651), 
	.D(n3685), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4683), 
	.D(n3684), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4715), 
	.D(n3683), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4747), 
	.Q(\UUT/regfile/reg_out[29][3] ), 
	.D(n3682), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4779), 
	.Q(\UUT/regfile/reg_out[28][3] ), 
	.D(n3681), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4811), 
	.D(n3680), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4843), 
	.D(n3679), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4875), 
	.Q(\UUT/regfile/reg_out[25][3] ), 
	.D(n3678), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4907), 
	.Q(\UUT/regfile/reg_out[24][3] ), 
	.D(n3677), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4939), 
	.D(n3676), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4971), 
	.D(n3675), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5003), 
	.Q(\UUT/regfile/reg_out[21][3] ), 
	.D(n3674), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5035), 
	.Q(\UUT/regfile/reg_out[20][3] ), 
	.D(n3673), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5067), 
	.D(n3672), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5099), 
	.Q(\UUT/regfile/reg_out[19][3] ), 
	.D(n3671), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5131), 
	.Q(\UUT/regfile/reg_out[18][3] ), 
	.D(n3670), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5163), 
	.D(n3669), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5195), 
	.D(n3668), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5227), 
	.D(n3667), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5259), 
	.D(n3666), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5291), 
	.D(n3665), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5323), 
	.D(n3664), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5355), 
	.D(n3663), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5387), 
	.D(n3662), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[3] ), 
	.D(n3660), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5627), 
	.D(n3659), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5626), 
	.Q(\UUT/Mpath/the_mult/acc_out[3] ), 
	.D(n3658), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5684), 
	.Q(\UUT/Mpath/the_mult/acc_out[35] ), 
	.D(n3657), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N78 ), 
	.Q(\UUT/Mpath/out_regB[3] ), 
	.D(n3656), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [3]), 
	.D(n3655), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[3]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2691), 
	.Q(\UUT/Mcontrol/f_currpc [3]), 
	.D(n3654), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5449), 
	.D(n3653), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4426), 
	.D(n3652), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4458), 
	.D(n3651), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4490), 
	.D(n3650), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4522), 
	.D(n3649), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4554), 
	.Q(\UUT/regfile/reg_out[5][4] ), 
	.D(n3648), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4586), 
	.Q(\UUT/regfile/reg_out[4][4] ), 
	.D(n3647), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4618), 
	.D(n3646), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4650), 
	.D(n3645), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4682), 
	.D(n3644), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4714), 
	.D(n3643), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4746), 
	.Q(\UUT/regfile/reg_out[29][4] ), 
	.D(n3642), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4778), 
	.Q(\UUT/regfile/reg_out[28][4] ), 
	.D(n3641), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4810), 
	.D(n3640), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4842), 
	.D(n3639), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4874), 
	.Q(\UUT/regfile/reg_out[25][4] ), 
	.D(n3638), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4906), 
	.Q(\UUT/regfile/reg_out[24][4] ), 
	.D(n3637), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4938), 
	.D(n3636), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4970), 
	.D(n3635), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5002), 
	.Q(\UUT/regfile/reg_out[21][4] ), 
	.D(n3634), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5034), 
	.Q(\UUT/regfile/reg_out[20][4] ), 
	.D(n3633), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5066), 
	.D(n3632), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5098), 
	.Q(\UUT/regfile/reg_out[19][4] ), 
	.D(n3631), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5130), 
	.Q(\UUT/regfile/reg_out[18][4] ), 
	.D(n3630), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5162), 
	.D(n3629), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5194), 
	.D(n3628), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5226), 
	.D(n3627), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5258), 
	.D(n3626), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5290), 
	.D(n3625), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5322), 
	.D(n3624), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5354), 
	.D(n3623), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5386), 
	.D(n3622), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[4] ), 
	.D(n3620), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5625), 
	.D(n3619), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5624), 
	.Q(\UUT/Mpath/the_mult/acc_out[4] ), 
	.D(n3618), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5683), 
	.Q(\UUT/Mpath/the_mult/acc_out[36] ), 
	.D(n3617), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N76 ), 
	.Q(\UUT/Mpath/out_regB[4] ), 
	.D(n3616), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [4]), 
	.D(n3615), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[4]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2688), 
	.Q(\UUT/Mcontrol/f_currpc [4]), 
	.D(n3614), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5446), 
	.D(n3613), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4425), 
	.D(n3612), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4457), 
	.D(n3611), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4489), 
	.D(n3610), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4521), 
	.D(n3609), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4553), 
	.Q(\UUT/regfile/reg_out[5][5] ), 
	.D(n3608), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4585), 
	.Q(\UUT/regfile/reg_out[4][5] ), 
	.D(n3607), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4617), 
	.D(n3606), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4649), 
	.D(n3605), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4681), 
	.D(n3604), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4713), 
	.D(n3603), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4745), 
	.Q(\UUT/regfile/reg_out[29][5] ), 
	.D(n3602), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4777), 
	.Q(\UUT/regfile/reg_out[28][5] ), 
	.D(n3601), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4809), 
	.D(n3600), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4841), 
	.D(n3599), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4873), 
	.Q(\UUT/regfile/reg_out[25][5] ), 
	.D(n3598), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4905), 
	.Q(\UUT/regfile/reg_out[24][5] ), 
	.D(n3597), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4937), 
	.D(n3596), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4969), 
	.D(n3595), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5001), 
	.Q(\UUT/regfile/reg_out[21][5] ), 
	.D(n3594), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5033), 
	.Q(\UUT/regfile/reg_out[20][5] ), 
	.D(n3593), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5065), 
	.D(n3592), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5097), 
	.Q(\UUT/regfile/reg_out[19][5] ), 
	.D(n3591), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5129), 
	.Q(\UUT/regfile/reg_out[18][5] ), 
	.D(n3590), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5161), 
	.D(n3589), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5193), 
	.D(n3588), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5225), 
	.D(n3587), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5257), 
	.D(n3586), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5289), 
	.D(n3585), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5321), 
	.D(n3584), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5353), 
	.D(n3583), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5385), 
	.D(n3582), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[5] ), 
	.D(n3580), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5623), 
	.D(n3579), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5622), 
	.Q(\UUT/Mpath/the_mult/acc_out[5] ), 
	.D(n3578), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5682), 
	.Q(\UUT/Mpath/the_mult/acc_out[37] ), 
	.D(n3577), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [5]), 
	.D(n3575), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5443), 
	.D(n3573), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4424), 
	.D(n3572), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4456), 
	.D(n3571), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4488), 
	.D(n3570), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4520), 
	.D(n3569), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4552), 
	.Q(\UUT/regfile/reg_out[5][6] ), 
	.D(n3568), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4584), 
	.Q(\UUT/regfile/reg_out[4][6] ), 
	.D(n3567), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4616), 
	.D(n3566), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4648), 
	.D(n3565), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4680), 
	.D(n3564), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4712), 
	.D(n3563), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4744), 
	.Q(\UUT/regfile/reg_out[29][6] ), 
	.D(n3562), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4776), 
	.Q(\UUT/regfile/reg_out[28][6] ), 
	.D(n3561), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4808), 
	.D(n3560), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4840), 
	.D(n3559), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4872), 
	.Q(\UUT/regfile/reg_out[25][6] ), 
	.D(n3558), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4904), 
	.Q(\UUT/regfile/reg_out[24][6] ), 
	.D(n3557), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4936), 
	.D(n3556), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4968), 
	.D(n3555), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5000), 
	.Q(\UUT/regfile/reg_out[21][6] ), 
	.D(n3554), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5032), 
	.Q(\UUT/regfile/reg_out[20][6] ), 
	.D(n3553), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5064), 
	.D(n3552), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5096), 
	.Q(\UUT/regfile/reg_out[19][6] ), 
	.D(n3551), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5128), 
	.Q(\UUT/regfile/reg_out[18][6] ), 
	.D(n3550), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5160), 
	.D(n3549), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5192), 
	.D(n3548), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5224), 
	.D(n3547), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5256), 
	.D(n3546), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5288), 
	.D(n3545), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5320), 
	.D(n3544), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5352), 
	.D(n3543), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5384), 
	.D(n3542), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[6] ), 
	.D(n3540), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5621), 
	.D(n3539), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5620), 
	.Q(\UUT/Mpath/the_mult/acc_out[6] ), 
	.D(n3538), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5681), 
	.Q(\UUT/Mpath/the_mult/acc_out[38] ), 
	.D(n3537), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N72 ), 
	.Q(\UUT/Mpath/out_regB[6] ), 
	.D(n3536), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [6]), 
	.D(n3535), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[6]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2682), 
	.Q(\UUT/Mcontrol/f_currpc [6]), 
	.D(n3534), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5440), 
	.D(n3533), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4423), 
	.D(n3532), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4455), 
	.D(n3531), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4487), 
	.D(n3530), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4519), 
	.D(n3529), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4551), 
	.Q(\UUT/regfile/reg_out[5][7] ), 
	.D(n3528), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4583), 
	.Q(\UUT/regfile/reg_out[4][7] ), 
	.D(n3527), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4615), 
	.D(n3526), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4647), 
	.D(n3525), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4679), 
	.D(n3524), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4711), 
	.D(n3523), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4743), 
	.Q(\UUT/regfile/reg_out[29][7] ), 
	.D(n3522), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4775), 
	.Q(\UUT/regfile/reg_out[28][7] ), 
	.D(n3521), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4807), 
	.D(n3520), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4839), 
	.D(n3519), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4871), 
	.Q(\UUT/regfile/reg_out[25][7] ), 
	.D(n3518), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4903), 
	.Q(\UUT/regfile/reg_out[24][7] ), 
	.D(n3517), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4935), 
	.D(n3516), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4967), 
	.D(n3515), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4999), 
	.Q(\UUT/regfile/reg_out[21][7] ), 
	.D(n3514), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5031), 
	.Q(\UUT/regfile/reg_out[20][7] ), 
	.D(n3513), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5063), 
	.D(n3512), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5095), 
	.Q(\UUT/regfile/reg_out[19][7] ), 
	.D(n3511), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5127), 
	.Q(\UUT/regfile/reg_out[18][7] ), 
	.D(n3510), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5159), 
	.D(n3509), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5191), 
	.D(n3508), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5223), 
	.D(n3507), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5255), 
	.D(n3506), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5287), 
	.D(n3505), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5319), 
	.D(n3504), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5351), 
	.D(n3503), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5383), 
	.D(n3502), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[7] ), 
	.D(n3500), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5619), 
	.D(n3499), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5618), 
	.Q(\UUT/Mpath/the_mult/acc_out[7] ), 
	.D(n3498), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5680), 
	.Q(\UUT/Mpath/the_mult/acc_out[39] ), 
	.D(n3497), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N70 ), 
	.Q(\UUT/Mpath/out_regB[7] ), 
	.D(n3496), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [7]), 
	.D(n3495), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[7]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2679), 
	.Q(\UUT/Mcontrol/f_currpc [7]), 
	.D(n3494), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5437), 
	.D(n3493), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[8] ), 
	.D(n3491), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5617), 
	.D(n3490), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5616), 
	.Q(\UUT/Mpath/the_mult/acc_out[8] ), 
	.D(n3489), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5679), 
	.Q(\UUT/Mpath/the_mult/acc_out[40] ), 
	.D(n3488), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[8]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2677), 
	.Q(\UUT/Mcontrol/f_currpc [8]), 
	.D(n3487), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5433), 
	.D(n3486), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4421), 
	.D(n3485), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4453), 
	.D(n3484), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4485), 
	.D(n3483), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4517), 
	.D(n3482), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4549), 
	.Q(\UUT/regfile/reg_out[5][9] ), 
	.D(n3481), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4581), 
	.Q(\UUT/regfile/reg_out[4][9] ), 
	.D(n3480), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4613), 
	.D(n3479), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4645), 
	.D(n3478), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4677), 
	.D(n3477), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4709), 
	.D(n3476), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4741), 
	.Q(\UUT/regfile/reg_out[29][9] ), 
	.D(n3475), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4773), 
	.Q(\UUT/regfile/reg_out[28][9] ), 
	.D(n3474), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4805), 
	.D(n3473), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4837), 
	.D(n3472), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4869), 
	.Q(\UUT/regfile/reg_out[25][9] ), 
	.D(n3471), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4901), 
	.Q(\UUT/regfile/reg_out[24][9] ), 
	.D(n3470), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4933), 
	.D(n3469), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4965), 
	.D(n3468), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4997), 
	.Q(\UUT/regfile/reg_out[21][9] ), 
	.D(n3467), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5029), 
	.Q(\UUT/regfile/reg_out[20][9] ), 
	.D(n3466), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5061), 
	.D(n3465), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5093), 
	.Q(\UUT/regfile/reg_out[19][9] ), 
	.D(n3464), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5125), 
	.Q(\UUT/regfile/reg_out[18][9] ), 
	.D(n3463), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5157), 
	.D(n3462), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5189), 
	.D(n3461), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5221), 
	.D(n3460), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5253), 
	.D(n3459), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5285), 
	.D(n3458), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5317), 
	.D(n3457), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5349), 
	.D(n3456), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5381), 
	.D(n3455), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[9] ), 
	.D(n3453), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5615), 
	.D(n3452), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5614), 
	.Q(\UUT/Mpath/the_mult/acc_out[9] ), 
	.D(n3451), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5678), 
	.Q(\UUT/Mpath/the_mult/acc_out[41] ), 
	.D(n3450), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N66 ), 
	.Q(\UUT/Mpath/out_regB[9] ), 
	.D(n3449), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [9]), 
	.D(n3448), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5524), 
	.D(n3447), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[10] ), 
	.D(n3445), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5675), 
	.D(n3444), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5674), 
	.Q(\UUT/Mpath/the_mult/acc_out[10] ), 
	.D(n3443), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5708), 
	.Q(\UUT/Mpath/the_mult/acc_out[42] ), 
	.D(n3442), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5521), 
	.D(n3441), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4450), 
	.D(n3440), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4482), 
	.D(n3439), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4514), 
	.D(n3438), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4546), 
	.D(n3437), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4578), 
	.Q(\UUT/regfile/reg_out[5][11] ), 
	.D(n3436), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4610), 
	.Q(\UUT/regfile/reg_out[4][11] ), 
	.D(n3435), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4642), 
	.D(n3434), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4674), 
	.D(n3433), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4706), 
	.D(n3432), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4738), 
	.D(n3431), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4770), 
	.Q(\UUT/regfile/reg_out[29][11] ), 
	.D(n3430), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4802), 
	.Q(\UUT/regfile/reg_out[28][11] ), 
	.D(n3429), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4834), 
	.D(n3428), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4866), 
	.D(n3427), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4898), 
	.Q(\UUT/regfile/reg_out[25][11] ), 
	.D(n3426), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4930), 
	.Q(\UUT/regfile/reg_out[24][11] ), 
	.D(n3425), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4962), 
	.D(n3424), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4994), 
	.D(n3423), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5026), 
	.Q(\UUT/regfile/reg_out[21][11] ), 
	.D(n3422), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5058), 
	.Q(\UUT/regfile/reg_out[20][11] ), 
	.D(n3421), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5090), 
	.D(n3420), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5122), 
	.Q(\UUT/regfile/reg_out[19][11] ), 
	.D(n3419), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5154), 
	.Q(\UUT/regfile/reg_out[18][11] ), 
	.D(n3418), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5186), 
	.D(n3417), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5218), 
	.D(n3416), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5250), 
	.D(n3415), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5282), 
	.D(n3414), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5314), 
	.D(n3413), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5346), 
	.D(n3412), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5378), 
	.D(n3411), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5410), 
	.D(n3410), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[11] ), 
	.D(n3408), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5673), 
	.D(n3407), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5672), 
	.Q(\UUT/Mpath/the_mult/acc_out[11] ), 
	.D(n3406), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5707), 
	.Q(\UUT/Mpath/the_mult/acc_out[43] ), 
	.D(n3405), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [11]), 
	.D(n3403), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[11]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2671), 
	.Q(\UUT/Mcontrol/f_currpc [11]), 
	.D(n3402), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5518), 
	.D(n3401), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4449), 
	.D(n3400), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4481), 
	.D(n3399), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4513), 
	.D(n3398), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4545), 
	.D(n3397), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4577), 
	.Q(\UUT/regfile/reg_out[5][12] ), 
	.D(n3396), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4609), 
	.Q(\UUT/regfile/reg_out[4][12] ), 
	.D(n3395), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4641), 
	.D(n3394), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4673), 
	.D(n3393), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4705), 
	.D(n3392), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4737), 
	.D(n3391), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4769), 
	.Q(\UUT/regfile/reg_out[29][12] ), 
	.D(n3390), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4801), 
	.Q(\UUT/regfile/reg_out[28][12] ), 
	.D(n3389), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4833), 
	.D(n3388), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4865), 
	.D(n3387), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4897), 
	.Q(\UUT/regfile/reg_out[25][12] ), 
	.D(n3386), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4929), 
	.Q(\UUT/regfile/reg_out[24][12] ), 
	.D(n3385), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4961), 
	.D(n3384), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4993), 
	.D(n3383), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5025), 
	.Q(\UUT/regfile/reg_out[21][12] ), 
	.D(n3382), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5057), 
	.Q(\UUT/regfile/reg_out[20][12] ), 
	.D(n3381), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5089), 
	.D(n3380), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5121), 
	.Q(\UUT/regfile/reg_out[19][12] ), 
	.D(n3379), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5153), 
	.Q(\UUT/regfile/reg_out[18][12] ), 
	.D(n3378), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5185), 
	.D(n3377), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5217), 
	.D(n3376), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5249), 
	.D(n3375), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5281), 
	.D(n3374), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5313), 
	.D(n3373), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5345), 
	.D(n3372), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5377), 
	.D(n3371), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5409), 
	.D(n3370), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[12] ), 
	.D(n3368), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5671), 
	.D(n3367), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5670), 
	.Q(\UUT/Mpath/the_mult/acc_out[12] ), 
	.D(n3366), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5706), 
	.Q(\UUT/Mpath/the_mult/acc_out[44] ), 
	.D(n3365), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [12]), 
	.D(n3363), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[12]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2668), 
	.Q(\UUT/Mcontrol/f_currpc [12]), 
	.D(n3362), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5515), 
	.D(n3361), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4448), 
	.D(n3360), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4480), 
	.D(n3359), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4512), 
	.D(n3358), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4544), 
	.D(n3357), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4576), 
	.Q(\UUT/regfile/reg_out[5][13] ), 
	.D(n3356), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4608), 
	.Q(\UUT/regfile/reg_out[4][13] ), 
	.D(n3355), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4640), 
	.D(n3354), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4672), 
	.D(n3353), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4704), 
	.D(n3352), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4736), 
	.D(n3351), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4768), 
	.Q(\UUT/regfile/reg_out[29][13] ), 
	.D(n3350), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4800), 
	.Q(\UUT/regfile/reg_out[28][13] ), 
	.D(n3349), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4832), 
	.D(n3348), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4864), 
	.D(n3347), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4896), 
	.Q(\UUT/regfile/reg_out[25][13] ), 
	.D(n3346), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4928), 
	.Q(\UUT/regfile/reg_out[24][13] ), 
	.D(n3345), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4960), 
	.D(n3344), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4992), 
	.D(n3343), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5024), 
	.Q(\UUT/regfile/reg_out[21][13] ), 
	.D(n3342), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5056), 
	.Q(\UUT/regfile/reg_out[20][13] ), 
	.D(n3341), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5088), 
	.D(n3340), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5120), 
	.Q(\UUT/regfile/reg_out[19][13] ), 
	.D(n3339), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5152), 
	.Q(\UUT/regfile/reg_out[18][13] ), 
	.D(n3338), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5184), 
	.D(n3337), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5216), 
	.D(n3336), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5248), 
	.D(n3335), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5280), 
	.D(n3334), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5312), 
	.D(n3333), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5344), 
	.D(n3332), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5376), 
	.D(n3331), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5408), 
	.D(n3330), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[13] ), 
	.D(n3328), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5669), 
	.D(n3327), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5668), 
	.Q(\UUT/Mpath/the_mult/acc_out[13] ), 
	.D(n3326), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5705), 
	.Q(\UUT/Mpath/the_mult/acc_out[45] ), 
	.D(n3325), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[13]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2666), 
	.Q(\UUT/Mcontrol/f_currpc [13]), 
	.D(n3323), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [13]), 
	.D(n3322), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5512), 
	.D(n3321), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4447), 
	.D(n3320), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4479), 
	.D(n3319), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4511), 
	.D(n3318), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4543), 
	.D(n3317), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4575), 
	.Q(\UUT/regfile/reg_out[5][14] ), 
	.D(n3316), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4607), 
	.Q(\UUT/regfile/reg_out[4][14] ), 
	.D(n3315), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4639), 
	.D(n3314), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4671), 
	.D(n3313), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4703), 
	.D(n3312), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4735), 
	.D(n3311), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4767), 
	.Q(\UUT/regfile/reg_out[29][14] ), 
	.D(n3310), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4799), 
	.Q(\UUT/regfile/reg_out[28][14] ), 
	.D(n3309), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4831), 
	.D(n3308), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4863), 
	.D(n3307), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4895), 
	.Q(\UUT/regfile/reg_out[25][14] ), 
	.D(n3306), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4927), 
	.Q(\UUT/regfile/reg_out[24][14] ), 
	.D(n3305), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4959), 
	.D(n3304), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4991), 
	.D(n3303), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5023), 
	.Q(\UUT/regfile/reg_out[21][14] ), 
	.D(n3302), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5055), 
	.Q(\UUT/regfile/reg_out[20][14] ), 
	.D(n3301), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5087), 
	.D(n3300), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5119), 
	.Q(\UUT/regfile/reg_out[19][14] ), 
	.D(n3299), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5151), 
	.Q(\UUT/regfile/reg_out[18][14] ), 
	.D(n3298), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5183), 
	.D(n3297), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5215), 
	.D(n3296), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5247), 
	.D(n3295), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5279), 
	.D(n3294), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5311), 
	.D(n3293), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5343), 
	.D(n3292), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5375), 
	.D(n3291), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5407), 
	.D(n3290), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[14] ), 
	.D(n3288), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5667), 
	.D(n3287), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5666), 
	.Q(\UUT/Mpath/the_mult/acc_out[14] ), 
	.D(n3286), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5704), 
	.Q(\UUT/Mpath/the_mult/acc_out[46] ), 
	.D(n3285), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[14]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2663), 
	.Q(\UUT/Mcontrol/f_currpc [14]), 
	.D(n3283), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [14]), 
	.D(n3282), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5509), 
	.D(n3281), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4446), 
	.D(n3280), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4478), 
	.D(n3279), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4510), 
	.D(n3278), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4542), 
	.D(n3277), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4574), 
	.Q(\UUT/regfile/reg_out[5][15] ), 
	.D(n3276), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4606), 
	.Q(\UUT/regfile/reg_out[4][15] ), 
	.D(n3275), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4638), 
	.D(n3274), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4670), 
	.D(n3273), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4702), 
	.D(n3272), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4734), 
	.D(n3271), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4766), 
	.Q(\UUT/regfile/reg_out[29][15] ), 
	.D(n3270), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4798), 
	.Q(\UUT/regfile/reg_out[28][15] ), 
	.D(n3269), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4830), 
	.D(n3268), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4862), 
	.D(n3267), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4894), 
	.Q(\UUT/regfile/reg_out[25][15] ), 
	.D(n3266), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4926), 
	.Q(\UUT/regfile/reg_out[24][15] ), 
	.D(n3265), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4958), 
	.D(n3264), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4990), 
	.D(n3263), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5022), 
	.Q(\UUT/regfile/reg_out[21][15] ), 
	.D(n3262), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5054), 
	.Q(\UUT/regfile/reg_out[20][15] ), 
	.D(n3261), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5086), 
	.D(n3260), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5118), 
	.Q(\UUT/regfile/reg_out[19][15] ), 
	.D(n3259), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5150), 
	.Q(\UUT/regfile/reg_out[18][15] ), 
	.D(n3258), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5182), 
	.D(n3257), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5214), 
	.D(n3256), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5246), 
	.D(n3255), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5278), 
	.D(n3254), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5310), 
	.D(n3253), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5342), 
	.D(n3252), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5374), 
	.D(n3251), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5406), 
	.D(n3250), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[15] ), 
	.D(n3248), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5665), 
	.D(n3247), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5664), 
	.Q(\UUT/Mpath/the_mult/acc_out[15] ), 
	.D(n3246), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5703), 
	.Q(\UUT/Mpath/the_mult/acc_out[47] ), 
	.D(n3245), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [15]), 
	.D(n3242), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5506), 
	.D(n3241), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4445), 
	.D(n3240), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4477), 
	.D(n3239), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4509), 
	.D(n3238), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4541), 
	.D(n3237), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4573), 
	.Q(\UUT/regfile/reg_out[5][16] ), 
	.D(n3236), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4605), 
	.Q(\UUT/regfile/reg_out[4][16] ), 
	.D(n3235), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4637), 
	.D(n3234), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4669), 
	.D(n3233), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4701), 
	.D(n3232), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4733), 
	.D(n3231), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4765), 
	.Q(\UUT/regfile/reg_out[29][16] ), 
	.D(n3230), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4797), 
	.Q(\UUT/regfile/reg_out[28][16] ), 
	.D(n3229), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4829), 
	.D(n3228), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4861), 
	.D(n3227), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4893), 
	.Q(\UUT/regfile/reg_out[25][16] ), 
	.D(n3226), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4925), 
	.Q(\UUT/regfile/reg_out[24][16] ), 
	.D(n3225), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4957), 
	.D(n3224), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4989), 
	.D(n3223), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5021), 
	.Q(\UUT/regfile/reg_out[21][16] ), 
	.D(n3222), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5053), 
	.Q(\UUT/regfile/reg_out[20][16] ), 
	.D(n3221), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5085), 
	.D(n3220), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5117), 
	.Q(\UUT/regfile/reg_out[19][16] ), 
	.D(n3219), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5149), 
	.Q(\UUT/regfile/reg_out[18][16] ), 
	.D(n3218), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5181), 
	.D(n3217), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5213), 
	.D(n3216), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5245), 
	.D(n3215), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5277), 
	.D(n3214), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5309), 
	.D(n3213), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5341), 
	.D(n3212), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5373), 
	.D(n3211), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5405), 
	.D(n3210), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[16] ), 
	.D(n3208), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5663), 
	.D(n3207), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5662), 
	.Q(\UUT/Mpath/the_mult/acc_out[16] ), 
	.D(n3206), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5702), 
	.Q(\UUT/Mpath/the_mult/acc_out[48] ), 
	.D(n3205), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[16]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2657), 
	.Q(\UUT/Mcontrol/f_currpc [16]), 
	.D(n3203), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [16]), 
	.D(n3202), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5503), 
	.D(n3201), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4444), 
	.D(n3200), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4476), 
	.D(n3199), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4508), 
	.D(n3198), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4540), 
	.D(n3197), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4572), 
	.Q(\UUT/regfile/reg_out[5][17] ), 
	.D(n3196), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4604), 
	.Q(\UUT/regfile/reg_out[4][17] ), 
	.D(n3195), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4636), 
	.D(n3194), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4668), 
	.D(n3193), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4700), 
	.D(n3192), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4732), 
	.D(n3191), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4764), 
	.Q(\UUT/regfile/reg_out[29][17] ), 
	.D(n3190), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4796), 
	.Q(\UUT/regfile/reg_out[28][17] ), 
	.D(n3189), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4828), 
	.D(n3188), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4860), 
	.D(n3187), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4892), 
	.Q(\UUT/regfile/reg_out[25][17] ), 
	.D(n3186), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4924), 
	.Q(\UUT/regfile/reg_out[24][17] ), 
	.D(n3185), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4956), 
	.D(n3184), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4988), 
	.D(n3183), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5020), 
	.Q(\UUT/regfile/reg_out[21][17] ), 
	.D(n3182), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5052), 
	.Q(\UUT/regfile/reg_out[20][17] ), 
	.D(n3181), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5084), 
	.D(n3180), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5116), 
	.Q(\UUT/regfile/reg_out[19][17] ), 
	.D(n3179), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5148), 
	.Q(\UUT/regfile/reg_out[18][17] ), 
	.D(n3178), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5180), 
	.D(n3177), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5212), 
	.D(n3176), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5244), 
	.D(n3175), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5276), 
	.D(n3174), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5308), 
	.D(n3173), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5340), 
	.D(n3172), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5372), 
	.D(n3171), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5404), 
	.D(n3170), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[17] ), 
	.D(n3168), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5661), 
	.D(n3167), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5660), 
	.Q(\UUT/Mpath/the_mult/acc_out[17] ), 
	.D(n3166), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5701), 
	.Q(\UUT/Mpath/the_mult/acc_out[49] ), 
	.D(n3165), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[17]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2654), 
	.Q(\UUT/Mcontrol/f_currpc [17]), 
	.D(n3163), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [17]), 
	.D(n3162), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5500), 
	.D(n3161), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4443), 
	.D(n3160), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4475), 
	.D(n3159), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4507), 
	.D(n3158), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4539), 
	.D(n3157), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4571), 
	.Q(\UUT/regfile/reg_out[5][18] ), 
	.D(n3156), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4603), 
	.Q(\UUT/regfile/reg_out[4][18] ), 
	.D(n3155), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4635), 
	.D(n3154), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4667), 
	.D(n3153), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4699), 
	.D(n3152), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4731), 
	.D(n3151), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4763), 
	.Q(\UUT/regfile/reg_out[29][18] ), 
	.D(n3150), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4795), 
	.Q(\UUT/regfile/reg_out[28][18] ), 
	.D(n3149), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4827), 
	.D(n3148), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4859), 
	.D(n3147), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4891), 
	.Q(\UUT/regfile/reg_out[25][18] ), 
	.D(n3146), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4923), 
	.Q(\UUT/regfile/reg_out[24][18] ), 
	.D(n3145), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4955), 
	.D(n3144), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4987), 
	.D(n3143), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5019), 
	.Q(\UUT/regfile/reg_out[21][18] ), 
	.D(n3142), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5051), 
	.Q(\UUT/regfile/reg_out[20][18] ), 
	.D(n3141), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5083), 
	.D(n3140), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5115), 
	.Q(\UUT/regfile/reg_out[19][18] ), 
	.D(n3139), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5147), 
	.Q(\UUT/regfile/reg_out[18][18] ), 
	.D(n3138), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5179), 
	.D(n3137), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5211), 
	.D(n3136), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5243), 
	.D(n3135), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5275), 
	.D(n3134), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5307), 
	.D(n3133), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5339), 
	.D(n3132), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5371), 
	.D(n3131), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5403), 
	.D(n3130), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[18] ), 
	.D(n3128), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5659), 
	.D(n3127), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5658), 
	.Q(\UUT/Mpath/the_mult/acc_out[18] ), 
	.D(n3126), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5700), 
	.Q(\UUT/Mpath/the_mult/acc_out[50] ), 
	.D(n3125), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [18]), 
	.D(n3122), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5497), 
	.D(n3121), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4442), 
	.D(n3120), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4474), 
	.D(n3119), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4506), 
	.D(n3118), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4538), 
	.D(n3117), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4570), 
	.Q(\UUT/regfile/reg_out[5][19] ), 
	.D(n3116), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4602), 
	.Q(\UUT/regfile/reg_out[4][19] ), 
	.D(n3115), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4634), 
	.D(n3114), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4666), 
	.D(n3113), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4698), 
	.D(n3112), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4730), 
	.D(n3111), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4762), 
	.Q(\UUT/regfile/reg_out[29][19] ), 
	.D(n3110), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4794), 
	.Q(\UUT/regfile/reg_out[28][19] ), 
	.D(n3109), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4826), 
	.D(n3108), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4858), 
	.D(n3107), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4890), 
	.Q(\UUT/regfile/reg_out[25][19] ), 
	.D(n3106), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4922), 
	.Q(\UUT/regfile/reg_out[24][19] ), 
	.D(n3105), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4954), 
	.D(n3104), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4986), 
	.D(n3103), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5018), 
	.Q(\UUT/regfile/reg_out[21][19] ), 
	.D(n3102), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5050), 
	.Q(\UUT/regfile/reg_out[20][19] ), 
	.D(n3101), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5082), 
	.D(n3100), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5114), 
	.Q(\UUT/regfile/reg_out[19][19] ), 
	.D(n3099), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5146), 
	.Q(\UUT/regfile/reg_out[18][19] ), 
	.D(n3098), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5178), 
	.D(n3097), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5210), 
	.D(n3096), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5242), 
	.D(n3095), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5274), 
	.D(n3094), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5306), 
	.D(n3093), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5338), 
	.D(n3092), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5370), 
	.D(n3091), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5402), 
	.D(n3090), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[19] ), 
	.D(n3088), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5657), 
	.D(n3087), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5656), 
	.Q(\UUT/Mpath/the_mult/acc_out[19] ), 
	.D(n3086), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5699), 
	.Q(\UUT/Mpath/the_mult/acc_out[51] ), 
	.D(n3085), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[19]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2648), 
	.Q(\UUT/Mcontrol/f_currpc [19]), 
	.D(n3083), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [19]), 
	.D(n3082), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5491), 
	.D(n3081), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4440), 
	.D(n3080), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4472), 
	.D(n3079), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4504), 
	.D(n3078), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4536), 
	.D(n3077), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4568), 
	.Q(\UUT/regfile/reg_out[5][20] ), 
	.D(n3076), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4600), 
	.Q(\UUT/regfile/reg_out[4][20] ), 
	.D(n3075), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4632), 
	.D(n3074), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4664), 
	.D(n3073), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4696), 
	.D(n3072), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4728), 
	.D(n3071), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4760), 
	.Q(\UUT/regfile/reg_out[29][20] ), 
	.D(n3070), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4792), 
	.Q(\UUT/regfile/reg_out[28][20] ), 
	.D(n3069), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4824), 
	.D(n3068), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4856), 
	.D(n3067), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4888), 
	.Q(\UUT/regfile/reg_out[25][20] ), 
	.D(n3066), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4920), 
	.Q(\UUT/regfile/reg_out[24][20] ), 
	.D(n3065), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4952), 
	.D(n3064), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4984), 
	.D(n3063), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5016), 
	.Q(\UUT/regfile/reg_out[21][20] ), 
	.D(n3062), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5048), 
	.Q(\UUT/regfile/reg_out[20][20] ), 
	.D(n3061), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5080), 
	.D(n3060), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5112), 
	.Q(\UUT/regfile/reg_out[19][20] ), 
	.D(n3059), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5144), 
	.Q(\UUT/regfile/reg_out[18][20] ), 
	.D(n3058), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5176), 
	.D(n3057), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5208), 
	.D(n3056), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5240), 
	.D(n3055), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5272), 
	.D(n3054), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5304), 
	.D(n3053), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5336), 
	.D(n3052), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5368), 
	.D(n3051), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5400), 
	.D(n3050), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[20] ), 
	.D(n3048), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5653), 
	.D(n3047), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5652), 
	.Q(\UUT/Mpath/the_mult/acc_out[20] ), 
	.D(n3046), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5697), 
	.Q(\UUT/Mpath/the_mult/acc_out[52] ), 
	.D(n3045), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[20]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2645), 
	.Q(\UUT/Mcontrol/f_currpc [20]), 
	.D(n3043), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [20]), 
	.D(n3042), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5488), 
	.D(n3041), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4439), 
	.D(n3040), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4471), 
	.D(n3039), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4503), 
	.D(n3038), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4535), 
	.D(n3037), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4567), 
	.Q(\UUT/regfile/reg_out[5][21] ), 
	.D(n3036), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4599), 
	.Q(\UUT/regfile/reg_out[4][21] ), 
	.D(n3035), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4631), 
	.D(n3034), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4663), 
	.D(n3033), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4695), 
	.D(n3032), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4727), 
	.D(n3031), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4759), 
	.Q(\UUT/regfile/reg_out[29][21] ), 
	.D(n3030), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4791), 
	.Q(\UUT/regfile/reg_out[28][21] ), 
	.D(n3029), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4823), 
	.D(n3028), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4855), 
	.D(n3027), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4887), 
	.Q(\UUT/regfile/reg_out[25][21] ), 
	.D(n3026), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4919), 
	.Q(\UUT/regfile/reg_out[24][21] ), 
	.D(n3025), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4951), 
	.D(n3024), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4983), 
	.D(n3023), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5015), 
	.Q(\UUT/regfile/reg_out[21][21] ), 
	.D(n3022), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5047), 
	.Q(\UUT/regfile/reg_out[20][21] ), 
	.D(n3021), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5079), 
	.D(n3020), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5111), 
	.Q(\UUT/regfile/reg_out[19][21] ), 
	.D(n3019), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5143), 
	.Q(\UUT/regfile/reg_out[18][21] ), 
	.D(n3018), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5175), 
	.D(n3017), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5207), 
	.D(n3016), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5239), 
	.D(n3015), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5271), 
	.D(n3014), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5303), 
	.D(n3013), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5335), 
	.D(n3012), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5367), 
	.D(n3011), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5399), 
	.D(n3010), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[21] ), 
	.D(n3008), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5651), 
	.D(n3007), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5650), 
	.Q(\UUT/Mpath/the_mult/acc_out[21] ), 
	.D(n3006), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5696), 
	.Q(\UUT/Mpath/the_mult/acc_out[53] ), 
	.D(n3005), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[21]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2642), 
	.Q(\UUT/Mcontrol/f_currpc [21]), 
	.D(n3003), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [21]), 
	.D(n3002), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5485), 
	.D(n3001), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4438), 
	.D(n3000), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4470), 
	.D(n2999), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4502), 
	.D(n2998), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4534), 
	.D(n2997), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4566), 
	.Q(\UUT/regfile/reg_out[5][22] ), 
	.D(n2996), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4598), 
	.Q(\UUT/regfile/reg_out[4][22] ), 
	.D(n2995), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4630), 
	.D(n2994), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4662), 
	.D(n2993), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4694), 
	.D(n2992), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4726), 
	.D(n2991), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4758), 
	.Q(\UUT/regfile/reg_out[29][22] ), 
	.D(n2990), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4790), 
	.Q(\UUT/regfile/reg_out[28][22] ), 
	.D(n2989), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4822), 
	.D(n2988), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4854), 
	.D(n2987), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4886), 
	.Q(\UUT/regfile/reg_out[25][22] ), 
	.D(n2986), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4918), 
	.Q(\UUT/regfile/reg_out[24][22] ), 
	.D(n2985), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4950), 
	.D(n2984), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4982), 
	.D(n2983), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5014), 
	.Q(\UUT/regfile/reg_out[21][22] ), 
	.D(n2982), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5046), 
	.Q(\UUT/regfile/reg_out[20][22] ), 
	.D(n2981), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5078), 
	.D(n2980), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5110), 
	.Q(\UUT/regfile/reg_out[19][22] ), 
	.D(n2979), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5142), 
	.Q(\UUT/regfile/reg_out[18][22] ), 
	.D(n2978), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5174), 
	.D(n2977), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5206), 
	.D(n2976), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5238), 
	.D(n2975), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5270), 
	.D(n2974), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5302), 
	.D(n2973), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5334), 
	.D(n2972), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5366), 
	.D(n2971), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5398), 
	.D(n2970), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[22] ), 
	.D(n2968), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5649), 
	.D(n2967), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5648), 
	.Q(\UUT/Mpath/the_mult/acc_out[22] ), 
	.D(n2966), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5695), 
	.Q(\UUT/Mpath/the_mult/acc_out[54] ), 
	.D(n2965), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[22]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2639), 
	.Q(\UUT/Mcontrol/f_currpc [22]), 
	.D(n2963), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [22]), 
	.D(n2962), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regM/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5479), 
	.D(n2961), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_9/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4436), 
	.D(n2960), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_8/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4468), 
	.D(n2959), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_7/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4500), 
	.D(n2958), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_6/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4532), 
	.D(n2957), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_5/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4564), 
	.Q(\UUT/regfile/reg_out[5][24] ), 
	.D(n2956), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_4/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4596), 
	.Q(\UUT/regfile/reg_out[4][24] ), 
	.D(n2955), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_3/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4628), 
	.D(n2954), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_31/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4660), 
	.D(n2953), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_30/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4692), 
	.D(n2952), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_2/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4724), 
	.D(n2951), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_29/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4756), 
	.Q(\UUT/regfile/reg_out[29][24] ), 
	.D(n2950), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_28/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4788), 
	.Q(\UUT/regfile/reg_out[28][24] ), 
	.D(n2949), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_27/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4820), 
	.D(n2948), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_26/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4852), 
	.D(n2947), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_25/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4884), 
	.Q(\UUT/regfile/reg_out[25][24] ), 
	.D(n2946), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_24/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4916), 
	.Q(\UUT/regfile/reg_out[24][24] ), 
	.D(n2945), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_23/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4948), 
	.D(n2944), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_22/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4980), 
	.D(n2943), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_21/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5012), 
	.Q(\UUT/regfile/reg_out[21][24] ), 
	.D(n2942), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_20/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5044), 
	.Q(\UUT/regfile/reg_out[20][24] ), 
	.D(n2941), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_1/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5076), 
	.D(n2940), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_19/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5108), 
	.Q(\UUT/regfile/reg_out[19][24] ), 
	.D(n2939), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_18/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5140), 
	.Q(\UUT/regfile/reg_out[18][24] ), 
	.D(n2938), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_17/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5172), 
	.D(n2937), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_16/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5204), 
	.D(n2936), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_15/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5236), 
	.D(n2935), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_14/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5268), 
	.D(n2934), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_13/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5300), 
	.D(n2933), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_12/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5332), 
	.D(n2932), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_11/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5364), 
	.D(n2931), 
	.CK(CLK));
   DFFR_X1 \UUT/regfile/rx_10/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5396), 
	.D(n2930), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[24] ), 
	.D(n2928), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5645), 
	.D(n2927), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5644), 
	.Q(\UUT/Mpath/the_mult/acc_out[24] ), 
	.D(n2926), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5693), 
	.Q(\UUT/Mpath/the_mult/acc_out[56] ), 
	.D(n2925), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [24]), 
	.D(n2923), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[25] ), 
	.D(n2922), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5643), 
	.D(n2921), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5642), 
	.Q(\UUT/Mpath/the_mult/acc_out[25] ), 
	.D(n2920), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5692), 
	.Q(\UUT/Mpath/the_mult/acc_out[57] ), 
	.D(n2919), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [25]), 
	.D(n2917), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[26] ), 
	.D(n2916), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5641), 
	.D(n2915), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5640), 
	.Q(\UUT/Mpath/the_mult/acc_out[26] ), 
	.D(n2914), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5691), 
	.Q(\UUT/Mpath/the_mult/acc_out[58] ), 
	.D(n2913), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [26]), 
	.D(n2911), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[27] ), 
	.D(n2910), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5639), 
	.D(n2909), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5638), 
	.Q(\UUT/Mpath/the_mult/acc_out[27] ), 
	.D(n2908), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5690), 
	.Q(\UUT/Mpath/the_mult/acc_out[59] ), 
	.D(n2907), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [27]), 
	.D(n2905), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[28] ), 
	.D(n2904), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5637), 
	.D(n2903), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5636), 
	.Q(\UUT/Mpath/the_mult/acc_out[28] ), 
	.D(n2902), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5689), 
	.Q(\UUT/Mpath/the_mult/acc_out[60] ), 
	.D(n2901), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [28]), 
	.D(n2899), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multa/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand1[29] ), 
	.D(n2898), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/Pipe_mtvalue_reg/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5635), 
	.D(n2897), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulLo_reg/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5634), 
	.Q(\UUT/Mpath/the_mult/acc_out[29] ), 
	.D(n2896), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5688), 
	.Q(\UUT/Mpath/the_mult/acc_out[61] ), 
	.D(n2895), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regB/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N26 ), 
	.Q(\UUT/Mpath/out_regB[29] ), 
	.D(n2894), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [29]), 
	.D(n2893), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [30]), 
	.D(n2892), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [23]), 
	.D(n2891), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2623), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[31] ), 
	.D(n2890), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2622), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[30] ), 
	.D(n2889), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2621), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[29] ), 
	.D(n2888), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2620), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[28] ), 
	.D(n2887), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2619), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[27] ), 
	.D(n2886), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2618), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[26] ), 
	.D(n2885), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2617), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[25] ), 
	.D(n2884), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2616), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[24] ), 
	.D(n2883), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2615), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[23] ), 
	.D(n2882), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2614), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[22] ), 
	.D(n2881), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2613), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[21] ), 
	.D(n2880), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2612), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[20] ), 
	.D(n2879), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2611), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[19] ), 
	.D(n2878), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2610), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[18] ), 
	.D(n2877), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2609), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[17] ), 
	.D(n2876), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2608), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[16] ), 
	.D(n2875), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2607), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
	.D(n2874), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2606), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
	.D(n2873), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2605), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
	.D(n2872), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2604), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
	.D(n2871), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2603), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
	.D(n2870), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2602), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
	.D(n2869), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2601), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[9] ), 
	.D(n2868), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2600), 
	.Q(\UUT/Mpath/the_memhandle/smdr_out[8] ), 
	.D(n2867), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4380), 
	.Q(D_DATA_OUTBUS[7]), 
	.D(n2866), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4381), 
	.Q(D_DATA_OUTBUS[6]), 
	.D(n2865), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4382), 
	.Q(D_DATA_OUTBUS[5]), 
	.D(n2864), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4383), 
	.Q(D_DATA_OUTBUS[4]), 
	.D(n2863), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4384), 
	.Q(D_DATA_OUTBUS[3]), 
	.D(n2862), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4387), 
	.Q(D_DATA_OUTBUS[2]), 
	.D(n2861), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4398), 
	.Q(D_DATA_OUTBUS[1]), 
	.D(n2860), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_memhandle/SMDR/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n4409), 
	.Q(D_DATA_OUTBUS[0]), 
	.D(n2859), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [8]), 
	.D(n2858), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [10]), 
	.D(n2857), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [31]), 
	.D(n2856), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/multb/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/x_operand2 [0]), 
	.D(n2855), 
	.CK(CLK));
   OAI221_X1 U3 (.ZN(n2855), 
	.C2(n71), 
	.C1(n70), 
	.B2(n69), 
	.B1(n68), 
	.A(n72));
   NAND2_X1 U4 (.ZN(n72), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN105_UUT_Mpath_the_mult_x_operand2_0_));
   OAI21_X1 U5 (.ZN(n2856), 
	.B2(FE_OFN8_n73), 
	.B1(n74), 
	.A(n75));
   NAND2_X1 U6 (.ZN(n75), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [31]));
   OAI221_X1 U7 (.ZN(n2857), 
	.C2(n71), 
	.C1(n77), 
	.B2(n69), 
	.B1(n76), 
	.A(n78));
   NAND2_X1 U8 (.ZN(n78), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [10]));
   OAI221_X1 U9 (.ZN(n2858), 
	.C2(n71), 
	.C1(n80), 
	.B2(n69), 
	.B1(n79), 
	.A(n81));
   NAND2_X1 U10 (.ZN(n81), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [8]));
   OAI22_X1 U11 (.ZN(n2859), 
	.B2(n83), 
	.B1(n70), 
	.A2(n82), 
	.A1(n4409));
   OAI22_X1 U12 (.ZN(n2860), 
	.B2(n83), 
	.B1(n84), 
	.A2(n82), 
	.A1(n4398));
   OAI22_X1 U13 (.ZN(n2861), 
	.B2(n83), 
	.B1(n85), 
	.A2(n82), 
	.A1(n4387));
   OAI22_X1 U14 (.ZN(n2862), 
	.B2(n83), 
	.B1(n86), 
	.A2(n82), 
	.A1(n4384));
   OAI22_X1 U15 (.ZN(n2863), 
	.B2(n83), 
	.B1(n87), 
	.A2(n82), 
	.A1(n4383));
   OAI22_X1 U16 (.ZN(n2864), 
	.B2(n83), 
	.B1(n88), 
	.A2(n82), 
	.A1(n4382));
   OAI22_X1 U48 (.ZN(n2865), 
	.B2(n83), 
	.B1(n89), 
	.A2(n82), 
	.A1(n4381));
   OAI22_X1 U49 (.ZN(n2866), 
	.B2(n83), 
	.B1(n90), 
	.A2(n82), 
	.A1(n4380));
   OAI22_X1 U50 (.ZN(n2867), 
	.B2(n83), 
	.B1(n80), 
	.A2(n2600), 
	.A1(n82));
   OAI22_X1 U51 (.ZN(n2868), 
	.B2(n83), 
	.B1(n91), 
	.A2(n2601), 
	.A1(n82));
   OAI22_X1 U52 (.ZN(n2869), 
	.B2(n83), 
	.B1(n77), 
	.A2(n2602), 
	.A1(n82));
   OAI22_X1 U53 (.ZN(n2870), 
	.B2(n83), 
	.B1(n92), 
	.A2(n2603), 
	.A1(n82));
   OAI22_X1 U54 (.ZN(n2871), 
	.B2(n83), 
	.B1(n93), 
	.A2(n2604), 
	.A1(n82));
   OAI22_X1 U55 (.ZN(n2872), 
	.B2(n83), 
	.B1(n94), 
	.A2(n2605), 
	.A1(n82));
   OAI22_X1 U56 (.ZN(n2873), 
	.B2(n83), 
	.B1(n95), 
	.A2(n2606), 
	.A1(n82));
   OAI22_X1 U57 (.ZN(n2874), 
	.B2(n83), 
	.B1(n96), 
	.A2(n2607), 
	.A1(n82));
   OAI22_X1 U58 (.ZN(n2875), 
	.B2(n83), 
	.B1(n97), 
	.A2(n2608), 
	.A1(n82));
   OAI22_X1 U59 (.ZN(n2876), 
	.B2(n83), 
	.B1(n98), 
	.A2(n2609), 
	.A1(n82));
   OAI22_X1 U60 (.ZN(n2877), 
	.B2(n83), 
	.B1(n99), 
	.A2(n2610), 
	.A1(n82));
   OAI22_X1 U61 (.ZN(n2878), 
	.B2(n83), 
	.B1(n100), 
	.A2(n2611), 
	.A1(n82));
   OAI22_X1 U62 (.ZN(n2879), 
	.B2(n83), 
	.B1(n101), 
	.A2(n2612), 
	.A1(n82));
   OAI22_X1 U63 (.ZN(n2880), 
	.B2(n83), 
	.B1(n102), 
	.A2(n2613), 
	.A1(n82));
   OAI22_X1 U64 (.ZN(n2881), 
	.B2(n83), 
	.B1(n103), 
	.A2(n2614), 
	.A1(n82));
   OAI22_X1 U65 (.ZN(n2882), 
	.B2(n83), 
	.B1(n104), 
	.A2(n2615), 
	.A1(n82));
   OAI22_X1 U66 (.ZN(n2883), 
	.B2(n83), 
	.B1(n105), 
	.A2(n2616), 
	.A1(n82));
   INV_X1 U67 (.ZN(n105), 
	.A(n106));
   OAI22_X1 U68 (.ZN(n2884), 
	.B2(n83), 
	.B1(n107), 
	.A2(n2617), 
	.A1(n82));
   INV_X1 U69 (.ZN(n107), 
	.A(n108));
   OAI22_X1 U70 (.ZN(n2885), 
	.B2(n83), 
	.B1(n109), 
	.A2(n2618), 
	.A1(n82));
   INV_X1 U71 (.ZN(n109), 
	.A(n110));
   OAI22_X1 U72 (.ZN(n2886), 
	.B2(n83), 
	.B1(n111), 
	.A2(n2619), 
	.A1(n82));
   OAI22_X1 U73 (.ZN(n2887), 
	.B2(n83), 
	.B1(n112), 
	.A2(n2620), 
	.A1(n82));
   OAI22_X1 U74 (.ZN(n2888), 
	.B2(n83), 
	.B1(n113), 
	.A2(n2621), 
	.A1(n82));
   OAI22_X1 U75 (.ZN(n2889), 
	.B2(n83), 
	.B1(n114), 
	.A2(n2622), 
	.A1(n82));
   OAI22_X1 U76 (.ZN(n2890), 
	.B2(n83), 
	.B1(n115), 
	.A2(n2623), 
	.A1(n82));
   OAI221_X1 U79 (.ZN(n2891), 
	.C2(n71), 
	.C1(n104), 
	.B2(n69), 
	.B1(FE_OFN102_n117), 
	.A(n118));
   NAND2_X1 U80 (.ZN(n118), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [23]));
   OAI221_X1 U81 (.ZN(n2892), 
	.C2(n71), 
	.C1(n114), 
	.B2(FE_OFN8_n73), 
	.B1(n119), 
	.A(n120));
   NAND2_X1 U82 (.ZN(n120), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [30]));
   OAI221_X1 U83 (.ZN(n2893), 
	.C2(n71), 
	.C1(n113), 
	.B2(FE_OFN8_n73), 
	.B1(n121), 
	.A(n122));
   NAND2_X1 U84 (.ZN(n122), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [29]));
   OAI222_X1 U85 (.ZN(n2894), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N26 ), 
	.B2(n121), 
	.B1(net54953), 
	.A2(n123), 
	.A1(n113));
   AOI21_X1 U86 (.ZN(n121), 
	.B2(n125), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [13]), 
	.A(n126));
   INV_X1 U87 (.ZN(n113), 
	.A(n127));
   OAI222_X1 U88 (.ZN(n127), 
	.C2(n132), 
	.C1(n5463), 
	.B2(n131), 
	.B1(n130), 
	.A2(n129), 
	.A1(FE_OFN24_n128));
   OAI221_X1 U91 (.ZN(n2896), 
	.C2(n142), 
	.C1(n5634), 
	.B2(n141), 
	.B1(n140), 
	.A(n143));
   AOI22_X1 U92 (.ZN(n143), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [29]), 
	.A2(n138), 
	.A1(n144));
   INV_X1 U93 (.ZN(n138), 
	.A(n5635));
   OAI22_X1 U94 (.ZN(n2897), 
	.B2(net54873), 
	.B1(n5635), 
	.A2(n146), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U95 (.ZN(n2898), 
	.B2(FE_OFN8_n73), 
	.B1(n148), 
	.A2(n146), 
	.A1(n147));
   INV_X1 U96 (.ZN(n146), 
	.A(FE_OFN113_UUT_Mpath_the_mult_x_operand1_29_));
   OAI221_X1 U97 (.ZN(n2899), 
	.C2(n71), 
	.C1(n112), 
	.B2(FE_OFN8_n73), 
	.B1(n149), 
	.A(n150));
   NAND2_X1 U98 (.ZN(n150), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [28]));
   OAI222_X1 U99 (.ZN(n2900), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N28 ), 
	.B2(n149), 
	.B1(net54953), 
	.A2(n123), 
	.A1(n112));
   AOI21_X1 U100 (.ZN(n149), 
	.B2(n125), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [12]), 
	.A(n126));
   INV_X1 U101 (.ZN(n112), 
	.A(n151));
   OAI222_X1 U102 (.ZN(n151), 
	.C2(n132), 
	.C1(n5466), 
	.B2(n131), 
	.B1(n153), 
	.A2(n129), 
	.A1(FE_OFN23_n152));
   OAI221_X1 U105 (.ZN(n2902), 
	.C2(n142), 
	.C1(n5636), 
	.B2(n157), 
	.B1(n140), 
	.A(n158));
   AOI22_X1 U106 (.ZN(n158), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [28]), 
	.A2(n156), 
	.A1(n144));
   INV_X1 U107 (.ZN(n156), 
	.A(n5637));
   OAI22_X1 U108 (.ZN(n2903), 
	.B2(net54875), 
	.B1(n5637), 
	.A2(n159), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U109 (.ZN(n2904), 
	.B2(FE_OFN8_n73), 
	.B1(n160), 
	.A2(n159), 
	.A1(n147));
   INV_X1 U110 (.ZN(n159), 
	.A(\UUT/Mpath/the_mult/x_operand1[28] ));
   OAI221_X1 U111 (.ZN(n2905), 
	.C2(n71), 
	.C1(n111), 
	.B2(FE_OFN8_n73), 
	.B1(n161), 
	.A(n162));
   NAND2_X1 U112 (.ZN(n162), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [27]));
   OAI222_X1 U113 (.ZN(n2906), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N30 ), 
	.B2(n161), 
	.B1(net54953), 
	.A2(n123), 
	.A1(n111));
   AOI21_X1 U114 (.ZN(n161), 
	.B2(n125), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [11]), 
	.A(n126));
   INV_X1 U115 (.ZN(n111), 
	.A(n163));
   OAI222_X1 U116 (.ZN(n163), 
	.C2(n132), 
	.C1(n5469), 
	.B2(n131), 
	.B1(n165), 
	.A2(n129), 
	.A1(FE_OFN22_n164));
   OAI221_X1 U117 (.ZN(n2907), 
	.C2(n135), 
	.C1(n5690), 
	.B2(n166), 
	.B1(n133), 
	.A(n167));
   AOI22_X1 U118 (.ZN(n167), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [59]), 
	.A2(n168), 
	.A1(n137));
   OAI221_X1 U119 (.ZN(n2908), 
	.C2(n142), 
	.C1(n5638), 
	.B2(n169), 
	.B1(n140), 
	.A(n170));
   AOI22_X1 U120 (.ZN(n170), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [27]), 
	.A2(n168), 
	.A1(n144));
   INV_X1 U121 (.ZN(n168), 
	.A(n5639));
   OAI22_X1 U122 (.ZN(n2909), 
	.B2(net54875), 
	.B1(n5639), 
	.A2(n171), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U123 (.ZN(n2910), 
	.B2(FE_OFN8_n73), 
	.B1(n172), 
	.A2(n171), 
	.A1(n147));
   INV_X1 U124 (.ZN(n171), 
	.A(FE_OFN117_UUT_Mpath_the_mult_x_operand1_27_));
   OAI21_X1 U125 (.ZN(n2911), 
	.B2(FE_OFN8_n73), 
	.B1(FE_OFN0_n173), 
	.A(n174));
   NAND2_X1 U126 (.ZN(n174), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [26]));
   OAI22_X1 U127 (.ZN(n2912), 
	.B2(FE_OFN0_n173), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N32 ));
   AOI211_X1 U128 (.ZN(n173), 
	.C2(n110), 
	.C1(n175), 
	.B(n177), 
	.A(n176));
   INV_X1 U129 (.ZN(n177), 
	.A(n178));
   AOI22_X1 U130 (.ZN(n178), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [10]), 
	.B1(n125), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [24]), 
	.A1(n179));
   OAI222_X1 U131 (.ZN(n110), 
	.C2(n132), 
	.C1(n5472), 
	.B2(n131), 
	.B1(n181), 
	.A2(n129), 
	.A1(FE_OFN26_n180));
   OAI221_X1 U132 (.ZN(n2913), 
	.C2(n135), 
	.C1(n5691), 
	.B2(n182), 
	.B1(n133), 
	.A(n183));
   AOI22_X1 U133 (.ZN(n183), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [58]), 
	.A2(n184), 
	.A1(n137));
   OAI221_X1 U134 (.ZN(n2914), 
	.C2(n142), 
	.C1(n5640), 
	.B2(n185), 
	.B1(n140), 
	.A(n186));
   AOI22_X1 U135 (.ZN(n186), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [26]), 
	.A2(n184), 
	.A1(n144));
   INV_X1 U136 (.ZN(n184), 
	.A(n5641));
   OAI22_X1 U137 (.ZN(n2915), 
	.B2(net54873), 
	.B1(n5641), 
	.A2(n187), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U138 (.ZN(n2916), 
	.B2(FE_OFN8_n73), 
	.B1(n188), 
	.A2(n187), 
	.A1(n147));
   INV_X1 U139 (.ZN(n187), 
	.A(\UUT/Mpath/the_mult/x_operand1[26] ));
   OAI21_X1 U140 (.ZN(n2917), 
	.B2(FE_OFN8_n73), 
	.B1(FE_OFN1_n189), 
	.A(n190));
   NAND2_X1 U141 (.ZN(n190), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN120_UUT_Mpath_the_mult_x_operand2_25_));
   OAI22_X1 U142 (.ZN(n2918), 
	.B2(FE_OFN1_n189), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N34 ));
   AOI211_X1 U143 (.ZN(n189), 
	.C2(n108), 
	.C1(n175), 
	.B(n191), 
	.A(n176));
   INV_X1 U144 (.ZN(n191), 
	.A(n192));
   AOI22_X1 U145 (.ZN(n192), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [9]), 
	.B1(n125), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [23]), 
	.A1(n179));
   OAI222_X1 U146 (.ZN(n108), 
	.C2(n132), 
	.C1(n5475), 
	.B2(n131), 
	.B1(n194), 
	.A2(n129), 
	.A1(FE_OFN21_n193));
   OAI221_X1 U147 (.ZN(n2919), 
	.C2(n135), 
	.C1(n5692), 
	.B2(n195), 
	.B1(n133), 
	.A(n196));
   AOI22_X1 U148 (.ZN(n196), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [57]), 
	.A2(n197), 
	.A1(n137));
   OAI221_X1 U149 (.ZN(n2920), 
	.C2(n142), 
	.C1(n5642), 
	.B2(n198), 
	.B1(n140), 
	.A(n199));
   AOI22_X1 U150 (.ZN(n199), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [25]), 
	.A2(n197), 
	.A1(n144));
   INV_X1 U151 (.ZN(n197), 
	.A(n5643));
   OAI22_X1 U152 (.ZN(n2921), 
	.B2(net54875), 
	.B1(n5643), 
	.A2(n200), 
	.A1(net54953));
   OAI22_X1 U153 (.ZN(n2922), 
	.B2(FE_OFN8_n73), 
	.B1(n201), 
	.A2(n200), 
	.A1(n147));
   INV_X1 U154 (.ZN(n200), 
	.A(FE_OFN121_UUT_Mpath_the_mult_x_operand1_25_));
   OAI21_X1 U155 (.ZN(n2923), 
	.B2(FE_OFN8_n73), 
	.B1(FE_OFN3_n202), 
	.A(n203));
   NAND2_X1 U156 (.ZN(n203), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [24]));
   OAI22_X1 U157 (.ZN(n2924), 
	.B2(FE_OFN3_n202), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N36 ));
   AOI211_X1 U158 (.ZN(n202), 
	.C2(n106), 
	.C1(n175), 
	.B(n204), 
	.A(n176));
   INV_X1 U159 (.ZN(n204), 
	.A(n205));
   AOI22_X1 U160 (.ZN(n205), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [8]), 
	.B1(n125), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [22]), 
	.A1(n179));
   NOR2_X1 U161 (.ZN(n179), 
	.A2(n5872), 
	.A1(n206));
   INV_X1 U162 (.ZN(n206), 
	.A(n207));
   OAI222_X1 U163 (.ZN(n106), 
	.C2(n132), 
	.C1(n5478), 
	.B2(n131), 
	.B1(n209), 
	.A2(n129), 
	.A1(FE_OFN192_n208));
   OAI221_X1 U164 (.ZN(n2925), 
	.C2(n135), 
	.C1(n5693), 
	.B2(n210), 
	.B1(n133), 
	.A(n211));
   AOI22_X1 U165 (.ZN(n211), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [56]), 
	.A2(n212), 
	.A1(n137));
   OAI221_X1 U166 (.ZN(n2926), 
	.C2(n142), 
	.C1(n5644), 
	.B2(n213), 
	.B1(n140), 
	.A(n214));
   AOI22_X1 U167 (.ZN(n214), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [24]), 
	.A2(n212), 
	.A1(n144));
   INV_X1 U168 (.ZN(n212), 
	.A(n5645));
   OAI22_X1 U169 (.ZN(n2927), 
	.B2(net54875), 
	.B1(n5645), 
	.A2(n215), 
	.A1(net54953));
   OAI22_X1 U170 (.ZN(n2928), 
	.B2(FE_OFN8_n73), 
	.B1(n216), 
	.A2(n215), 
	.A1(n147));
   INV_X1 U171 (.ZN(n215), 
	.A(\UUT/Mpath/the_mult/x_operand1[24] ));
   OAI22_X1 U172 (.ZN(n2929), 
	.B2(n216), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N35 ));
   INV_X1 U173 (.ZN(n216), 
	.A(n217));
   OAI222_X1 U174 (.ZN(n217), 
	.C2(n5421), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN192_n208), 
	.B1(n5528), 
	.A2(n209), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U175 (.ZN(n2930), 
	.B2(n219), 
	.B1(n209), 
	.A2(n6407), 
	.A1(n5396));
   OAI22_X1 U176 (.ZN(n2931), 
	.B2(n221), 
	.B1(n209), 
	.A2(n6410), 
	.A1(n5364));
   OAI22_X1 U177 (.ZN(n2932), 
	.B2(n223), 
	.B1(n209), 
	.A2(n6401), 
	.A1(n5332));
   OAI22_X1 U178 (.ZN(n2933), 
	.B2(n225), 
	.B1(n209), 
	.A2(n6406), 
	.A1(n5300));
   OAI22_X1 U179 (.ZN(n2934), 
	.B2(n227), 
	.B1(n209), 
	.A2(n6399), 
	.A1(n5268));
   OAI22_X1 U180 (.ZN(n2935), 
	.B2(n229), 
	.B1(n209), 
	.A2(n6404), 
	.A1(n5236));
   OAI22_X1 U181 (.ZN(n2936), 
	.B2(n231), 
	.B1(n209), 
	.A2(n6398), 
	.A1(n5204));
   OAI22_X1 U182 (.ZN(n2937), 
	.B2(n233), 
	.B1(n209), 
	.A2(n6396), 
	.A1(n5172));
   OAI22_X1 U183 (.ZN(n2938), 
	.B2(n235), 
	.B1(n209), 
	.A2(n6393), 
	.A1(n5140));
   OAI22_X1 U184 (.ZN(n2939), 
	.B2(n237), 
	.B1(n209), 
	.A2(n6391), 
	.A1(n5108));
   OAI22_X1 U185 (.ZN(n2940), 
	.B2(n239), 
	.B1(n209), 
	.A2(n6390), 
	.A1(n5076));
   OAI22_X1 U186 (.ZN(n2941), 
	.B2(n241), 
	.B1(n209), 
	.A2(n6388), 
	.A1(n5044));
   OAI22_X1 U187 (.ZN(n2942), 
	.B2(n243), 
	.B1(n209), 
	.A2(n6385), 
	.A1(n5012));
   OAI22_X1 U188 (.ZN(n2943), 
	.B2(n245), 
	.B1(n209), 
	.A2(n6383), 
	.A1(n4980));
   OAI22_X1 U189 (.ZN(n2944), 
	.B2(n247), 
	.B1(n209), 
	.A2(n6382), 
	.A1(n4948));
   OAI22_X1 U190 (.ZN(n2945), 
	.B2(n249), 
	.B1(n209), 
	.A2(n6380), 
	.A1(n4916));
   OAI22_X1 U191 (.ZN(n2946), 
	.B2(n251), 
	.B1(n209), 
	.A2(n6384), 
	.A1(n4884));
   OAI22_X1 U192 (.ZN(n2947), 
	.B2(n253), 
	.B1(n209), 
	.A2(n6381), 
	.A1(n4852));
   OAI22_X1 U193 (.ZN(n2948), 
	.B2(n255), 
	.B1(n209), 
	.A2(n6387), 
	.A1(n4820));
   OAI22_X1 U194 (.ZN(n2949), 
	.B2(n257), 
	.B1(n209), 
	.A2(n6386), 
	.A1(n4788));
   OAI22_X1 U195 (.ZN(n2950), 
	.B2(n259), 
	.B1(n209), 
	.A2(n6392), 
	.A1(n4756));
   OAI22_X1 U196 (.ZN(n2951), 
	.B2(n261), 
	.B1(n209), 
	.A2(n6394), 
	.A1(n4724));
   OAI22_X1 U197 (.ZN(n2952), 
	.B2(n263), 
	.B1(n209), 
	.A2(n6389), 
	.A1(n4692));
   OAI22_X1 U198 (.ZN(n2953), 
	.B2(n265), 
	.B1(n209), 
	.A2(n6395), 
	.A1(n4660));
   OAI22_X1 U199 (.ZN(n2954), 
	.B2(n267), 
	.B1(n209), 
	.A2(n6400), 
	.A1(n4628));
   OAI22_X1 U200 (.ZN(n2955), 
	.B2(n269), 
	.B1(n209), 
	.A2(n6402), 
	.A1(n4596));
   OAI22_X1 U201 (.ZN(n2956), 
	.B2(n271), 
	.B1(n209), 
	.A2(n6397), 
	.A1(n4564));
   OAI22_X1 U202 (.ZN(n2957), 
	.B2(n273), 
	.B1(n209), 
	.A2(n6403), 
	.A1(n4532));
   OAI22_X1 U203 (.ZN(n2958), 
	.B2(n275), 
	.B1(n209), 
	.A2(n6408), 
	.A1(n4500));
   OAI22_X1 U204 (.ZN(n2959), 
	.B2(n277), 
	.B1(n209), 
	.A2(n6405), 
	.A1(n4468));
   OAI22_X1 U205 (.ZN(n2960), 
	.B2(n279), 
	.B1(n209), 
	.A2(n6411), 
	.A1(n4436));
   OAI22_X1 U208 (.ZN(n2961), 
	.B2(FE_OFN192_n208), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5479));
   AOI221_X1 U209 (.ZN(n208), 
	.C2(FE_OFN91_n285), 
	.C1(n5605), 
	.B2(n284), 
	.B1(n283), 
	.A(n286));
   INV_X1 U210 (.ZN(n286), 
	.A(n287));
   AOI222_X1 U211 (.ZN(n287), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[24] ), 
	.B2(n5606), 
	.B1(FE_OFN89_n290), 
	.A2(n289), 
	.A1(n288));
   INV_X1 U212 (.ZN(n289), 
	.A(n5644));
   INV_X1 U213 (.ZN(n283), 
	.A(n5693));
   OAI221_X1 U214 (.ZN(n2962), 
	.C2(n71), 
	.C1(n103), 
	.B2(n69), 
	.B1(FE_OFN101_n292), 
	.A(n293));
   NAND2_X1 U215 (.ZN(n293), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [22]));
   OAI222_X1 U218 (.ZN(n2964), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N40 ), 
	.B2(n300), 
	.B1(FE_OFN101_n292), 
	.A2(n123), 
	.A1(n103));
   INV_X1 U219 (.ZN(n103), 
	.A(n301));
   OAI222_X1 U220 (.ZN(n301), 
	.C2(n132), 
	.C1(n5484), 
	.B2(n131), 
	.B1(n303), 
	.A2(n129), 
	.A1(n302));
   OAI221_X1 U221 (.ZN(n2965), 
	.C2(n135), 
	.C1(n5695), 
	.B2(n304), 
	.B1(n133), 
	.A(n305));
   AOI22_X1 U222 (.ZN(n305), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [54]), 
	.A2(n306), 
	.A1(n137));
   OAI221_X1 U223 (.ZN(n2966), 
	.C2(n142), 
	.C1(n5648), 
	.B2(n307), 
	.B1(n140), 
	.A(n308));
   AOI22_X1 U224 (.ZN(n308), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [22]), 
	.A2(n306), 
	.A1(n144));
   INV_X1 U225 (.ZN(n306), 
	.A(n5649));
   OAI22_X1 U226 (.ZN(n2967), 
	.B2(net54873), 
	.B1(n5649), 
	.A2(n309), 
	.A1(net54953));
   OAI221_X1 U227 (.ZN(n2968), 
	.C2(n309), 
	.C1(n147), 
	.B2(n310), 
	.B1(n302), 
	.A(n311));
   AOI22_X1 U228 (.ZN(n311), 
	.B2(n315), 
	.B1(FE_OFN6_n314), 
	.A2(n313), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U229 (.ZN(n309), 
	.A(\UUT/Mpath/the_mult/x_operand1[22] ));
   OAI221_X1 U230 (.ZN(n2969), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N39 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n302), 
	.A(n317));
   AOI22_X1 U231 (.ZN(n317), 
	.B2(n315), 
	.B1(FE_OFN4_n319), 
	.A2(n313), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U232 (.ZN(n2970), 
	.B2(n219), 
	.B1(n303), 
	.A2(n6407), 
	.A1(n5398));
   OAI22_X1 U233 (.ZN(n2971), 
	.B2(n221), 
	.B1(n303), 
	.A2(n6410), 
	.A1(n5366));
   OAI22_X1 U234 (.ZN(n2972), 
	.B2(n223), 
	.B1(n303), 
	.A2(n6401), 
	.A1(n5334));
   OAI22_X1 U235 (.ZN(n2973), 
	.B2(n225), 
	.B1(n303), 
	.A2(n6406), 
	.A1(n5302));
   OAI22_X1 U236 (.ZN(n2974), 
	.B2(n227), 
	.B1(n303), 
	.A2(n6399), 
	.A1(n5270));
   OAI22_X1 U237 (.ZN(n2975), 
	.B2(n229), 
	.B1(n303), 
	.A2(n6404), 
	.A1(n5238));
   OAI22_X1 U238 (.ZN(n2976), 
	.B2(n231), 
	.B1(n303), 
	.A2(n6398), 
	.A1(n5206));
   OAI22_X1 U239 (.ZN(n2977), 
	.B2(n233), 
	.B1(n303), 
	.A2(n6396), 
	.A1(n5174));
   OAI22_X1 U240 (.ZN(n2978), 
	.B2(n235), 
	.B1(n303), 
	.A2(n6393), 
	.A1(n5142));
   OAI22_X1 U241 (.ZN(n2979), 
	.B2(n237), 
	.B1(n303), 
	.A2(n6391), 
	.A1(n5110));
   OAI22_X1 U242 (.ZN(n2980), 
	.B2(n239), 
	.B1(n303), 
	.A2(n6390), 
	.A1(n5078));
   OAI22_X1 U243 (.ZN(n2981), 
	.B2(n241), 
	.B1(n303), 
	.A2(n6388), 
	.A1(n5046));
   OAI22_X1 U244 (.ZN(n2982), 
	.B2(n243), 
	.B1(n303), 
	.A2(n6385), 
	.A1(n5014));
   OAI22_X1 U245 (.ZN(n2983), 
	.B2(n245), 
	.B1(n303), 
	.A2(n6383), 
	.A1(n4982));
   OAI22_X1 U246 (.ZN(n2984), 
	.B2(n247), 
	.B1(n303), 
	.A2(n6382), 
	.A1(n4950));
   OAI22_X1 U247 (.ZN(n2985), 
	.B2(n249), 
	.B1(n303), 
	.A2(n6380), 
	.A1(n4918));
   OAI22_X1 U248 (.ZN(n2986), 
	.B2(n251), 
	.B1(n303), 
	.A2(n6384), 
	.A1(n4886));
   OAI22_X1 U249 (.ZN(n2987), 
	.B2(n253), 
	.B1(n303), 
	.A2(n6381), 
	.A1(n4854));
   OAI22_X1 U250 (.ZN(n2988), 
	.B2(n255), 
	.B1(n303), 
	.A2(n6387), 
	.A1(n4822));
   OAI22_X1 U251 (.ZN(n2989), 
	.B2(n257), 
	.B1(n303), 
	.A2(n6386), 
	.A1(n4790));
   OAI22_X1 U252 (.ZN(n2990), 
	.B2(n259), 
	.B1(n303), 
	.A2(n6392), 
	.A1(n4758));
   OAI22_X1 U253 (.ZN(n2991), 
	.B2(n261), 
	.B1(n303), 
	.A2(n6394), 
	.A1(n4726));
   OAI22_X1 U254 (.ZN(n2992), 
	.B2(n263), 
	.B1(n303), 
	.A2(n6389), 
	.A1(n4694));
   OAI22_X1 U255 (.ZN(n2993), 
	.B2(n265), 
	.B1(n303), 
	.A2(n6395), 
	.A1(n4662));
   OAI22_X1 U256 (.ZN(n2994), 
	.B2(n267), 
	.B1(n303), 
	.A2(n6400), 
	.A1(n4630));
   OAI22_X1 U257 (.ZN(n2995), 
	.B2(n269), 
	.B1(n303), 
	.A2(n6402), 
	.A1(n4598));
   OAI22_X1 U258 (.ZN(n2996), 
	.B2(n271), 
	.B1(n303), 
	.A2(n6397), 
	.A1(n4566));
   OAI22_X1 U259 (.ZN(n2997), 
	.B2(n273), 
	.B1(n303), 
	.A2(n6403), 
	.A1(n4534));
   OAI22_X1 U260 (.ZN(n2998), 
	.B2(n275), 
	.B1(n303), 
	.A2(n6408), 
	.A1(n4502));
   OAI22_X1 U261 (.ZN(n2999), 
	.B2(n277), 
	.B1(n303), 
	.A2(n6405), 
	.A1(n4470));
   OAI22_X1 U262 (.ZN(n3000), 
	.B2(n279), 
	.B1(n303), 
	.A2(n6411), 
	.A1(n4438));
   OAI221_X1 U264 (.ZN(n315), 
	.C2(n5485), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5772), 
	.A(n282));
   OAI22_X1 U265 (.ZN(n3001), 
	.B2(n302), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5485));
   INV_X1 U266 (.ZN(n302), 
	.A(n320));
   OAI211_X1 U267 (.ZN(n320), 
	.C2(n321), 
	.C1(n5648), 
	.B(n323), 
	.A(n322));
   AOI222_X1 U268 (.ZN(n323), 
	.C2(n326), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[22] ), 
	.A2(n324), 
	.A1(FE_OFN91_n285));
   INV_X1 U269 (.ZN(n326), 
	.A(n5695));
   AOI22_X1 U270 (.ZN(n322), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[22] ), 
	.A2(n6100), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U271 (.ZN(n3002), 
	.C2(n71), 
	.C1(n102), 
	.B2(n69), 
	.B1(FE_OFN100_n327), 
	.A(n328));
   NAND2_X1 U272 (.ZN(n328), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [21]));
   OAI222_X1 U275 (.ZN(n3004), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N42 ), 
	.B2(n300), 
	.B1(FE_OFN100_n327), 
	.A2(n123), 
	.A1(n102));
   INV_X1 U276 (.ZN(n102), 
	.A(n330));
   OAI222_X1 U277 (.ZN(n330), 
	.C2(n132), 
	.C1(n5487), 
	.B2(n131), 
	.B1(n332), 
	.A2(n129), 
	.A1(n331));
   OAI221_X1 U278 (.ZN(n3005), 
	.C2(n135), 
	.C1(n5696), 
	.B2(n333), 
	.B1(n133), 
	.A(n334));
   AOI22_X1 U279 (.ZN(n334), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [53]), 
	.A2(n335), 
	.A1(n137));
   OAI221_X1 U280 (.ZN(n3006), 
	.C2(n142), 
	.C1(n5650), 
	.B2(n336), 
	.B1(n140), 
	.A(n337));
   AOI22_X1 U281 (.ZN(n337), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [21]), 
	.A2(n335), 
	.A1(n144));
   INV_X1 U282 (.ZN(n335), 
	.A(n5651));
   OAI22_X1 U283 (.ZN(n3007), 
	.B2(net54875), 
	.B1(n5651), 
	.A2(n338), 
	.A1(FE_OFN11_net54953));
   OAI221_X1 U284 (.ZN(n3008), 
	.C2(n338), 
	.C1(n147), 
	.B2(n310), 
	.B1(n331), 
	.A(n339));
   AOI22_X1 U285 (.ZN(n339), 
	.B2(n341), 
	.B1(FE_OFN6_n314), 
	.A2(n340), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U286 (.ZN(n338), 
	.A(FE_OFCN204_FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_));
   OAI221_X1 U287 (.ZN(n3009), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N41 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n331), 
	.A(n342));
   AOI22_X1 U288 (.ZN(n342), 
	.B2(n341), 
	.B1(FE_OFN4_n319), 
	.A2(n340), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U289 (.ZN(n3010), 
	.B2(n219), 
	.B1(n332), 
	.A2(n218), 
	.A1(n5399));
   OAI22_X1 U290 (.ZN(n3011), 
	.B2(n221), 
	.B1(n332), 
	.A2(n220), 
	.A1(n5367));
   OAI22_X1 U291 (.ZN(n3012), 
	.B2(n223), 
	.B1(n332), 
	.A2(n222), 
	.A1(n5335));
   OAI22_X1 U292 (.ZN(n3013), 
	.B2(n225), 
	.B1(n332), 
	.A2(n224), 
	.A1(n5303));
   OAI22_X1 U293 (.ZN(n3014), 
	.B2(n227), 
	.B1(n332), 
	.A2(n226), 
	.A1(n5271));
   OAI22_X1 U294 (.ZN(n3015), 
	.B2(n229), 
	.B1(n332), 
	.A2(n228), 
	.A1(n5239));
   OAI22_X1 U295 (.ZN(n3016), 
	.B2(n231), 
	.B1(n332), 
	.A2(n230), 
	.A1(n5207));
   OAI22_X1 U296 (.ZN(n3017), 
	.B2(n233), 
	.B1(n332), 
	.A2(n232), 
	.A1(n5175));
   OAI22_X1 U297 (.ZN(n3018), 
	.B2(n235), 
	.B1(n332), 
	.A2(n234), 
	.A1(n5143));
   OAI22_X1 U298 (.ZN(n3019), 
	.B2(n237), 
	.B1(n332), 
	.A2(n236), 
	.A1(n5111));
   OAI22_X1 U299 (.ZN(n3020), 
	.B2(n239), 
	.B1(n332), 
	.A2(n238), 
	.A1(n5079));
   OAI22_X1 U300 (.ZN(n3021), 
	.B2(n241), 
	.B1(n332), 
	.A2(n240), 
	.A1(n5047));
   OAI22_X1 U301 (.ZN(n3022), 
	.B2(n243), 
	.B1(n332), 
	.A2(n242), 
	.A1(n5015));
   OAI22_X1 U302 (.ZN(n3023), 
	.B2(n245), 
	.B1(n332), 
	.A2(n244), 
	.A1(n4983));
   OAI22_X1 U303 (.ZN(n3024), 
	.B2(n247), 
	.B1(n332), 
	.A2(n246), 
	.A1(n4951));
   OAI22_X1 U304 (.ZN(n3025), 
	.B2(n249), 
	.B1(n332), 
	.A2(n248), 
	.A1(n4919));
   OAI22_X1 U305 (.ZN(n3026), 
	.B2(n251), 
	.B1(n332), 
	.A2(n250), 
	.A1(n4887));
   OAI22_X1 U306 (.ZN(n3027), 
	.B2(n253), 
	.B1(n332), 
	.A2(n252), 
	.A1(n4855));
   OAI22_X1 U307 (.ZN(n3028), 
	.B2(n255), 
	.B1(n332), 
	.A2(n254), 
	.A1(n4823));
   OAI22_X1 U308 (.ZN(n3029), 
	.B2(n257), 
	.B1(n332), 
	.A2(n256), 
	.A1(n4791));
   OAI22_X1 U309 (.ZN(n3030), 
	.B2(n259), 
	.B1(n332), 
	.A2(n258), 
	.A1(n4759));
   OAI22_X1 U310 (.ZN(n3031), 
	.B2(n261), 
	.B1(n332), 
	.A2(n260), 
	.A1(n4727));
   OAI22_X1 U311 (.ZN(n3032), 
	.B2(n263), 
	.B1(n332), 
	.A2(n262), 
	.A1(n4695));
   OAI22_X1 U312 (.ZN(n3033), 
	.B2(n265), 
	.B1(n332), 
	.A2(n264), 
	.A1(n4663));
   OAI22_X1 U313 (.ZN(n3034), 
	.B2(n267), 
	.B1(n332), 
	.A2(n266), 
	.A1(n4631));
   OAI22_X1 U314 (.ZN(n3035), 
	.B2(n269), 
	.B1(n332), 
	.A2(n268), 
	.A1(n4599));
   OAI22_X1 U315 (.ZN(n3036), 
	.B2(n271), 
	.B1(n332), 
	.A2(n270), 
	.A1(n4567));
   OAI22_X1 U316 (.ZN(n3037), 
	.B2(n273), 
	.B1(n332), 
	.A2(n272), 
	.A1(n4535));
   OAI22_X1 U317 (.ZN(n3038), 
	.B2(n275), 
	.B1(n332), 
	.A2(n274), 
	.A1(n4503));
   OAI22_X1 U318 (.ZN(n3039), 
	.B2(n277), 
	.B1(n332), 
	.A2(n276), 
	.A1(n4471));
   OAI22_X1 U319 (.ZN(n3040), 
	.B2(n279), 
	.B1(n332), 
	.A2(n278), 
	.A1(n4439));
   OAI221_X1 U321 (.ZN(n341), 
	.C2(n5488), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5789), 
	.A(n282));
   OAI22_X1 U322 (.ZN(n3041), 
	.B2(n331), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5488));
   INV_X1 U323 (.ZN(n331), 
	.A(n343));
   OAI211_X1 U324 (.ZN(n343), 
	.C2(n321), 
	.C1(n5650), 
	.B(n345), 
	.A(n344));
   AOI222_X1 U325 (.ZN(n345), 
	.C2(n347), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[21] ), 
	.A2(n346), 
	.A1(FE_OFN91_n285));
   INV_X1 U326 (.ZN(n347), 
	.A(n5696));
   AOI22_X1 U327 (.ZN(n344), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[21] ), 
	.A2(n6107), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U328 (.ZN(n3042), 
	.C2(n71), 
	.C1(n101), 
	.B2(n69), 
	.B1(FE_OFN99_n348), 
	.A(n349));
   NAND2_X1 U329 (.ZN(n349), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [20]));
   OAI222_X1 U332 (.ZN(n3044), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N44 ), 
	.B2(n300), 
	.B1(FE_OFN99_n348), 
	.A2(n123), 
	.A1(n101));
   INV_X1 U333 (.ZN(n101), 
	.A(n351));
   OAI222_X1 U334 (.ZN(n351), 
	.C2(n132), 
	.C1(n5490), 
	.B2(n131), 
	.B1(n353), 
	.A2(n129), 
	.A1(n352));
   OAI221_X1 U335 (.ZN(n3045), 
	.C2(n135), 
	.C1(n5697), 
	.B2(n354), 
	.B1(n133), 
	.A(n355));
   AOI22_X1 U336 (.ZN(n355), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [52]), 
	.A2(n356), 
	.A1(n137));
   OAI221_X1 U337 (.ZN(n3046), 
	.C2(n142), 
	.C1(n5652), 
	.B2(n357), 
	.B1(n140), 
	.A(n358));
   AOI22_X1 U338 (.ZN(n358), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [20]), 
	.A2(n356), 
	.A1(n144));
   INV_X1 U339 (.ZN(n356), 
	.A(n5653));
   OAI22_X1 U340 (.ZN(n3047), 
	.B2(net54873), 
	.B1(n5653), 
	.A2(n359), 
	.A1(net54953));
   OAI221_X1 U341 (.ZN(n3048), 
	.C2(n359), 
	.C1(n147), 
	.B2(n310), 
	.B1(n352), 
	.A(n360));
   AOI22_X1 U342 (.ZN(n360), 
	.B2(n362), 
	.B1(FE_OFN6_n314), 
	.A2(n361), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U343 (.ZN(n359), 
	.A(\UUT/Mpath/the_mult/x_operand1[20] ));
   OAI221_X1 U344 (.ZN(n3049), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N43 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n352), 
	.A(n363));
   AOI22_X1 U345 (.ZN(n363), 
	.B2(n362), 
	.B1(FE_OFN4_n319), 
	.A2(n361), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U346 (.ZN(n3050), 
	.B2(n219), 
	.B1(n353), 
	.A2(n6407), 
	.A1(n5400));
   OAI22_X1 U347 (.ZN(n3051), 
	.B2(n221), 
	.B1(n353), 
	.A2(n6410), 
	.A1(n5368));
   OAI22_X1 U348 (.ZN(n3052), 
	.B2(n223), 
	.B1(n353), 
	.A2(n6401), 
	.A1(n5336));
   OAI22_X1 U349 (.ZN(n3053), 
	.B2(n225), 
	.B1(n353), 
	.A2(n6406), 
	.A1(n5304));
   OAI22_X1 U350 (.ZN(n3054), 
	.B2(n227), 
	.B1(n353), 
	.A2(n6399), 
	.A1(n5272));
   OAI22_X1 U351 (.ZN(n3055), 
	.B2(n229), 
	.B1(n353), 
	.A2(n6404), 
	.A1(n5240));
   OAI22_X1 U352 (.ZN(n3056), 
	.B2(n231), 
	.B1(n353), 
	.A2(n6398), 
	.A1(n5208));
   OAI22_X1 U353 (.ZN(n3057), 
	.B2(n233), 
	.B1(n353), 
	.A2(n6396), 
	.A1(n5176));
   OAI22_X1 U354 (.ZN(n3058), 
	.B2(n235), 
	.B1(n353), 
	.A2(n6393), 
	.A1(n5144));
   OAI22_X1 U355 (.ZN(n3059), 
	.B2(n237), 
	.B1(n353), 
	.A2(n6391), 
	.A1(n5112));
   OAI22_X1 U356 (.ZN(n3060), 
	.B2(n239), 
	.B1(n353), 
	.A2(n6390), 
	.A1(n5080));
   OAI22_X1 U357 (.ZN(n3061), 
	.B2(n241), 
	.B1(n353), 
	.A2(n6388), 
	.A1(n5048));
   OAI22_X1 U358 (.ZN(n3062), 
	.B2(n243), 
	.B1(n353), 
	.A2(n6385), 
	.A1(n5016));
   OAI22_X1 U359 (.ZN(n3063), 
	.B2(n245), 
	.B1(n353), 
	.A2(n6383), 
	.A1(n4984));
   OAI22_X1 U360 (.ZN(n3064), 
	.B2(n247), 
	.B1(n353), 
	.A2(n6382), 
	.A1(n4952));
   OAI22_X1 U361 (.ZN(n3065), 
	.B2(n249), 
	.B1(n353), 
	.A2(n6380), 
	.A1(n4920));
   OAI22_X1 U362 (.ZN(n3066), 
	.B2(n251), 
	.B1(n353), 
	.A2(n6384), 
	.A1(n4888));
   OAI22_X1 U363 (.ZN(n3067), 
	.B2(n253), 
	.B1(n353), 
	.A2(n6381), 
	.A1(n4856));
   OAI22_X1 U364 (.ZN(n3068), 
	.B2(n255), 
	.B1(n353), 
	.A2(n6387), 
	.A1(n4824));
   OAI22_X1 U365 (.ZN(n3069), 
	.B2(n257), 
	.B1(n353), 
	.A2(n6386), 
	.A1(n4792));
   OAI22_X1 U366 (.ZN(n3070), 
	.B2(n259), 
	.B1(n353), 
	.A2(n6392), 
	.A1(n4760));
   OAI22_X1 U367 (.ZN(n3071), 
	.B2(n261), 
	.B1(n353), 
	.A2(n6394), 
	.A1(n4728));
   OAI22_X1 U368 (.ZN(n3072), 
	.B2(n263), 
	.B1(n353), 
	.A2(n6389), 
	.A1(n4696));
   OAI22_X1 U369 (.ZN(n3073), 
	.B2(n265), 
	.B1(n353), 
	.A2(n6395), 
	.A1(n4664));
   OAI22_X1 U370 (.ZN(n3074), 
	.B2(n267), 
	.B1(n353), 
	.A2(n6400), 
	.A1(n4632));
   OAI22_X1 U371 (.ZN(n3075), 
	.B2(n269), 
	.B1(n353), 
	.A2(n6402), 
	.A1(n4600));
   OAI22_X1 U372 (.ZN(n3076), 
	.B2(n271), 
	.B1(n353), 
	.A2(n6397), 
	.A1(n4568));
   OAI22_X1 U373 (.ZN(n3077), 
	.B2(n273), 
	.B1(n353), 
	.A2(n6403), 
	.A1(n4536));
   OAI22_X1 U374 (.ZN(n3078), 
	.B2(n275), 
	.B1(n353), 
	.A2(n6408), 
	.A1(n4504));
   OAI22_X1 U375 (.ZN(n3079), 
	.B2(n277), 
	.B1(n353), 
	.A2(n6405), 
	.A1(n4472));
   OAI22_X1 U376 (.ZN(n3080), 
	.B2(n279), 
	.B1(n353), 
	.A2(n6411), 
	.A1(n4440));
   OAI221_X1 U378 (.ZN(n362), 
	.C2(n5491), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5802), 
	.A(n282));
   OAI22_X1 U379 (.ZN(n3081), 
	.B2(n352), 
	.B1(FE_OFN11_net54953), 
	.A2(net54883), 
	.A1(n5491));
   INV_X1 U380 (.ZN(n352), 
	.A(n364));
   OAI211_X1 U381 (.ZN(n364), 
	.C2(n321), 
	.C1(n5652), 
	.B(n366), 
	.A(n365));
   AOI222_X1 U382 (.ZN(n366), 
	.C2(n368), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[20] ), 
	.A2(n367), 
	.A1(FE_OFN91_n285));
   INV_X1 U383 (.ZN(n368), 
	.A(n5697));
   AOI22_X1 U384 (.ZN(n365), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[20] ), 
	.A2(n6114), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U385 (.ZN(n3082), 
	.C2(n71), 
	.C1(n100), 
	.B2(n69), 
	.B1(n369), 
	.A(n370));
   NAND2_X1 U386 (.ZN(n370), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN129_UUT_Mpath_the_mult_x_operand2_19_));
   INV_X1 U387 (.ZN(n100), 
	.A(n371));
   INV_X1 U390 (.ZN(n369), 
	.A(\UUT/break_code[19] ));
   OAI211_X1 U391 (.ZN(n3084), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N46 ), 
	.B(n374), 
	.A(n373));
   AOI222_X1 U392 (.ZN(n374), 
	.C2(n6126), 
	.C1(n377), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [3]), 
	.B1(n376), 
	.A2(n371), 
	.A1(n375));
   OAI222_X1 U393 (.ZN(n371), 
	.C2(n132), 
	.C1(n5496), 
	.B2(n131), 
	.B1(n379), 
	.A2(n129), 
	.A1(n378));
   OAI221_X1 U394 (.ZN(n3085), 
	.C2(n135), 
	.C1(n5699), 
	.B2(n380), 
	.B1(n133), 
	.A(n381));
   AOI22_X1 U395 (.ZN(n381), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [51]), 
	.A2(n382), 
	.A1(n137));
   OAI221_X1 U396 (.ZN(n3086), 
	.C2(n142), 
	.C1(n5656), 
	.B2(n383), 
	.B1(n140), 
	.A(n384));
   AOI22_X1 U397 (.ZN(n384), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [19]), 
	.A2(n382), 
	.A1(n144));
   INV_X1 U398 (.ZN(n382), 
	.A(n5657));
   OAI22_X1 U399 (.ZN(n3087), 
	.B2(net54873), 
	.B1(n5657), 
	.A2(n385), 
	.A1(net54953));
   OAI221_X1 U400 (.ZN(n3088), 
	.C2(n385), 
	.C1(n147), 
	.B2(n310), 
	.B1(n378), 
	.A(n386));
   AOI22_X1 U401 (.ZN(n386), 
	.B2(n388), 
	.B1(FE_OFN6_n314), 
	.A2(n387), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U402 (.ZN(n385), 
	.A(FE_OFN130_UUT_Mpath_the_mult_x_operand1_19_));
   OAI221_X1 U403 (.ZN(n3089), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N45 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n378), 
	.A(n389));
   AOI22_X1 U404 (.ZN(n389), 
	.B2(n388), 
	.B1(FE_OFN4_n319), 
	.A2(n387), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U405 (.ZN(n3090), 
	.B2(n219), 
	.B1(n379), 
	.A2(n218), 
	.A1(n5402));
   OAI22_X1 U406 (.ZN(n3091), 
	.B2(n221), 
	.B1(n379), 
	.A2(n220), 
	.A1(n5370));
   OAI22_X1 U407 (.ZN(n3092), 
	.B2(n223), 
	.B1(n379), 
	.A2(n222), 
	.A1(n5338));
   OAI22_X1 U408 (.ZN(n3093), 
	.B2(n225), 
	.B1(n379), 
	.A2(n224), 
	.A1(n5306));
   OAI22_X1 U409 (.ZN(n3094), 
	.B2(n227), 
	.B1(n379), 
	.A2(n226), 
	.A1(n5274));
   OAI22_X1 U410 (.ZN(n3095), 
	.B2(n229), 
	.B1(n379), 
	.A2(n228), 
	.A1(n5242));
   OAI22_X1 U411 (.ZN(n3096), 
	.B2(n231), 
	.B1(n379), 
	.A2(n230), 
	.A1(n5210));
   OAI22_X1 U412 (.ZN(n3097), 
	.B2(n233), 
	.B1(n379), 
	.A2(n232), 
	.A1(n5178));
   OAI22_X1 U413 (.ZN(n3098), 
	.B2(n235), 
	.B1(n379), 
	.A2(n234), 
	.A1(n5146));
   OAI22_X1 U414 (.ZN(n3099), 
	.B2(n237), 
	.B1(n379), 
	.A2(n236), 
	.A1(n5114));
   OAI22_X1 U415 (.ZN(n3100), 
	.B2(n239), 
	.B1(n379), 
	.A2(n238), 
	.A1(n5082));
   OAI22_X1 U416 (.ZN(n3101), 
	.B2(n241), 
	.B1(n379), 
	.A2(n240), 
	.A1(n5050));
   OAI22_X1 U417 (.ZN(n3102), 
	.B2(n243), 
	.B1(n379), 
	.A2(n242), 
	.A1(n5018));
   OAI22_X1 U418 (.ZN(n3103), 
	.B2(n245), 
	.B1(n379), 
	.A2(n244), 
	.A1(n4986));
   OAI22_X1 U419 (.ZN(n3104), 
	.B2(n247), 
	.B1(n379), 
	.A2(n246), 
	.A1(n4954));
   OAI22_X1 U420 (.ZN(n3105), 
	.B2(n249), 
	.B1(n379), 
	.A2(n248), 
	.A1(n4922));
   OAI22_X1 U421 (.ZN(n3106), 
	.B2(n251), 
	.B1(n379), 
	.A2(n250), 
	.A1(n4890));
   OAI22_X1 U422 (.ZN(n3107), 
	.B2(n253), 
	.B1(n379), 
	.A2(n252), 
	.A1(n4858));
   OAI22_X1 U423 (.ZN(n3108), 
	.B2(n255), 
	.B1(n379), 
	.A2(n254), 
	.A1(n4826));
   OAI22_X1 U424 (.ZN(n3109), 
	.B2(n257), 
	.B1(n379), 
	.A2(n256), 
	.A1(n4794));
   OAI22_X1 U425 (.ZN(n3110), 
	.B2(n259), 
	.B1(n379), 
	.A2(n258), 
	.A1(n4762));
   OAI22_X1 U426 (.ZN(n3111), 
	.B2(n261), 
	.B1(n379), 
	.A2(n260), 
	.A1(n4730));
   OAI22_X1 U427 (.ZN(n3112), 
	.B2(n263), 
	.B1(n379), 
	.A2(n262), 
	.A1(n4698));
   OAI22_X1 U428 (.ZN(n3113), 
	.B2(n265), 
	.B1(n379), 
	.A2(n264), 
	.A1(n4666));
   OAI22_X1 U429 (.ZN(n3114), 
	.B2(n267), 
	.B1(n379), 
	.A2(n266), 
	.A1(n4634));
   OAI22_X1 U430 (.ZN(n3115), 
	.B2(n269), 
	.B1(n379), 
	.A2(n268), 
	.A1(n4602));
   OAI22_X1 U431 (.ZN(n3116), 
	.B2(n271), 
	.B1(n379), 
	.A2(n270), 
	.A1(n4570));
   OAI22_X1 U432 (.ZN(n3117), 
	.B2(n273), 
	.B1(n379), 
	.A2(n272), 
	.A1(n4538));
   OAI22_X1 U433 (.ZN(n3118), 
	.B2(n275), 
	.B1(n379), 
	.A2(n274), 
	.A1(n4506));
   OAI22_X1 U434 (.ZN(n3119), 
	.B2(n277), 
	.B1(n379), 
	.A2(n276), 
	.A1(n4474));
   OAI22_X1 U435 (.ZN(n3120), 
	.B2(n279), 
	.B1(n379), 
	.A2(n278), 
	.A1(n4442));
   OAI221_X1 U437 (.ZN(n388), 
	.C2(n5497), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5815), 
	.A(n282));
   OAI22_X1 U438 (.ZN(n3121), 
	.B2(n378), 
	.B1(FE_OFN11_net54953), 
	.A2(net54883), 
	.A1(n5497));
   INV_X1 U439 (.ZN(n378), 
	.A(n390));
   OAI211_X1 U440 (.ZN(n390), 
	.C2(n321), 
	.C1(n5656), 
	.B(n392), 
	.A(n391));
   AOI222_X1 U441 (.ZN(n392), 
	.C2(n394), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[19] ), 
	.A2(n393), 
	.A1(FE_OFN91_n285));
   INV_X1 U442 (.ZN(n394), 
	.A(n5699));
   AOI22_X1 U443 (.ZN(n391), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[19] ), 
	.A2(n6124), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U444 (.ZN(n3122), 
	.C2(n71), 
	.C1(n99), 
	.B2(n69), 
	.B1(n395), 
	.A(n396));
   NAND2_X1 U445 (.ZN(n396), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [18]));
   INV_X1 U446 (.ZN(n99), 
	.A(n397));
   INV_X1 U449 (.ZN(n395), 
	.A(\UUT/break_code[18] ));
   OAI211_X1 U450 (.ZN(n3124), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N48 ), 
	.B(n399), 
	.A(n373));
   AOI222_X1 U451 (.ZN(n399), 
	.C2(n377), 
	.C1(n6135), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [2]), 
	.B1(n376), 
	.A2(n397), 
	.A1(n375));
   OAI222_X1 U452 (.ZN(n397), 
	.C2(n132), 
	.C1(n5499), 
	.B2(n131), 
	.B1(n401), 
	.A2(n129), 
	.A1(n400));
   OAI221_X1 U453 (.ZN(n3125), 
	.C2(n135), 
	.C1(n5700), 
	.B2(n402), 
	.B1(n133), 
	.A(n403));
   AOI22_X1 U454 (.ZN(n403), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [50]), 
	.A2(n404), 
	.A1(n137));
   OAI221_X1 U455 (.ZN(n3126), 
	.C2(n142), 
	.C1(n5658), 
	.B2(n405), 
	.B1(n140), 
	.A(n406));
   AOI22_X1 U456 (.ZN(n406), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [18]), 
	.A2(n404), 
	.A1(n144));
   INV_X1 U457 (.ZN(n404), 
	.A(n5659));
   OAI22_X1 U458 (.ZN(n3127), 
	.B2(net54873), 
	.B1(n5659), 
	.A2(n407), 
	.A1(FE_OFN10_net54953));
   OAI221_X1 U459 (.ZN(n3128), 
	.C2(n407), 
	.C1(n147), 
	.B2(n310), 
	.B1(n400), 
	.A(n408));
   AOI22_X1 U460 (.ZN(n408), 
	.B2(n410), 
	.B1(FE_OFN6_n314), 
	.A2(n409), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U461 (.ZN(n407), 
	.A(\UUT/Mpath/the_mult/x_operand1[18] ));
   OAI221_X1 U462 (.ZN(n3129), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N47 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n400), 
	.A(n411));
   AOI22_X1 U463 (.ZN(n411), 
	.B2(n410), 
	.B1(FE_OFN4_n319), 
	.A2(n409), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U464 (.ZN(n3130), 
	.B2(n219), 
	.B1(n401), 
	.A2(n6407), 
	.A1(n5403));
   OAI22_X1 U465 (.ZN(n3131), 
	.B2(n221), 
	.B1(n401), 
	.A2(n6410), 
	.A1(n5371));
   OAI22_X1 U466 (.ZN(n3132), 
	.B2(n223), 
	.B1(n401), 
	.A2(n6401), 
	.A1(n5339));
   OAI22_X1 U467 (.ZN(n3133), 
	.B2(n225), 
	.B1(n401), 
	.A2(n6406), 
	.A1(n5307));
   OAI22_X1 U468 (.ZN(n3134), 
	.B2(n227), 
	.B1(n401), 
	.A2(n6399), 
	.A1(n5275));
   OAI22_X1 U469 (.ZN(n3135), 
	.B2(n229), 
	.B1(n401), 
	.A2(n6404), 
	.A1(n5243));
   OAI22_X1 U470 (.ZN(n3136), 
	.B2(n231), 
	.B1(n401), 
	.A2(n6398), 
	.A1(n5211));
   OAI22_X1 U471 (.ZN(n3137), 
	.B2(n233), 
	.B1(n401), 
	.A2(n6396), 
	.A1(n5179));
   OAI22_X1 U472 (.ZN(n3138), 
	.B2(n235), 
	.B1(n401), 
	.A2(n6393), 
	.A1(n5147));
   OAI22_X1 U473 (.ZN(n3139), 
	.B2(n237), 
	.B1(n401), 
	.A2(n6391), 
	.A1(n5115));
   OAI22_X1 U474 (.ZN(n3140), 
	.B2(n239), 
	.B1(n401), 
	.A2(n6390), 
	.A1(n5083));
   OAI22_X1 U475 (.ZN(n3141), 
	.B2(n241), 
	.B1(n401), 
	.A2(n6388), 
	.A1(n5051));
   OAI22_X1 U476 (.ZN(n3142), 
	.B2(n243), 
	.B1(n401), 
	.A2(n6385), 
	.A1(n5019));
   OAI22_X1 U477 (.ZN(n3143), 
	.B2(n245), 
	.B1(n401), 
	.A2(n6383), 
	.A1(n4987));
   OAI22_X1 U478 (.ZN(n3144), 
	.B2(n247), 
	.B1(n401), 
	.A2(n6382), 
	.A1(n4955));
   OAI22_X1 U479 (.ZN(n3145), 
	.B2(n249), 
	.B1(n401), 
	.A2(n6380), 
	.A1(n4923));
   OAI22_X1 U480 (.ZN(n3146), 
	.B2(n251), 
	.B1(n401), 
	.A2(n6384), 
	.A1(n4891));
   OAI22_X1 U481 (.ZN(n3147), 
	.B2(n253), 
	.B1(n401), 
	.A2(n6381), 
	.A1(n4859));
   OAI22_X1 U482 (.ZN(n3148), 
	.B2(n255), 
	.B1(n401), 
	.A2(n6387), 
	.A1(n4827));
   OAI22_X1 U483 (.ZN(n3149), 
	.B2(n257), 
	.B1(n401), 
	.A2(n6386), 
	.A1(n4795));
   OAI22_X1 U484 (.ZN(n3150), 
	.B2(n259), 
	.B1(n401), 
	.A2(n6392), 
	.A1(n4763));
   OAI22_X1 U485 (.ZN(n3151), 
	.B2(n261), 
	.B1(n401), 
	.A2(n6394), 
	.A1(n4731));
   OAI22_X1 U486 (.ZN(n3152), 
	.B2(n263), 
	.B1(n401), 
	.A2(n6389), 
	.A1(n4699));
   OAI22_X1 U487 (.ZN(n3153), 
	.B2(n265), 
	.B1(n401), 
	.A2(n6395), 
	.A1(n4667));
   OAI22_X1 U488 (.ZN(n3154), 
	.B2(n267), 
	.B1(n401), 
	.A2(n6400), 
	.A1(n4635));
   OAI22_X1 U489 (.ZN(n3155), 
	.B2(n269), 
	.B1(n401), 
	.A2(n6402), 
	.A1(n4603));
   OAI22_X1 U490 (.ZN(n3156), 
	.B2(n271), 
	.B1(n401), 
	.A2(n6397), 
	.A1(n4571));
   OAI22_X1 U491 (.ZN(n3157), 
	.B2(n273), 
	.B1(n401), 
	.A2(n6403), 
	.A1(n4539));
   OAI22_X1 U492 (.ZN(n3158), 
	.B2(n275), 
	.B1(n401), 
	.A2(n6408), 
	.A1(n4507));
   OAI22_X1 U493 (.ZN(n3159), 
	.B2(n277), 
	.B1(n401), 
	.A2(n6405), 
	.A1(n4475));
   OAI22_X1 U494 (.ZN(n3160), 
	.B2(n279), 
	.B1(n401), 
	.A2(n6411), 
	.A1(n4443));
   OAI221_X1 U496 (.ZN(n410), 
	.C2(n5500), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5841), 
	.A(n282));
   OAI22_X1 U497 (.ZN(n3161), 
	.B2(n400), 
	.B1(FE_OFN11_net54953), 
	.A2(net54883), 
	.A1(n5500));
   INV_X1 U498 (.ZN(n400), 
	.A(n412));
   OAI211_X1 U499 (.ZN(n412), 
	.C2(n321), 
	.C1(n5658), 
	.B(n414), 
	.A(n413));
   AOI222_X1 U500 (.ZN(n414), 
	.C2(n416), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[18] ), 
	.A2(n415), 
	.A1(FE_OFN91_n285));
   INV_X1 U501 (.ZN(n416), 
	.A(n5700));
   AOI22_X1 U502 (.ZN(n413), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[18] ), 
	.A2(n6134), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U503 (.ZN(n3162), 
	.C2(n71), 
	.C1(n98), 
	.B2(n69), 
	.B1(n417), 
	.A(n418));
   NAND2_X1 U504 (.ZN(n418), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN133_UUT_Mpath_the_mult_x_operand2_17_));
   INV_X1 U505 (.ZN(n98), 
	.A(n419));
   INV_X1 U508 (.ZN(n417), 
	.A(\UUT/break_code[17] ));
   OAI211_X1 U509 (.ZN(n3164), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N50 ), 
	.B(n421), 
	.A(n373));
   AOI222_X1 U510 (.ZN(n421), 
	.C2(n377), 
	.C1(n6153), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [1]), 
	.B1(n376), 
	.A2(n419), 
	.A1(n375));
   OAI222_X1 U511 (.ZN(n419), 
	.C2(n132), 
	.C1(n5502), 
	.B2(n131), 
	.B1(n423), 
	.A2(n129), 
	.A1(n422));
   OAI221_X1 U512 (.ZN(n3165), 
	.C2(n135), 
	.C1(n5701), 
	.B2(n424), 
	.B1(n133), 
	.A(n425));
   AOI22_X1 U513 (.ZN(n425), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [49]), 
	.A2(n426), 
	.A1(n137));
   OAI221_X1 U514 (.ZN(n3166), 
	.C2(n142), 
	.C1(n5660), 
	.B2(n427), 
	.B1(n140), 
	.A(n428));
   AOI22_X1 U515 (.ZN(n428), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [17]), 
	.A2(n426), 
	.A1(n144));
   INV_X1 U516 (.ZN(n426), 
	.A(n5661));
   OAI22_X1 U517 (.ZN(n3167), 
	.B2(net54873), 
	.B1(n5661), 
	.A2(n429), 
	.A1(FE_OFN10_net54953));
   OAI221_X1 U518 (.ZN(n3168), 
	.C2(n429), 
	.C1(n147), 
	.B2(n310), 
	.B1(n422), 
	.A(n430));
   AOI22_X1 U519 (.ZN(n430), 
	.B2(n432), 
	.B1(FE_OFN6_n314), 
	.A2(n431), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U520 (.ZN(n429), 
	.A(FE_OFN134_UUT_Mpath_the_mult_x_operand1_17_));
   OAI221_X1 U521 (.ZN(n3169), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N49 ), 
	.B2(n316), 
	.B1(n422), 
	.A(n433));
   AOI22_X1 U522 (.ZN(n433), 
	.B2(n432), 
	.B1(FE_OFN4_n319), 
	.A2(n431), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U523 (.ZN(n3170), 
	.B2(n219), 
	.B1(n423), 
	.A2(n6407), 
	.A1(n5404));
   OAI22_X1 U524 (.ZN(n3171), 
	.B2(n221), 
	.B1(n423), 
	.A2(n6410), 
	.A1(n5372));
   OAI22_X1 U525 (.ZN(n3172), 
	.B2(n223), 
	.B1(n423), 
	.A2(n6401), 
	.A1(n5340));
   OAI22_X1 U526 (.ZN(n3173), 
	.B2(n225), 
	.B1(n423), 
	.A2(n6406), 
	.A1(n5308));
   OAI22_X1 U527 (.ZN(n3174), 
	.B2(n227), 
	.B1(n423), 
	.A2(n6399), 
	.A1(n5276));
   OAI22_X1 U528 (.ZN(n3175), 
	.B2(n229), 
	.B1(n423), 
	.A2(n6404), 
	.A1(n5244));
   OAI22_X1 U529 (.ZN(n3176), 
	.B2(n231), 
	.B1(n423), 
	.A2(n6398), 
	.A1(n5212));
   OAI22_X1 U530 (.ZN(n3177), 
	.B2(n233), 
	.B1(n423), 
	.A2(n6396), 
	.A1(n5180));
   OAI22_X1 U531 (.ZN(n3178), 
	.B2(n235), 
	.B1(n423), 
	.A2(n6393), 
	.A1(n5148));
   OAI22_X1 U532 (.ZN(n3179), 
	.B2(n237), 
	.B1(n423), 
	.A2(n6391), 
	.A1(n5116));
   OAI22_X1 U533 (.ZN(n3180), 
	.B2(n239), 
	.B1(n423), 
	.A2(n6390), 
	.A1(n5084));
   OAI22_X1 U534 (.ZN(n3181), 
	.B2(n241), 
	.B1(n423), 
	.A2(n6388), 
	.A1(n5052));
   OAI22_X1 U535 (.ZN(n3182), 
	.B2(n243), 
	.B1(n423), 
	.A2(n6385), 
	.A1(n5020));
   OAI22_X1 U536 (.ZN(n3183), 
	.B2(n245), 
	.B1(n423), 
	.A2(n6383), 
	.A1(n4988));
   OAI22_X1 U537 (.ZN(n3184), 
	.B2(n247), 
	.B1(n423), 
	.A2(n6382), 
	.A1(n4956));
   OAI22_X1 U538 (.ZN(n3185), 
	.B2(n249), 
	.B1(n423), 
	.A2(n6380), 
	.A1(n4924));
   OAI22_X1 U539 (.ZN(n3186), 
	.B2(n251), 
	.B1(n423), 
	.A2(n6384), 
	.A1(n4892));
   OAI22_X1 U540 (.ZN(n3187), 
	.B2(n253), 
	.B1(n423), 
	.A2(n6381), 
	.A1(n4860));
   OAI22_X1 U541 (.ZN(n3188), 
	.B2(n255), 
	.B1(n423), 
	.A2(n6387), 
	.A1(n4828));
   OAI22_X1 U542 (.ZN(n3189), 
	.B2(n257), 
	.B1(n423), 
	.A2(n6386), 
	.A1(n4796));
   OAI22_X1 U543 (.ZN(n3190), 
	.B2(n259), 
	.B1(n423), 
	.A2(n6392), 
	.A1(n4764));
   OAI22_X1 U544 (.ZN(n3191), 
	.B2(n261), 
	.B1(n423), 
	.A2(n6394), 
	.A1(n4732));
   OAI22_X1 U545 (.ZN(n3192), 
	.B2(n263), 
	.B1(n423), 
	.A2(n6389), 
	.A1(n4700));
   OAI22_X1 U546 (.ZN(n3193), 
	.B2(n265), 
	.B1(n423), 
	.A2(n6395), 
	.A1(n4668));
   OAI22_X1 U547 (.ZN(n3194), 
	.B2(n267), 
	.B1(n423), 
	.A2(n6400), 
	.A1(n4636));
   OAI22_X1 U548 (.ZN(n3195), 
	.B2(n269), 
	.B1(n423), 
	.A2(n6402), 
	.A1(n4604));
   OAI22_X1 U549 (.ZN(n3196), 
	.B2(n271), 
	.B1(n423), 
	.A2(n6397), 
	.A1(n4572));
   OAI22_X1 U550 (.ZN(n3197), 
	.B2(n273), 
	.B1(n423), 
	.A2(n6403), 
	.A1(n4540));
   OAI22_X1 U551 (.ZN(n3198), 
	.B2(n275), 
	.B1(n423), 
	.A2(n6408), 
	.A1(n4508));
   OAI22_X1 U552 (.ZN(n3199), 
	.B2(n277), 
	.B1(n423), 
	.A2(n6405), 
	.A1(n4476));
   OAI22_X1 U553 (.ZN(n3200), 
	.B2(n279), 
	.B1(n423), 
	.A2(n6411), 
	.A1(n4444));
   OAI221_X1 U555 (.ZN(n432), 
	.C2(n5503), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5919), 
	.A(n282));
   OAI22_X1 U556 (.ZN(n3201), 
	.B2(n422), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5503));
   INV_X1 U557 (.ZN(n422), 
	.A(n434));
   OAI211_X1 U558 (.ZN(n434), 
	.C2(n321), 
	.C1(n5660), 
	.B(n436), 
	.A(n435));
   AOI222_X1 U559 (.ZN(n436), 
	.C2(n438), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[17] ), 
	.A2(n437), 
	.A1(FE_OFN91_n285));
   INV_X1 U560 (.ZN(n438), 
	.A(n5701));
   AOI22_X1 U561 (.ZN(n435), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[17] ), 
	.A2(n6152), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U562 (.ZN(n3202), 
	.C2(n71), 
	.C1(n97), 
	.B2(n69), 
	.B1(n439), 
	.A(n440));
   NAND2_X1 U563 (.ZN(n440), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN136_UUT_Mpath_the_mult_x_operand2_16_));
   INV_X1 U564 (.ZN(n97), 
	.A(n441));
   INV_X1 U567 (.ZN(n439), 
	.A(\UUT/break_code[16] ));
   OAI211_X1 U568 (.ZN(n3204), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N52 ), 
	.B(n443), 
	.A(n373));
   AOI222_X1 U569 (.ZN(n443), 
	.C2(n377), 
	.C1(n6162), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [0]), 
	.B1(n376), 
	.A2(n441), 
	.A1(n375));
   AND2_X1 U570 (.ZN(n377), 
	.A2(n445), 
	.A1(n444));
   AND2_X1 U571 (.ZN(n376), 
	.A2(net54895), 
	.A1(n125));
   OAI222_X1 U572 (.ZN(n441), 
	.C2(n132), 
	.C1(n5505), 
	.B2(n131), 
	.B1(n447), 
	.A2(n129), 
	.A1(n446));
   INV_X1 U573 (.ZN(n375), 
	.A(n123));
   AOI22_X1 U574 (.ZN(n373), 
	.B2(n444), 
	.B1(n6127), 
	.A2(n449), 
	.A1(n448));
   NOR3_X1 U575 (.ZN(n444), 
	.A3(n450), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U576 (.ZN(n3205), 
	.C2(n135), 
	.C1(n5702), 
	.B2(n451), 
	.B1(n133), 
	.A(n452));
   AOI22_X1 U577 (.ZN(n452), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [48]), 
	.A2(n453), 
	.A1(n137));
   OAI221_X1 U578 (.ZN(n3206), 
	.C2(n142), 
	.C1(n5662), 
	.B2(n454), 
	.B1(n140), 
	.A(n455));
   AOI22_X1 U579 (.ZN(n455), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [16]), 
	.A2(n453), 
	.A1(n144));
   INV_X1 U580 (.ZN(n453), 
	.A(n5663));
   OAI22_X1 U581 (.ZN(n3207), 
	.B2(net54873), 
	.B1(n5663), 
	.A2(n456), 
	.A1(net54953));
   OAI221_X1 U582 (.ZN(n3208), 
	.C2(n456), 
	.C1(n147), 
	.B2(n310), 
	.B1(n446), 
	.A(n457));
   AOI22_X1 U583 (.ZN(n457), 
	.B2(n459), 
	.B1(FE_OFN6_n314), 
	.A2(n458), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U584 (.ZN(n456), 
	.A(\UUT/Mpath/the_mult/x_operand1[16] ));
   OAI221_X1 U585 (.ZN(n3209), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N51 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n446), 
	.A(n460));
   AOI22_X1 U586 (.ZN(n460), 
	.B2(n459), 
	.B1(FE_OFN4_n319), 
	.A2(n458), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U587 (.ZN(n3210), 
	.B2(n219), 
	.B1(n447), 
	.A2(n6407), 
	.A1(n5405));
   OAI22_X1 U588 (.ZN(n3211), 
	.B2(n221), 
	.B1(n447), 
	.A2(n6410), 
	.A1(n5373));
   OAI22_X1 U589 (.ZN(n3212), 
	.B2(n223), 
	.B1(n447), 
	.A2(n6401), 
	.A1(n5341));
   OAI22_X1 U590 (.ZN(n3213), 
	.B2(n225), 
	.B1(n447), 
	.A2(n6406), 
	.A1(n5309));
   OAI22_X1 U591 (.ZN(n3214), 
	.B2(n227), 
	.B1(n447), 
	.A2(n6399), 
	.A1(n5277));
   OAI22_X1 U592 (.ZN(n3215), 
	.B2(n229), 
	.B1(n447), 
	.A2(n6404), 
	.A1(n5245));
   OAI22_X1 U593 (.ZN(n3216), 
	.B2(n231), 
	.B1(n447), 
	.A2(n6398), 
	.A1(n5213));
   OAI22_X1 U594 (.ZN(n3217), 
	.B2(n233), 
	.B1(n447), 
	.A2(n6396), 
	.A1(n5181));
   OAI22_X1 U595 (.ZN(n3218), 
	.B2(n235), 
	.B1(n447), 
	.A2(n6393), 
	.A1(n5149));
   OAI22_X1 U596 (.ZN(n3219), 
	.B2(n237), 
	.B1(n447), 
	.A2(n6391), 
	.A1(n5117));
   OAI22_X1 U597 (.ZN(n3220), 
	.B2(n239), 
	.B1(n447), 
	.A2(n6390), 
	.A1(n5085));
   OAI22_X1 U598 (.ZN(n3221), 
	.B2(n241), 
	.B1(n447), 
	.A2(n6388), 
	.A1(n5053));
   OAI22_X1 U599 (.ZN(n3222), 
	.B2(n243), 
	.B1(n447), 
	.A2(n6385), 
	.A1(n5021));
   OAI22_X1 U600 (.ZN(n3223), 
	.B2(n245), 
	.B1(n447), 
	.A2(n6383), 
	.A1(n4989));
   OAI22_X1 U601 (.ZN(n3224), 
	.B2(n247), 
	.B1(n447), 
	.A2(n6382), 
	.A1(n4957));
   OAI22_X1 U602 (.ZN(n3225), 
	.B2(n249), 
	.B1(n447), 
	.A2(n6380), 
	.A1(n4925));
   OAI22_X1 U603 (.ZN(n3226), 
	.B2(n251), 
	.B1(n447), 
	.A2(n6384), 
	.A1(n4893));
   OAI22_X1 U604 (.ZN(n3227), 
	.B2(n253), 
	.B1(n447), 
	.A2(n6381), 
	.A1(n4861));
   OAI22_X1 U605 (.ZN(n3228), 
	.B2(n255), 
	.B1(n447), 
	.A2(n6387), 
	.A1(n4829));
   OAI22_X1 U606 (.ZN(n3229), 
	.B2(n257), 
	.B1(n447), 
	.A2(n6386), 
	.A1(n4797));
   OAI22_X1 U607 (.ZN(n3230), 
	.B2(n259), 
	.B1(n447), 
	.A2(n6392), 
	.A1(n4765));
   OAI22_X1 U608 (.ZN(n3231), 
	.B2(n261), 
	.B1(n447), 
	.A2(n6394), 
	.A1(n4733));
   OAI22_X1 U609 (.ZN(n3232), 
	.B2(n263), 
	.B1(n447), 
	.A2(n6389), 
	.A1(n4701));
   OAI22_X1 U610 (.ZN(n3233), 
	.B2(n265), 
	.B1(n447), 
	.A2(n6395), 
	.A1(n4669));
   OAI22_X1 U611 (.ZN(n3234), 
	.B2(n267), 
	.B1(n447), 
	.A2(n6400), 
	.A1(n4637));
   OAI22_X1 U612 (.ZN(n3235), 
	.B2(n269), 
	.B1(n447), 
	.A2(n6402), 
	.A1(n4605));
   OAI22_X1 U613 (.ZN(n3236), 
	.B2(n271), 
	.B1(n447), 
	.A2(n6397), 
	.A1(n4573));
   OAI22_X1 U614 (.ZN(n3237), 
	.B2(n273), 
	.B1(n447), 
	.A2(n6403), 
	.A1(n4541));
   OAI22_X1 U615 (.ZN(n3238), 
	.B2(n275), 
	.B1(n447), 
	.A2(n6408), 
	.A1(n4509));
   OAI22_X1 U616 (.ZN(n3239), 
	.B2(n277), 
	.B1(n447), 
	.A2(n6405), 
	.A1(n4477));
   OAI22_X1 U617 (.ZN(n3240), 
	.B2(n279), 
	.B1(n447), 
	.A2(n6411), 
	.A1(n4445));
   OAI221_X1 U619 (.ZN(n459), 
	.C2(n5506), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5944), 
	.A(n282));
   OAI22_X1 U620 (.ZN(n3241), 
	.B2(n446), 
	.B1(FE_OFN11_net54953), 
	.A2(net54885), 
	.A1(n5506));
   INV_X1 U621 (.ZN(n446), 
	.A(n461));
   OAI211_X1 U622 (.ZN(n461), 
	.C2(n321), 
	.C1(n5662), 
	.B(n463), 
	.A(n462));
   AOI222_X1 U623 (.ZN(n463), 
	.C2(n465), 
	.C1(n284), 
	.B2(n325), 
	.B1(\UUT/Mpath/out_jar[16] ), 
	.A2(n464), 
	.A1(FE_OFN91_n285));
   INV_X1 U624 (.ZN(n465), 
	.A(n5702));
   AOI22_X1 U625 (.ZN(n462), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[16] ), 
	.A2(n6161), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U626 (.ZN(n3242), 
	.C2(n71), 
	.C1(n96), 
	.B2(n466), 
	.B1(n69), 
	.A(n467));
   NAND2_X1 U627 (.ZN(n467), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN137_UUT_Mpath_the_mult_x_operand2_15_));
   OAI222_X1 U630 (.ZN(n3244), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N54 ), 
	.B2(n466), 
	.B1(n300), 
	.A2(n123), 
	.A1(n96));
   INV_X1 U631 (.ZN(n96), 
	.A(n469));
   OAI222_X1 U632 (.ZN(n469), 
	.C2(n132), 
	.C1(n5508), 
	.B2(n131), 
	.B1(n471), 
	.A2(n129), 
	.A1(n470));
   OAI221_X1 U633 (.ZN(n3245), 
	.C2(n135), 
	.C1(n5703), 
	.B2(n472), 
	.B1(n133), 
	.A(n473));
   AOI22_X1 U634 (.ZN(n473), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [47]), 
	.A2(n474), 
	.A1(n137));
   OAI221_X1 U635 (.ZN(n3246), 
	.C2(n142), 
	.C1(n5664), 
	.B2(n475), 
	.B1(n140), 
	.A(n476));
   AOI22_X1 U636 (.ZN(n476), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [15]), 
	.A2(n474), 
	.A1(n144));
   INV_X1 U637 (.ZN(n474), 
	.A(n5665));
   OAI22_X1 U638 (.ZN(n3247), 
	.B2(net54873), 
	.B1(n5665), 
	.A2(n477), 
	.A1(net54953));
   OAI221_X1 U639 (.ZN(n3248), 
	.C2(n477), 
	.C1(n147), 
	.B2(n310), 
	.B1(n470), 
	.A(n478));
   AOI22_X1 U640 (.ZN(n478), 
	.B2(n480), 
	.B1(FE_OFN6_n314), 
	.A2(n479), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U641 (.ZN(n477), 
	.A(FE_OFN138_UUT_Mpath_the_mult_x_operand1_15_));
   OAI221_X1 U642 (.ZN(n3249), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N53 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n470), 
	.A(n481));
   AOI22_X1 U643 (.ZN(n481), 
	.B2(n480), 
	.B1(FE_OFN4_n319), 
	.A2(n479), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U644 (.ZN(n3250), 
	.B2(n219), 
	.B1(n471), 
	.A2(n6407), 
	.A1(n5406));
   OAI22_X1 U645 (.ZN(n3251), 
	.B2(n221), 
	.B1(n471), 
	.A2(n6410), 
	.A1(n5374));
   OAI22_X1 U646 (.ZN(n3252), 
	.B2(n223), 
	.B1(n471), 
	.A2(n6401), 
	.A1(n5342));
   OAI22_X1 U647 (.ZN(n3253), 
	.B2(n225), 
	.B1(n471), 
	.A2(n6406), 
	.A1(n5310));
   OAI22_X1 U648 (.ZN(n3254), 
	.B2(n227), 
	.B1(n471), 
	.A2(n6399), 
	.A1(n5278));
   OAI22_X1 U649 (.ZN(n3255), 
	.B2(n229), 
	.B1(n471), 
	.A2(n6404), 
	.A1(n5246));
   OAI22_X1 U650 (.ZN(n3256), 
	.B2(n231), 
	.B1(n471), 
	.A2(n6398), 
	.A1(n5214));
   OAI22_X1 U651 (.ZN(n3257), 
	.B2(n233), 
	.B1(n471), 
	.A2(n6396), 
	.A1(n5182));
   OAI22_X1 U652 (.ZN(n3258), 
	.B2(n235), 
	.B1(n471), 
	.A2(n6393), 
	.A1(n5150));
   OAI22_X1 U653 (.ZN(n3259), 
	.B2(n237), 
	.B1(n471), 
	.A2(n6391), 
	.A1(n5118));
   OAI22_X1 U654 (.ZN(n3260), 
	.B2(n239), 
	.B1(n471), 
	.A2(n6390), 
	.A1(n5086));
   OAI22_X1 U655 (.ZN(n3261), 
	.B2(n241), 
	.B1(n471), 
	.A2(n6388), 
	.A1(n5054));
   OAI22_X1 U656 (.ZN(n3262), 
	.B2(n243), 
	.B1(n471), 
	.A2(n6385), 
	.A1(n5022));
   OAI22_X1 U657 (.ZN(n3263), 
	.B2(n245), 
	.B1(n471), 
	.A2(n6383), 
	.A1(n4990));
   OAI22_X1 U658 (.ZN(n3264), 
	.B2(n247), 
	.B1(n471), 
	.A2(n6382), 
	.A1(n4958));
   OAI22_X1 U659 (.ZN(n3265), 
	.B2(n249), 
	.B1(n471), 
	.A2(n6380), 
	.A1(n4926));
   OAI22_X1 U660 (.ZN(n3266), 
	.B2(n251), 
	.B1(n471), 
	.A2(n6384), 
	.A1(n4894));
   OAI22_X1 U661 (.ZN(n3267), 
	.B2(n253), 
	.B1(n471), 
	.A2(n6381), 
	.A1(n4862));
   OAI22_X1 U662 (.ZN(n3268), 
	.B2(n255), 
	.B1(n471), 
	.A2(n6387), 
	.A1(n4830));
   OAI22_X1 U663 (.ZN(n3269), 
	.B2(n257), 
	.B1(n471), 
	.A2(n6386), 
	.A1(n4798));
   OAI22_X1 U664 (.ZN(n3270), 
	.B2(n259), 
	.B1(n471), 
	.A2(n6392), 
	.A1(n4766));
   OAI22_X1 U665 (.ZN(n3271), 
	.B2(n261), 
	.B1(n471), 
	.A2(n6394), 
	.A1(n4734));
   OAI22_X1 U666 (.ZN(n3272), 
	.B2(n263), 
	.B1(n471), 
	.A2(n6389), 
	.A1(n4702));
   OAI22_X1 U667 (.ZN(n3273), 
	.B2(n265), 
	.B1(n471), 
	.A2(n6395), 
	.A1(n4670));
   OAI22_X1 U668 (.ZN(n3274), 
	.B2(n267), 
	.B1(n471), 
	.A2(n6400), 
	.A1(n4638));
   OAI22_X1 U669 (.ZN(n3275), 
	.B2(n269), 
	.B1(n471), 
	.A2(n6402), 
	.A1(n4606));
   OAI22_X1 U670 (.ZN(n3276), 
	.B2(n271), 
	.B1(n471), 
	.A2(n6397), 
	.A1(n4574));
   OAI22_X1 U671 (.ZN(n3277), 
	.B2(n273), 
	.B1(n471), 
	.A2(n6403), 
	.A1(n4542));
   OAI22_X1 U672 (.ZN(n3278), 
	.B2(n275), 
	.B1(n471), 
	.A2(n6408), 
	.A1(n4510));
   OAI22_X1 U673 (.ZN(n3279), 
	.B2(n277), 
	.B1(n471), 
	.A2(n6405), 
	.A1(n4478));
   OAI22_X1 U674 (.ZN(n3280), 
	.B2(n279), 
	.B1(n471), 
	.A2(n6411), 
	.A1(n4446));
   OAI211_X1 U676 (.ZN(n480), 
	.C2(n483), 
	.C1(n482), 
	.B(n485), 
	.A(n484));
   AOI22_X1 U677 (.ZN(n485), 
	.B2(n489), 
	.B1(n488), 
	.A2(n487), 
	.A1(n486));
   INV_X1 U678 (.ZN(n488), 
	.A(n5509));
   INV_X1 U679 (.ZN(n483), 
	.A(n5756));
   OAI22_X1 U680 (.ZN(n3281), 
	.B2(n470), 
	.B1(FE_OFN11_net54953), 
	.A2(net54883), 
	.A1(n5509));
   INV_X1 U681 (.ZN(n470), 
	.A(n490));
   OAI211_X1 U682 (.ZN(n490), 
	.C2(n321), 
	.C1(n5664), 
	.B(n492), 
	.A(n491));
   AOI222_X1 U683 (.ZN(n492), 
	.C2(n494), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[15] ), 
	.A2(n493), 
	.A1(FE_OFN91_n285));
   INV_X1 U684 (.ZN(n494), 
	.A(n5703));
   AOI22_X1 U685 (.ZN(n491), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[15] ), 
	.A2(n6169), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U686 (.ZN(n3282), 
	.C2(n71), 
	.C1(n95), 
	.B2(n69), 
	.B1(n495), 
	.A(n496));
   NAND2_X1 U687 (.ZN(n496), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN140_UUT_Mpath_the_mult_x_operand2_14_));
   OAI222_X1 U690 (.ZN(n3284), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N56 ), 
	.B2(n300), 
	.B1(n495), 
	.A2(n123), 
	.A1(n95));
   INV_X1 U691 (.ZN(n495), 
	.A(\UUT/break_code[14] ));
   INV_X1 U692 (.ZN(n95), 
	.A(n498));
   OAI222_X1 U693 (.ZN(n498), 
	.C2(n132), 
	.C1(n5511), 
	.B2(n131), 
	.B1(n500), 
	.A2(n129), 
	.A1(n499));
   OAI221_X1 U694 (.ZN(n3285), 
	.C2(n135), 
	.C1(n5704), 
	.B2(n501), 
	.B1(n133), 
	.A(n502));
   AOI22_X1 U695 (.ZN(n502), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [46]), 
	.A2(n503), 
	.A1(n137));
   OAI221_X1 U696 (.ZN(n3286), 
	.C2(n142), 
	.C1(n5666), 
	.B2(n504), 
	.B1(n140), 
	.A(n505));
   AOI22_X1 U697 (.ZN(n505), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [14]), 
	.A2(n503), 
	.A1(n144));
   INV_X1 U698 (.ZN(n503), 
	.A(n5667));
   OAI22_X1 U699 (.ZN(n3287), 
	.B2(net54873), 
	.B1(n5667), 
	.A2(n506), 
	.A1(net54953));
   OAI221_X1 U700 (.ZN(n3288), 
	.C2(n506), 
	.C1(n147), 
	.B2(n310), 
	.B1(n499), 
	.A(n507));
   AOI22_X1 U701 (.ZN(n507), 
	.B2(n509), 
	.B1(FE_OFN6_n314), 
	.A2(n508), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U702 (.ZN(n506), 
	.A(\UUT/Mpath/the_mult/x_operand1[14] ));
   OAI221_X1 U703 (.ZN(n3289), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N55 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n499), 
	.A(n510));
   AOI22_X1 U704 (.ZN(n510), 
	.B2(n509), 
	.B1(FE_OFN4_n319), 
	.A2(n508), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U705 (.ZN(n3290), 
	.B2(n219), 
	.B1(n500), 
	.A2(n6407), 
	.A1(n5407));
   OAI22_X1 U706 (.ZN(n3291), 
	.B2(n221), 
	.B1(n500), 
	.A2(n6410), 
	.A1(n5375));
   OAI22_X1 U707 (.ZN(n3292), 
	.B2(n223), 
	.B1(n500), 
	.A2(n6401), 
	.A1(n5343));
   OAI22_X1 U708 (.ZN(n3293), 
	.B2(n225), 
	.B1(n500), 
	.A2(n6406), 
	.A1(n5311));
   OAI22_X1 U709 (.ZN(n3294), 
	.B2(n227), 
	.B1(n500), 
	.A2(n6399), 
	.A1(n5279));
   OAI22_X1 U710 (.ZN(n3295), 
	.B2(n229), 
	.B1(n500), 
	.A2(n6404), 
	.A1(n5247));
   OAI22_X1 U711 (.ZN(n3296), 
	.B2(n231), 
	.B1(n500), 
	.A2(n6398), 
	.A1(n5215));
   OAI22_X1 U712 (.ZN(n3297), 
	.B2(n233), 
	.B1(n500), 
	.A2(n6396), 
	.A1(n5183));
   OAI22_X1 U713 (.ZN(n3298), 
	.B2(n235), 
	.B1(n500), 
	.A2(n6393), 
	.A1(n5151));
   OAI22_X1 U714 (.ZN(n3299), 
	.B2(n237), 
	.B1(n500), 
	.A2(n6391), 
	.A1(n5119));
   OAI22_X1 U715 (.ZN(n3300), 
	.B2(n239), 
	.B1(n500), 
	.A2(n6390), 
	.A1(n5087));
   OAI22_X1 U716 (.ZN(n3301), 
	.B2(n241), 
	.B1(n500), 
	.A2(n6388), 
	.A1(n5055));
   OAI22_X1 U717 (.ZN(n3302), 
	.B2(n243), 
	.B1(n500), 
	.A2(n6385), 
	.A1(n5023));
   OAI22_X1 U718 (.ZN(n3303), 
	.B2(n245), 
	.B1(n500), 
	.A2(n6383), 
	.A1(n4991));
   OAI22_X1 U719 (.ZN(n3304), 
	.B2(n247), 
	.B1(n500), 
	.A2(n6382), 
	.A1(n4959));
   OAI22_X1 U720 (.ZN(n3305), 
	.B2(n249), 
	.B1(n500), 
	.A2(n6380), 
	.A1(n4927));
   OAI22_X1 U721 (.ZN(n3306), 
	.B2(n251), 
	.B1(n500), 
	.A2(n6384), 
	.A1(n4895));
   OAI22_X1 U722 (.ZN(n3307), 
	.B2(n253), 
	.B1(n500), 
	.A2(n6381), 
	.A1(n4863));
   OAI22_X1 U723 (.ZN(n3308), 
	.B2(n255), 
	.B1(n500), 
	.A2(n6387), 
	.A1(n4831));
   OAI22_X1 U724 (.ZN(n3309), 
	.B2(n257), 
	.B1(n500), 
	.A2(n6386), 
	.A1(n4799));
   OAI22_X1 U725 (.ZN(n3310), 
	.B2(n259), 
	.B1(n500), 
	.A2(n6392), 
	.A1(n4767));
   OAI22_X1 U726 (.ZN(n3311), 
	.B2(n261), 
	.B1(n500), 
	.A2(n6394), 
	.A1(n4735));
   OAI22_X1 U727 (.ZN(n3312), 
	.B2(n263), 
	.B1(n500), 
	.A2(n6389), 
	.A1(n4703));
   OAI22_X1 U728 (.ZN(n3313), 
	.B2(n265), 
	.B1(n500), 
	.A2(n6395), 
	.A1(n4671));
   OAI22_X1 U729 (.ZN(n3314), 
	.B2(n267), 
	.B1(n500), 
	.A2(n6400), 
	.A1(n4639));
   OAI22_X1 U730 (.ZN(n3315), 
	.B2(n269), 
	.B1(n500), 
	.A2(n6402), 
	.A1(n4607));
   OAI22_X1 U731 (.ZN(n3316), 
	.B2(n271), 
	.B1(n500), 
	.A2(n6397), 
	.A1(n4575));
   OAI22_X1 U732 (.ZN(n3317), 
	.B2(n273), 
	.B1(n500), 
	.A2(n6403), 
	.A1(n4543));
   OAI22_X1 U733 (.ZN(n3318), 
	.B2(n275), 
	.B1(n500), 
	.A2(n6408), 
	.A1(n4511));
   OAI22_X1 U734 (.ZN(n3319), 
	.B2(n277), 
	.B1(n500), 
	.A2(n6405), 
	.A1(n4479));
   OAI22_X1 U735 (.ZN(n3320), 
	.B2(n279), 
	.B1(n500), 
	.A2(n6411), 
	.A1(n4447));
   OAI211_X1 U737 (.ZN(n509), 
	.C2(n511), 
	.C1(n482), 
	.B(n512), 
	.A(n484));
   AOI22_X1 U738 (.ZN(n512), 
	.B2(n489), 
	.B1(n514), 
	.A2(n513), 
	.A1(n486));
   INV_X1 U739 (.ZN(n514), 
	.A(n5512));
   INV_X1 U740 (.ZN(n511), 
	.A(n5769));
   OAI22_X1 U741 (.ZN(n3321), 
	.B2(n499), 
	.B1(FE_OFN12_net54953), 
	.A2(net54881), 
	.A1(n5512));
   INV_X1 U742 (.ZN(n499), 
	.A(n515));
   OAI211_X1 U743 (.ZN(n515), 
	.C2(n321), 
	.C1(n5666), 
	.B(n517), 
	.A(n516));
   AOI222_X1 U744 (.ZN(n517), 
	.C2(n519), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[14] ), 
	.A2(n518), 
	.A1(FE_OFN91_n285));
   INV_X1 U745 (.ZN(n519), 
	.A(n5704));
   AOI22_X1 U746 (.ZN(n516), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[14] ), 
	.A2(n6180), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U747 (.ZN(n3322), 
	.C2(n71), 
	.C1(n94), 
	.B2(n69), 
	.B1(n520), 
	.A(n521));
   NAND2_X1 U748 (.ZN(n521), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [13]));
   OAI222_X1 U751 (.ZN(n3324), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N58 ), 
	.B2(n300), 
	.B1(n520), 
	.A2(n123), 
	.A1(n94));
   INV_X1 U752 (.ZN(n520), 
	.A(\UUT/break_code[13] ));
   INV_X1 U753 (.ZN(n94), 
	.A(n523));
   OAI222_X1 U754 (.ZN(n523), 
	.C2(n132), 
	.C1(n5514), 
	.B2(n131), 
	.B1(n525), 
	.A2(n129), 
	.A1(n524));
   OAI221_X1 U755 (.ZN(n3325), 
	.C2(n135), 
	.C1(n5705), 
	.B2(n526), 
	.B1(n133), 
	.A(n527));
   AOI22_X1 U756 (.ZN(n527), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [45]), 
	.A2(n528), 
	.A1(n137));
   OAI221_X1 U757 (.ZN(n3326), 
	.C2(n142), 
	.C1(n5668), 
	.B2(n529), 
	.B1(n140), 
	.A(n530));
   AOI22_X1 U758 (.ZN(n530), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [13]), 
	.A2(n528), 
	.A1(n144));
   INV_X1 U759 (.ZN(n528), 
	.A(n5669));
   OAI22_X1 U760 (.ZN(n3327), 
	.B2(net54871), 
	.B1(n5669), 
	.A2(n531), 
	.A1(net54953));
   OAI221_X1 U761 (.ZN(n3328), 
	.C2(n531), 
	.C1(n147), 
	.B2(n310), 
	.B1(n524), 
	.A(n532));
   AOI22_X1 U762 (.ZN(n532), 
	.B2(n534), 
	.B1(FE_OFN6_n314), 
	.A2(n533), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U763 (.ZN(n531), 
	.A(FE_OFN142_UUT_Mpath_the_mult_x_operand1_13_));
   OAI221_X1 U764 (.ZN(n3329), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N57 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n524), 
	.A(n535));
   AOI22_X1 U765 (.ZN(n535), 
	.B2(n534), 
	.B1(FE_OFN4_n319), 
	.A2(n533), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U766 (.ZN(n3330), 
	.B2(n219), 
	.B1(n525), 
	.A2(n6407), 
	.A1(n5408));
   OAI22_X1 U767 (.ZN(n3331), 
	.B2(n221), 
	.B1(n525), 
	.A2(n6410), 
	.A1(n5376));
   OAI22_X1 U768 (.ZN(n3332), 
	.B2(n223), 
	.B1(n525), 
	.A2(n6401), 
	.A1(n5344));
   OAI22_X1 U769 (.ZN(n3333), 
	.B2(n225), 
	.B1(n525), 
	.A2(n6406), 
	.A1(n5312));
   OAI22_X1 U770 (.ZN(n3334), 
	.B2(n227), 
	.B1(n525), 
	.A2(n6399), 
	.A1(n5280));
   OAI22_X1 U771 (.ZN(n3335), 
	.B2(n229), 
	.B1(n525), 
	.A2(n6404), 
	.A1(n5248));
   OAI22_X1 U772 (.ZN(n3336), 
	.B2(n231), 
	.B1(n525), 
	.A2(n6398), 
	.A1(n5216));
   OAI22_X1 U773 (.ZN(n3337), 
	.B2(n233), 
	.B1(n525), 
	.A2(n6396), 
	.A1(n5184));
   OAI22_X1 U774 (.ZN(n3338), 
	.B2(n235), 
	.B1(n525), 
	.A2(n6393), 
	.A1(n5152));
   OAI22_X1 U775 (.ZN(n3339), 
	.B2(n237), 
	.B1(n525), 
	.A2(n6391), 
	.A1(n5120));
   OAI22_X1 U776 (.ZN(n3340), 
	.B2(n239), 
	.B1(n525), 
	.A2(n6390), 
	.A1(n5088));
   OAI22_X1 U777 (.ZN(n3341), 
	.B2(n241), 
	.B1(n525), 
	.A2(n6388), 
	.A1(n5056));
   OAI22_X1 U778 (.ZN(n3342), 
	.B2(n243), 
	.B1(n525), 
	.A2(n6385), 
	.A1(n5024));
   OAI22_X1 U779 (.ZN(n3343), 
	.B2(n245), 
	.B1(n525), 
	.A2(n6383), 
	.A1(n4992));
   OAI22_X1 U780 (.ZN(n3344), 
	.B2(n247), 
	.B1(n525), 
	.A2(n6382), 
	.A1(n4960));
   OAI22_X1 U781 (.ZN(n3345), 
	.B2(n249), 
	.B1(n525), 
	.A2(n6380), 
	.A1(n4928));
   OAI22_X1 U782 (.ZN(n3346), 
	.B2(n251), 
	.B1(n525), 
	.A2(n6384), 
	.A1(n4896));
   OAI22_X1 U783 (.ZN(n3347), 
	.B2(n253), 
	.B1(n525), 
	.A2(n6381), 
	.A1(n4864));
   OAI22_X1 U784 (.ZN(n3348), 
	.B2(n255), 
	.B1(n525), 
	.A2(n6387), 
	.A1(n4832));
   OAI22_X1 U785 (.ZN(n3349), 
	.B2(n257), 
	.B1(n525), 
	.A2(n6386), 
	.A1(n4800));
   OAI22_X1 U786 (.ZN(n3350), 
	.B2(n259), 
	.B1(n525), 
	.A2(n6392), 
	.A1(n4768));
   OAI22_X1 U787 (.ZN(n3351), 
	.B2(n261), 
	.B1(n525), 
	.A2(n6394), 
	.A1(n4736));
   OAI22_X1 U788 (.ZN(n3352), 
	.B2(n263), 
	.B1(n525), 
	.A2(n6389), 
	.A1(n4704));
   OAI22_X1 U789 (.ZN(n3353), 
	.B2(n265), 
	.B1(n525), 
	.A2(n6395), 
	.A1(n4672));
   OAI22_X1 U790 (.ZN(n3354), 
	.B2(n267), 
	.B1(n525), 
	.A2(n6400), 
	.A1(n4640));
   OAI22_X1 U791 (.ZN(n3355), 
	.B2(n269), 
	.B1(n525), 
	.A2(n6402), 
	.A1(n4608));
   OAI22_X1 U792 (.ZN(n3356), 
	.B2(n271), 
	.B1(n525), 
	.A2(n6397), 
	.A1(n4576));
   OAI22_X1 U793 (.ZN(n3357), 
	.B2(n273), 
	.B1(n525), 
	.A2(n6403), 
	.A1(n4544));
   OAI22_X1 U794 (.ZN(n3358), 
	.B2(n275), 
	.B1(n525), 
	.A2(n6408), 
	.A1(n4512));
   OAI22_X1 U795 (.ZN(n3359), 
	.B2(n277), 
	.B1(n525), 
	.A2(n6405), 
	.A1(n4480));
   OAI22_X1 U796 (.ZN(n3360), 
	.B2(n279), 
	.B1(n525), 
	.A2(n6411), 
	.A1(n4448));
   OAI211_X1 U798 (.ZN(n534), 
	.C2(n536), 
	.C1(n482), 
	.B(n537), 
	.A(n484));
   AOI22_X1 U799 (.ZN(n537), 
	.B2(n489), 
	.B1(n539), 
	.A2(n538), 
	.A1(n486));
   INV_X1 U800 (.ZN(n539), 
	.A(n5515));
   INV_X1 U801 (.ZN(n536), 
	.A(n5786));
   OAI22_X1 U802 (.ZN(n3361), 
	.B2(n524), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5515));
   INV_X1 U803 (.ZN(n524), 
	.A(n540));
   OAI211_X1 U804 (.ZN(n540), 
	.C2(n321), 
	.C1(n5668), 
	.B(n542), 
	.A(n541));
   AOI222_X1 U805 (.ZN(n542), 
	.C2(n544), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[13] ), 
	.A2(n543), 
	.A1(FE_OFN91_n285));
   INV_X1 U806 (.ZN(n544), 
	.A(n5705));
   AOI22_X1 U807 (.ZN(n541), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[13] ), 
	.A2(n6187), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U808 (.ZN(n3362), 
	.B2(n2668), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n545));
   OAI221_X1 U809 (.ZN(n3363), 
	.C2(n71), 
	.C1(n93), 
	.B2(n69), 
	.B1(n547), 
	.A(n548));
   NAND2_X1 U810 (.ZN(n548), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [12]));
   OAI222_X1 U811 (.ZN(n3364), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N60 ), 
	.B2(n300), 
	.B1(n547), 
	.A2(n123), 
	.A1(n93));
   INV_X1 U812 (.ZN(n547), 
	.A(\UUT/break_code[12] ));
   INV_X1 U813 (.ZN(n93), 
	.A(n549));
   OAI222_X1 U814 (.ZN(n549), 
	.C2(n132), 
	.C1(n5517), 
	.B2(n131), 
	.B1(n551), 
	.A2(n129), 
	.A1(n550));
   OAI221_X1 U815 (.ZN(n3365), 
	.C2(n135), 
	.C1(n5706), 
	.B2(n552), 
	.B1(n133), 
	.A(n553));
   AOI22_X1 U816 (.ZN(n553), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [44]), 
	.A2(n554), 
	.A1(n137));
   OAI221_X1 U817 (.ZN(n3366), 
	.C2(n142), 
	.C1(n5670), 
	.B2(n555), 
	.B1(n140), 
	.A(n556));
   AOI22_X1 U818 (.ZN(n556), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [12]), 
	.A2(n554), 
	.A1(n144));
   INV_X1 U819 (.ZN(n554), 
	.A(n5671));
   OAI22_X1 U820 (.ZN(n3367), 
	.B2(net54871), 
	.B1(n5671), 
	.A2(n557), 
	.A1(net54953));
   OAI221_X1 U821 (.ZN(n3368), 
	.C2(n557), 
	.C1(n147), 
	.B2(n310), 
	.B1(n550), 
	.A(n558));
   AOI22_X1 U822 (.ZN(n558), 
	.B2(n560), 
	.B1(FE_OFN6_n314), 
	.A2(n559), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U823 (.ZN(n557), 
	.A(\UUT/Mpath/the_mult/x_operand1[12] ));
   OAI221_X1 U824 (.ZN(n3369), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N59 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n550), 
	.A(n561));
   AOI22_X1 U825 (.ZN(n561), 
	.B2(n560), 
	.B1(FE_OFN4_n319), 
	.A2(n559), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U826 (.ZN(n3370), 
	.B2(n219), 
	.B1(n551), 
	.A2(n6407), 
	.A1(n5409));
   OAI22_X1 U827 (.ZN(n3371), 
	.B2(n221), 
	.B1(n551), 
	.A2(n6410), 
	.A1(n5377));
   OAI22_X1 U828 (.ZN(n3372), 
	.B2(n223), 
	.B1(n551), 
	.A2(n6401), 
	.A1(n5345));
   OAI22_X1 U829 (.ZN(n3373), 
	.B2(n225), 
	.B1(n551), 
	.A2(n6406), 
	.A1(n5313));
   OAI22_X1 U830 (.ZN(n3374), 
	.B2(n227), 
	.B1(n551), 
	.A2(n6399), 
	.A1(n5281));
   OAI22_X1 U831 (.ZN(n3375), 
	.B2(n229), 
	.B1(n551), 
	.A2(n6404), 
	.A1(n5249));
   OAI22_X1 U832 (.ZN(n3376), 
	.B2(n231), 
	.B1(n551), 
	.A2(n6398), 
	.A1(n5217));
   OAI22_X1 U833 (.ZN(n3377), 
	.B2(n233), 
	.B1(n551), 
	.A2(n6396), 
	.A1(n5185));
   OAI22_X1 U834 (.ZN(n3378), 
	.B2(n235), 
	.B1(n551), 
	.A2(n6393), 
	.A1(n5153));
   OAI22_X1 U835 (.ZN(n3379), 
	.B2(n237), 
	.B1(n551), 
	.A2(n6391), 
	.A1(n5121));
   OAI22_X1 U836 (.ZN(n3380), 
	.B2(n239), 
	.B1(n551), 
	.A2(n6390), 
	.A1(n5089));
   OAI22_X1 U837 (.ZN(n3381), 
	.B2(n241), 
	.B1(n551), 
	.A2(n6388), 
	.A1(n5057));
   OAI22_X1 U838 (.ZN(n3382), 
	.B2(n243), 
	.B1(n551), 
	.A2(n6385), 
	.A1(n5025));
   OAI22_X1 U839 (.ZN(n3383), 
	.B2(n245), 
	.B1(n551), 
	.A2(n6383), 
	.A1(n4993));
   OAI22_X1 U840 (.ZN(n3384), 
	.B2(n247), 
	.B1(n551), 
	.A2(n6382), 
	.A1(n4961));
   OAI22_X1 U841 (.ZN(n3385), 
	.B2(n249), 
	.B1(n551), 
	.A2(n6380), 
	.A1(n4929));
   OAI22_X1 U842 (.ZN(n3386), 
	.B2(n251), 
	.B1(n551), 
	.A2(n6384), 
	.A1(n4897));
   OAI22_X1 U843 (.ZN(n3387), 
	.B2(n253), 
	.B1(n551), 
	.A2(n6381), 
	.A1(n4865));
   OAI22_X1 U844 (.ZN(n3388), 
	.B2(n255), 
	.B1(n551), 
	.A2(n6387), 
	.A1(n4833));
   OAI22_X1 U845 (.ZN(n3389), 
	.B2(n257), 
	.B1(n551), 
	.A2(n6386), 
	.A1(n4801));
   OAI22_X1 U846 (.ZN(n3390), 
	.B2(n259), 
	.B1(n551), 
	.A2(n6392), 
	.A1(n4769));
   OAI22_X1 U847 (.ZN(n3391), 
	.B2(n261), 
	.B1(n551), 
	.A2(n6394), 
	.A1(n4737));
   OAI22_X1 U848 (.ZN(n3392), 
	.B2(n263), 
	.B1(n551), 
	.A2(n6389), 
	.A1(n4705));
   OAI22_X1 U849 (.ZN(n3393), 
	.B2(n265), 
	.B1(n551), 
	.A2(n6395), 
	.A1(n4673));
   OAI22_X1 U850 (.ZN(n3394), 
	.B2(n267), 
	.B1(n551), 
	.A2(n6400), 
	.A1(n4641));
   OAI22_X1 U851 (.ZN(n3395), 
	.B2(n269), 
	.B1(n551), 
	.A2(n6402), 
	.A1(n4609));
   OAI22_X1 U852 (.ZN(n3396), 
	.B2(n271), 
	.B1(n551), 
	.A2(n6397), 
	.A1(n4577));
   OAI22_X1 U853 (.ZN(n3397), 
	.B2(n273), 
	.B1(n551), 
	.A2(n6403), 
	.A1(n4545));
   OAI22_X1 U854 (.ZN(n3398), 
	.B2(n275), 
	.B1(n551), 
	.A2(n6408), 
	.A1(n4513));
   OAI22_X1 U855 (.ZN(n3399), 
	.B2(n277), 
	.B1(n551), 
	.A2(n6405), 
	.A1(n4481));
   OAI22_X1 U856 (.ZN(n3400), 
	.B2(n279), 
	.B1(n551), 
	.A2(n6411), 
	.A1(n4449));
   OAI211_X1 U858 (.ZN(n560), 
	.C2(n562), 
	.C1(n482), 
	.B(n563), 
	.A(n484));
   AOI22_X1 U859 (.ZN(n563), 
	.B2(n489), 
	.B1(n565), 
	.A2(n564), 
	.A1(n486));
   INV_X1 U860 (.ZN(n565), 
	.A(n5518));
   INV_X1 U861 (.ZN(n562), 
	.A(n5799));
   OAI22_X1 U862 (.ZN(n3401), 
	.B2(n550), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5518));
   INV_X1 U863 (.ZN(n550), 
	.A(n566));
   OAI211_X1 U864 (.ZN(n566), 
	.C2(n321), 
	.C1(n5670), 
	.B(n568), 
	.A(n567));
   AOI222_X1 U865 (.ZN(n568), 
	.C2(n570), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[12] ), 
	.A2(n569), 
	.A1(FE_OFN91_n285));
   INV_X1 U866 (.ZN(n570), 
	.A(n5706));
   AOI22_X1 U867 (.ZN(n567), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[12] ), 
	.A2(n6203), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U868 (.ZN(n3402), 
	.B2(n2671), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n571));
   OAI221_X1 U869 (.ZN(n3403), 
	.C2(n71), 
	.C1(n92), 
	.B2(n69), 
	.B1(n572), 
	.A(n573));
   NAND2_X1 U870 (.ZN(n573), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [11]));
   OAI222_X1 U871 (.ZN(n3404), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N62 ), 
	.B2(n300), 
	.B1(n572), 
	.A2(n123), 
	.A1(n92));
   INV_X1 U872 (.ZN(n572), 
	.A(\UUT/break_code[11] ));
   INV_X1 U873 (.ZN(n92), 
	.A(n574));
   OAI222_X1 U874 (.ZN(n574), 
	.C2(n132), 
	.C1(n5520), 
	.B2(n131), 
	.B1(n576), 
	.A2(n129), 
	.A1(n575));
   OAI221_X1 U875 (.ZN(n3405), 
	.C2(n135), 
	.C1(n5707), 
	.B2(n577), 
	.B1(n133), 
	.A(n578));
   AOI22_X1 U876 (.ZN(n578), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [43]), 
	.A2(n579), 
	.A1(n137));
   OAI221_X1 U877 (.ZN(n3406), 
	.C2(n142), 
	.C1(n5672), 
	.B2(n580), 
	.B1(n140), 
	.A(n581));
   AOI22_X1 U878 (.ZN(n581), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [11]), 
	.A2(n579), 
	.A1(n144));
   INV_X1 U879 (.ZN(n579), 
	.A(n5673));
   OAI22_X1 U880 (.ZN(n3407), 
	.B2(net54873), 
	.B1(n5673), 
	.A2(n582), 
	.A1(net54953));
   OAI221_X1 U881 (.ZN(n3408), 
	.C2(n582), 
	.C1(n147), 
	.B2(n310), 
	.B1(n575), 
	.A(n583));
   AOI22_X1 U882 (.ZN(n583), 
	.B2(n585), 
	.B1(FE_OFN6_n314), 
	.A2(n584), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U883 (.ZN(n582), 
	.A(FE_OFN146_UUT_Mpath_the_mult_x_operand1_11_));
   OAI221_X1 U884 (.ZN(n3409), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N61 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n575), 
	.A(n586));
   AOI22_X1 U885 (.ZN(n586), 
	.B2(n585), 
	.B1(FE_OFN4_n319), 
	.A2(n584), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U886 (.ZN(n3410), 
	.B2(n219), 
	.B1(n576), 
	.A2(n6407), 
	.A1(n5410));
   OAI22_X1 U887 (.ZN(n3411), 
	.B2(n221), 
	.B1(n576), 
	.A2(n6410), 
	.A1(n5378));
   OAI22_X1 U888 (.ZN(n3412), 
	.B2(n223), 
	.B1(n576), 
	.A2(n6401), 
	.A1(n5346));
   OAI22_X1 U889 (.ZN(n3413), 
	.B2(n225), 
	.B1(n576), 
	.A2(n6406), 
	.A1(n5314));
   OAI22_X1 U890 (.ZN(n3414), 
	.B2(n227), 
	.B1(n576), 
	.A2(n6399), 
	.A1(n5282));
   OAI22_X1 U891 (.ZN(n3415), 
	.B2(n229), 
	.B1(n576), 
	.A2(n6404), 
	.A1(n5250));
   OAI22_X1 U892 (.ZN(n3416), 
	.B2(n231), 
	.B1(n576), 
	.A2(n6398), 
	.A1(n5218));
   OAI22_X1 U893 (.ZN(n3417), 
	.B2(n233), 
	.B1(n576), 
	.A2(n6396), 
	.A1(n5186));
   OAI22_X1 U894 (.ZN(n3418), 
	.B2(n235), 
	.B1(n576), 
	.A2(n6393), 
	.A1(n5154));
   OAI22_X1 U895 (.ZN(n3419), 
	.B2(n237), 
	.B1(n576), 
	.A2(n6391), 
	.A1(n5122));
   OAI22_X1 U896 (.ZN(n3420), 
	.B2(n239), 
	.B1(n576), 
	.A2(n6390), 
	.A1(n5090));
   OAI22_X1 U897 (.ZN(n3421), 
	.B2(n241), 
	.B1(n576), 
	.A2(n6388), 
	.A1(n5058));
   OAI22_X1 U898 (.ZN(n3422), 
	.B2(n243), 
	.B1(n576), 
	.A2(n6385), 
	.A1(n5026));
   OAI22_X1 U899 (.ZN(n3423), 
	.B2(n245), 
	.B1(n576), 
	.A2(n6383), 
	.A1(n4994));
   OAI22_X1 U900 (.ZN(n3424), 
	.B2(n247), 
	.B1(n576), 
	.A2(n6382), 
	.A1(n4962));
   OAI22_X1 U901 (.ZN(n3425), 
	.B2(n249), 
	.B1(n576), 
	.A2(n6380), 
	.A1(n4930));
   OAI22_X1 U902 (.ZN(n3426), 
	.B2(n251), 
	.B1(n576), 
	.A2(n6384), 
	.A1(n4898));
   OAI22_X1 U903 (.ZN(n3427), 
	.B2(n253), 
	.B1(n576), 
	.A2(n6381), 
	.A1(n4866));
   OAI22_X1 U904 (.ZN(n3428), 
	.B2(n255), 
	.B1(n576), 
	.A2(n6387), 
	.A1(n4834));
   OAI22_X1 U905 (.ZN(n3429), 
	.B2(n257), 
	.B1(n576), 
	.A2(n6386), 
	.A1(n4802));
   OAI22_X1 U906 (.ZN(n3430), 
	.B2(n259), 
	.B1(n576), 
	.A2(n6392), 
	.A1(n4770));
   OAI22_X1 U907 (.ZN(n3431), 
	.B2(n261), 
	.B1(n576), 
	.A2(n6394), 
	.A1(n4738));
   OAI22_X1 U908 (.ZN(n3432), 
	.B2(n263), 
	.B1(n576), 
	.A2(n6389), 
	.A1(n4706));
   OAI22_X1 U909 (.ZN(n3433), 
	.B2(n265), 
	.B1(n576), 
	.A2(n6395), 
	.A1(n4674));
   OAI22_X1 U910 (.ZN(n3434), 
	.B2(n267), 
	.B1(n576), 
	.A2(n6400), 
	.A1(n4642));
   OAI22_X1 U911 (.ZN(n3435), 
	.B2(n269), 
	.B1(n576), 
	.A2(n6402), 
	.A1(n4610));
   OAI22_X1 U912 (.ZN(n3436), 
	.B2(n271), 
	.B1(n576), 
	.A2(n6397), 
	.A1(n4578));
   OAI22_X1 U913 (.ZN(n3437), 
	.B2(n273), 
	.B1(n576), 
	.A2(n6403), 
	.A1(n4546));
   OAI22_X1 U914 (.ZN(n3438), 
	.B2(n275), 
	.B1(n576), 
	.A2(n6408), 
	.A1(n4514));
   OAI22_X1 U915 (.ZN(n3439), 
	.B2(n277), 
	.B1(n576), 
	.A2(n6405), 
	.A1(n4482));
   OAI22_X1 U916 (.ZN(n3440), 
	.B2(n279), 
	.B1(n576), 
	.A2(n6411), 
	.A1(n4450));
   OAI211_X1 U918 (.ZN(n585), 
	.C2(n587), 
	.C1(n482), 
	.B(n588), 
	.A(n484));
   AOI22_X1 U919 (.ZN(n588), 
	.B2(n489), 
	.B1(n590), 
	.A2(n589), 
	.A1(n486));
   INV_X1 U920 (.ZN(n590), 
	.A(n5521));
   INV_X1 U921 (.ZN(n587), 
	.A(n5812));
   OAI22_X1 U922 (.ZN(n3441), 
	.B2(n575), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5521));
   INV_X1 U923 (.ZN(n575), 
	.A(n591));
   OAI211_X1 U924 (.ZN(n591), 
	.C2(n321), 
	.C1(n5672), 
	.B(n593), 
	.A(n592));
   AOI222_X1 U925 (.ZN(n593), 
	.C2(n595), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[11] ), 
	.A2(n594), 
	.A1(FE_OFN91_n285));
   INV_X1 U926 (.ZN(n595), 
	.A(n5707));
   AOI22_X1 U927 (.ZN(n592), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[11] ), 
	.A2(n6204), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U928 (.ZN(n3442), 
	.C2(n135), 
	.C1(n5708), 
	.B2(n596), 
	.B1(n133), 
	.A(n597));
   AOI22_X1 U929 (.ZN(n597), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [42]), 
	.A2(n598), 
	.A1(n137));
   OAI221_X1 U930 (.ZN(n3443), 
	.C2(n142), 
	.C1(n5674), 
	.B2(n599), 
	.B1(n140), 
	.A(n600));
   AOI22_X1 U931 (.ZN(n600), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [10]), 
	.A2(n598), 
	.A1(n144));
   INV_X1 U932 (.ZN(n598), 
	.A(n5675));
   OAI22_X1 U933 (.ZN(n3444), 
	.B2(net54871), 
	.B1(n5675), 
	.A2(n601), 
	.A1(net54953));
   OAI221_X1 U934 (.ZN(n3445), 
	.C2(n601), 
	.C1(n147), 
	.B2(n310), 
	.B1(n602), 
	.A(n603));
   AOI22_X1 U935 (.ZN(n603), 
	.B2(n605), 
	.B1(FE_OFN6_n314), 
	.A2(n604), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U936 (.ZN(n601), 
	.A(\UUT/Mpath/the_mult/x_operand1[10] ));
   OAI221_X1 U937 (.ZN(n3446), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N63 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n602), 
	.A(n606));
   AOI22_X1 U938 (.ZN(n606), 
	.B2(n605), 
	.B1(FE_OFN4_n319), 
	.A2(n604), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U939 (.ZN(n3447), 
	.B2(n602), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5524));
   OAI221_X1 U940 (.ZN(n3448), 
	.C2(n71), 
	.C1(n91), 
	.B2(n69), 
	.B1(n607), 
	.A(n608));
   NAND2_X1 U941 (.ZN(n608), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [9]));
   OAI222_X1 U942 (.ZN(n3449), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N66 ), 
	.B2(n300), 
	.B1(n607), 
	.A2(n123), 
	.A1(n91));
   INV_X1 U943 (.ZN(n607), 
	.A(\UUT/break_code[9] ));
   INV_X1 U944 (.ZN(n91), 
	.A(n609));
   OAI222_X1 U945 (.ZN(n609), 
	.C2(n132), 
	.C1(n5431), 
	.B2(n131), 
	.B1(n611), 
	.A2(n129), 
	.A1(n610));
   OAI221_X1 U946 (.ZN(n3450), 
	.C2(n135), 
	.C1(n5678), 
	.B2(n612), 
	.B1(n133), 
	.A(n613));
   AOI22_X1 U947 (.ZN(n613), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [41]), 
	.A2(n614), 
	.A1(n137));
   OAI221_X1 U948 (.ZN(n3451), 
	.C2(n142), 
	.C1(n5614), 
	.B2(n615), 
	.B1(n140), 
	.A(n616));
   AOI22_X1 U949 (.ZN(n616), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [9]), 
	.A2(n614), 
	.A1(n144));
   INV_X1 U950 (.ZN(n614), 
	.A(n5615));
   OAI22_X1 U951 (.ZN(n3452), 
	.B2(net54871), 
	.B1(n5615), 
	.A2(n617), 
	.A1(net54953));
   OAI221_X1 U952 (.ZN(n3453), 
	.C2(n617), 
	.C1(n147), 
	.B2(n310), 
	.B1(n610), 
	.A(n618));
   AOI22_X1 U953 (.ZN(n618), 
	.B2(n620), 
	.B1(FE_OFN6_n314), 
	.A2(n619), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U954 (.ZN(n617), 
	.A(FE_OFN149_UUT_Mpath_the_mult_x_operand1_9_));
   OAI221_X1 U955 (.ZN(n3454), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N65 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n610), 
	.A(n621));
   AOI22_X1 U956 (.ZN(n621), 
	.B2(n620), 
	.B1(FE_OFN4_n319), 
	.A2(n619), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U957 (.ZN(n3455), 
	.B2(n219), 
	.B1(n611), 
	.A2(n6407), 
	.A1(n5381));
   OAI22_X1 U958 (.ZN(n3456), 
	.B2(n221), 
	.B1(n611), 
	.A2(n6410), 
	.A1(n5349));
   OAI22_X1 U959 (.ZN(n3457), 
	.B2(n223), 
	.B1(n611), 
	.A2(n6401), 
	.A1(n5317));
   OAI22_X1 U960 (.ZN(n3458), 
	.B2(n225), 
	.B1(n611), 
	.A2(n6406), 
	.A1(n5285));
   OAI22_X1 U961 (.ZN(n3459), 
	.B2(n227), 
	.B1(n611), 
	.A2(n6399), 
	.A1(n5253));
   OAI22_X1 U962 (.ZN(n3460), 
	.B2(n229), 
	.B1(n611), 
	.A2(n6404), 
	.A1(n5221));
   OAI22_X1 U963 (.ZN(n3461), 
	.B2(n231), 
	.B1(n611), 
	.A2(n6398), 
	.A1(n5189));
   OAI22_X1 U964 (.ZN(n3462), 
	.B2(n233), 
	.B1(n611), 
	.A2(n6396), 
	.A1(n5157));
   OAI22_X1 U965 (.ZN(n3463), 
	.B2(n235), 
	.B1(n611), 
	.A2(n6393), 
	.A1(n5125));
   OAI22_X1 U966 (.ZN(n3464), 
	.B2(n237), 
	.B1(n611), 
	.A2(n6391), 
	.A1(n5093));
   OAI22_X1 U967 (.ZN(n3465), 
	.B2(n239), 
	.B1(n611), 
	.A2(n6390), 
	.A1(n5061));
   OAI22_X1 U968 (.ZN(n3466), 
	.B2(n241), 
	.B1(n611), 
	.A2(n6388), 
	.A1(n5029));
   OAI22_X1 U969 (.ZN(n3467), 
	.B2(n243), 
	.B1(n611), 
	.A2(n6385), 
	.A1(n4997));
   OAI22_X1 U970 (.ZN(n3468), 
	.B2(n245), 
	.B1(n611), 
	.A2(n6383), 
	.A1(n4965));
   OAI22_X1 U971 (.ZN(n3469), 
	.B2(n247), 
	.B1(n611), 
	.A2(n6382), 
	.A1(n4933));
   OAI22_X1 U972 (.ZN(n3470), 
	.B2(n249), 
	.B1(n611), 
	.A2(n6380), 
	.A1(n4901));
   OAI22_X1 U973 (.ZN(n3471), 
	.B2(n251), 
	.B1(n611), 
	.A2(n6384), 
	.A1(n4869));
   OAI22_X1 U974 (.ZN(n3472), 
	.B2(n253), 
	.B1(n611), 
	.A2(n6381), 
	.A1(n4837));
   OAI22_X1 U975 (.ZN(n3473), 
	.B2(n255), 
	.B1(n611), 
	.A2(n6387), 
	.A1(n4805));
   OAI22_X1 U976 (.ZN(n3474), 
	.B2(n257), 
	.B1(n611), 
	.A2(n6386), 
	.A1(n4773));
   OAI22_X1 U977 (.ZN(n3475), 
	.B2(n259), 
	.B1(n611), 
	.A2(n6392), 
	.A1(n4741));
   OAI22_X1 U978 (.ZN(n3476), 
	.B2(n261), 
	.B1(n611), 
	.A2(n6394), 
	.A1(n4709));
   OAI22_X1 U979 (.ZN(n3477), 
	.B2(n263), 
	.B1(n611), 
	.A2(n6389), 
	.A1(n4677));
   OAI22_X1 U980 (.ZN(n3478), 
	.B2(n265), 
	.B1(n611), 
	.A2(n6395), 
	.A1(n4645));
   OAI22_X1 U981 (.ZN(n3479), 
	.B2(n267), 
	.B1(n611), 
	.A2(n6400), 
	.A1(n4613));
   OAI22_X1 U982 (.ZN(n3480), 
	.B2(n269), 
	.B1(n611), 
	.A2(n6402), 
	.A1(n4581));
   OAI22_X1 U983 (.ZN(n3481), 
	.B2(n271), 
	.B1(n611), 
	.A2(n6397), 
	.A1(n4549));
   OAI22_X1 U984 (.ZN(n3482), 
	.B2(n273), 
	.B1(n611), 
	.A2(n6403), 
	.A1(n4517));
   OAI22_X1 U985 (.ZN(n3483), 
	.B2(n275), 
	.B1(n611), 
	.A2(n6408), 
	.A1(n4485));
   OAI22_X1 U986 (.ZN(n3484), 
	.B2(n277), 
	.B1(n611), 
	.A2(n6405), 
	.A1(n4453));
   OAI22_X1 U987 (.ZN(n3485), 
	.B2(n279), 
	.B1(n611), 
	.A2(n6411), 
	.A1(n4421));
   OAI211_X1 U989 (.ZN(n620), 
	.C2(n622), 
	.C1(n482), 
	.B(n623), 
	.A(n484));
   AOI22_X1 U990 (.ZN(n623), 
	.B2(n489), 
	.B1(n625), 
	.A2(n624), 
	.A1(n486));
   INV_X1 U991 (.ZN(n625), 
	.A(n5433));
   INV_X1 U992 (.ZN(n622), 
	.A(n5712));
   OAI22_X1 U993 (.ZN(n3486), 
	.B2(n610), 
	.B1(FE_OFN12_net54953), 
	.A2(net54877), 
	.A1(n5433));
   INV_X1 U994 (.ZN(n610), 
	.A(n626));
   OAI211_X1 U995 (.ZN(n626), 
	.C2(n321), 
	.C1(n5614), 
	.B(n628), 
	.A(n627));
   AOI222_X1 U996 (.ZN(n628), 
	.C2(n630), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[9] ), 
	.A2(n629), 
	.A1(FE_OFN91_n285));
   INV_X1 U997 (.ZN(n630), 
	.A(n5678));
   AOI22_X1 U998 (.ZN(n627), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[9] ), 
	.A2(n6189), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U999 (.ZN(n3487), 
	.B2(n2677), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n631));
   OAI221_X1 U1000 (.ZN(n3488), 
	.C2(n135), 
	.C1(n5679), 
	.B2(n632), 
	.B1(n133), 
	.A(n633));
   AOI22_X1 U1001 (.ZN(n633), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [40]), 
	.A2(n634), 
	.A1(n137));
   OAI221_X1 U1002 (.ZN(n3489), 
	.C2(n142), 
	.C1(n5616), 
	.B2(n635), 
	.B1(n140), 
	.A(n636));
   AOI22_X1 U1003 (.ZN(n636), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [8]), 
	.A2(n634), 
	.A1(n144));
   INV_X1 U1004 (.ZN(n634), 
	.A(n5617));
   OAI22_X1 U1005 (.ZN(n3490), 
	.B2(net54875), 
	.B1(n5617), 
	.A2(n637), 
	.A1(net54953));
   OAI221_X1 U1006 (.ZN(n3491), 
	.C2(n637), 
	.C1(n147), 
	.B2(n310), 
	.B1(n638), 
	.A(n639));
   AOI22_X1 U1007 (.ZN(n639), 
	.B2(n641), 
	.B1(FE_OFN6_n314), 
	.A2(n640), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1008 (.ZN(n637), 
	.A(\UUT/Mpath/the_mult/x_operand1[8] ));
   OAI221_X1 U1009 (.ZN(n3492), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N67 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n638), 
	.A(n642));
   AOI22_X1 U1010 (.ZN(n642), 
	.B2(n641), 
	.B1(FE_OFN4_n319), 
	.A2(n640), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1011 (.ZN(n3493), 
	.B2(n638), 
	.B1(FE_OFN12_net54953), 
	.A2(net54879), 
	.A1(n5437));
   OAI22_X1 U1012 (.ZN(n3494), 
	.B2(n2679), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n643));
   OAI221_X1 U1013 (.ZN(n3495), 
	.C2(n71), 
	.C1(n90), 
	.B2(n69), 
	.B1(n644), 
	.A(n645));
   NAND2_X1 U1014 (.ZN(n645), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [7]));
   OAI222_X1 U1015 (.ZN(n3496), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N70 ), 
	.B2(n300), 
	.B1(n644), 
	.A2(n123), 
	.A1(n90));
   INV_X1 U1016 (.ZN(n644), 
	.A(\UUT/break_code[7] ));
   INV_X1 U1017 (.ZN(n90), 
	.A(n646));
   OAI222_X1 U1018 (.ZN(n646), 
	.C2(n132), 
	.C1(n5439), 
	.B2(n131), 
	.B1(n648), 
	.A2(n129), 
	.A1(n647));
   OAI221_X1 U1019 (.ZN(n3497), 
	.C2(n135), 
	.C1(n5680), 
	.B2(n649), 
	.B1(n133), 
	.A(n650));
   AOI22_X1 U1020 (.ZN(n650), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [39]), 
	.A2(n651), 
	.A1(n137));
   OAI221_X1 U1021 (.ZN(n3498), 
	.C2(n142), 
	.C1(n5618), 
	.B2(n652), 
	.B1(n140), 
	.A(n653));
   AOI22_X1 U1022 (.ZN(n653), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [7]), 
	.A2(n651), 
	.A1(n144));
   INV_X1 U1023 (.ZN(n651), 
	.A(n5619));
   OAI22_X1 U1024 (.ZN(n3499), 
	.B2(net54871), 
	.B1(n5619), 
	.A2(n654), 
	.A1(net54953));
   OAI221_X1 U1025 (.ZN(n3500), 
	.C2(n654), 
	.C1(n147), 
	.B2(n310), 
	.B1(n647), 
	.A(n655));
   AOI22_X1 U1026 (.ZN(n655), 
	.B2(n657), 
	.B1(FE_OFN6_n314), 
	.A2(n656), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1027 (.ZN(n654), 
	.A(FE_OFN152_UUT_Mpath_the_mult_x_operand1_7_));
   OAI221_X1 U1028 (.ZN(n3501), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N69 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n647), 
	.A(n658));
   AOI22_X1 U1029 (.ZN(n658), 
	.B2(n657), 
	.B1(FE_OFN4_n319), 
	.A2(n656), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1030 (.ZN(n3502), 
	.B2(n219), 
	.B1(n648), 
	.A2(n6407), 
	.A1(n5383));
   OAI22_X1 U1031 (.ZN(n3503), 
	.B2(n221), 
	.B1(n648), 
	.A2(n6410), 
	.A1(n5351));
   OAI22_X1 U1032 (.ZN(n3504), 
	.B2(n223), 
	.B1(n648), 
	.A2(n6401), 
	.A1(n5319));
   OAI22_X1 U1033 (.ZN(n3505), 
	.B2(n225), 
	.B1(n648), 
	.A2(n6406), 
	.A1(n5287));
   OAI22_X1 U1034 (.ZN(n3506), 
	.B2(n227), 
	.B1(n648), 
	.A2(n6399), 
	.A1(n5255));
   OAI22_X1 U1035 (.ZN(n3507), 
	.B2(n229), 
	.B1(n648), 
	.A2(n6404), 
	.A1(n5223));
   OAI22_X1 U1036 (.ZN(n3508), 
	.B2(n231), 
	.B1(n648), 
	.A2(n6398), 
	.A1(n5191));
   OAI22_X1 U1037 (.ZN(n3509), 
	.B2(n233), 
	.B1(n648), 
	.A2(n6396), 
	.A1(n5159));
   OAI22_X1 U1038 (.ZN(n3510), 
	.B2(n235), 
	.B1(n648), 
	.A2(n6393), 
	.A1(n5127));
   OAI22_X1 U1039 (.ZN(n3511), 
	.B2(n237), 
	.B1(n648), 
	.A2(n6391), 
	.A1(n5095));
   OAI22_X1 U1040 (.ZN(n3512), 
	.B2(n239), 
	.B1(n648), 
	.A2(n6390), 
	.A1(n5063));
   OAI22_X1 U1041 (.ZN(n3513), 
	.B2(n241), 
	.B1(n648), 
	.A2(n6388), 
	.A1(n5031));
   OAI22_X1 U1042 (.ZN(n3514), 
	.B2(n243), 
	.B1(n648), 
	.A2(n6385), 
	.A1(n4999));
   OAI22_X1 U1043 (.ZN(n3515), 
	.B2(n245), 
	.B1(n648), 
	.A2(n6383), 
	.A1(n4967));
   OAI22_X1 U1044 (.ZN(n3516), 
	.B2(n247), 
	.B1(n648), 
	.A2(n6382), 
	.A1(n4935));
   OAI22_X1 U1045 (.ZN(n3517), 
	.B2(n249), 
	.B1(n648), 
	.A2(n6380), 
	.A1(n4903));
   OAI22_X1 U1046 (.ZN(n3518), 
	.B2(n251), 
	.B1(n648), 
	.A2(n6384), 
	.A1(n4871));
   OAI22_X1 U1047 (.ZN(n3519), 
	.B2(n253), 
	.B1(n648), 
	.A2(n6381), 
	.A1(n4839));
   OAI22_X1 U1048 (.ZN(n3520), 
	.B2(n255), 
	.B1(n648), 
	.A2(n6387), 
	.A1(n4807));
   OAI22_X1 U1049 (.ZN(n3521), 
	.B2(n257), 
	.B1(n648), 
	.A2(n6386), 
	.A1(n4775));
   OAI22_X1 U1050 (.ZN(n3522), 
	.B2(n259), 
	.B1(n648), 
	.A2(n6392), 
	.A1(n4743));
   OAI22_X1 U1051 (.ZN(n3523), 
	.B2(n261), 
	.B1(n648), 
	.A2(n6394), 
	.A1(n4711));
   OAI22_X1 U1052 (.ZN(n3524), 
	.B2(n263), 
	.B1(n648), 
	.A2(n6389), 
	.A1(n4679));
   OAI22_X1 U1053 (.ZN(n3525), 
	.B2(n265), 
	.B1(n648), 
	.A2(n6395), 
	.A1(n4647));
   OAI22_X1 U1054 (.ZN(n3526), 
	.B2(n267), 
	.B1(n648), 
	.A2(n6400), 
	.A1(n4615));
   OAI22_X1 U1055 (.ZN(n3527), 
	.B2(n269), 
	.B1(n648), 
	.A2(n6402), 
	.A1(n4583));
   OAI22_X1 U1056 (.ZN(n3528), 
	.B2(n271), 
	.B1(n648), 
	.A2(n6397), 
	.A1(n4551));
   OAI22_X1 U1057 (.ZN(n3529), 
	.B2(n273), 
	.B1(n648), 
	.A2(n6403), 
	.A1(n4519));
   OAI22_X1 U1058 (.ZN(n3530), 
	.B2(n275), 
	.B1(n648), 
	.A2(n6408), 
	.A1(n4487));
   OAI22_X1 U1059 (.ZN(n3531), 
	.B2(n277), 
	.B1(n648), 
	.A2(n6405), 
	.A1(n4455));
   OAI22_X1 U1060 (.ZN(n3532), 
	.B2(n279), 
	.B1(n648), 
	.A2(n6411), 
	.A1(n4423));
   OAI222_X1 U1062 (.ZN(n657), 
	.C2(n5440), 
	.C1(n5710), 
	.B2(n660), 
	.B1(n659), 
	.A2(n489), 
	.A1(n5754));
   AOI221_X1 U1063 (.ZN(n659), 
	.C2(n5755), 
	.C1(n5756), 
	.B2(n487), 
	.B1(n5757), 
	.A(n5759));
   INV_X1 U1064 (.ZN(n487), 
	.A(n5957));
   OAI22_X1 U1065 (.ZN(n3533), 
	.B2(n647), 
	.B1(FE_OFN12_net54953), 
	.A2(net54881), 
	.A1(n5440));
   INV_X1 U1066 (.ZN(n647), 
	.A(n661));
   OAI211_X1 U1067 (.ZN(n661), 
	.C2(n321), 
	.C1(n5618), 
	.B(n663), 
	.A(n662));
   AOI222_X1 U1068 (.ZN(n663), 
	.C2(n665), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[7] ), 
	.A2(n664), 
	.A1(FE_OFN91_n285));
   INV_X1 U1069 (.ZN(n665), 
	.A(n5680));
   AOI22_X1 U1070 (.ZN(n662), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[7] ), 
	.A2(n6191), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1071 (.ZN(n3534), 
	.B2(n2682), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n666));
   OAI221_X1 U1072 (.ZN(n3535), 
	.C2(n71), 
	.C1(n89), 
	.B2(n69), 
	.B1(n667), 
	.A(n668));
   NAND2_X1 U1073 (.ZN(n668), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [6]));
   OAI222_X1 U1074 (.ZN(n3536), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N72 ), 
	.B2(n300), 
	.B1(n667), 
	.A2(n123), 
	.A1(n89));
   INV_X1 U1075 (.ZN(n667), 
	.A(\UUT/break_code[6] ));
   INV_X1 U1076 (.ZN(n89), 
	.A(n669));
   OAI222_X1 U1077 (.ZN(n669), 
	.C2(n132), 
	.C1(n5442), 
	.B2(n131), 
	.B1(n671), 
	.A2(n129), 
	.A1(n670));
   OAI221_X1 U1078 (.ZN(n3537), 
	.C2(n135), 
	.C1(n5681), 
	.B2(n672), 
	.B1(n133), 
	.A(n673));
   AOI22_X1 U1079 (.ZN(n673), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [38]), 
	.A2(n674), 
	.A1(n137));
   OAI221_X1 U1080 (.ZN(n3538), 
	.C2(n142), 
	.C1(n5620), 
	.B2(n675), 
	.B1(n140), 
	.A(n676));
   AOI22_X1 U1081 (.ZN(n676), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [6]), 
	.A2(n674), 
	.A1(n144));
   INV_X1 U1082 (.ZN(n674), 
	.A(n5621));
   OAI22_X1 U1083 (.ZN(n3539), 
	.B2(net54869), 
	.B1(n5621), 
	.A2(n677), 
	.A1(net54953));
   OAI221_X1 U1084 (.ZN(n3540), 
	.C2(n677), 
	.C1(n147), 
	.B2(n310), 
	.B1(n670), 
	.A(n678));
   AOI22_X1 U1085 (.ZN(n678), 
	.B2(n680), 
	.B1(FE_OFN6_n314), 
	.A2(n679), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1086 (.ZN(n677), 
	.A(\UUT/Mpath/the_mult/x_operand1[6] ));
   OAI221_X1 U1087 (.ZN(n3541), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N71 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n670), 
	.A(n681));
   AOI22_X1 U1088 (.ZN(n681), 
	.B2(n680), 
	.B1(FE_OFN4_n319), 
	.A2(n679), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1089 (.ZN(n3542), 
	.B2(n219), 
	.B1(n671), 
	.A2(n6407), 
	.A1(n5384));
   OAI22_X1 U1090 (.ZN(n3543), 
	.B2(n221), 
	.B1(n671), 
	.A2(n6410), 
	.A1(n5352));
   OAI22_X1 U1091 (.ZN(n3544), 
	.B2(n223), 
	.B1(n671), 
	.A2(n6401), 
	.A1(n5320));
   OAI22_X1 U1092 (.ZN(n3545), 
	.B2(n225), 
	.B1(n671), 
	.A2(n6406), 
	.A1(n5288));
   OAI22_X1 U1093 (.ZN(n3546), 
	.B2(n227), 
	.B1(n671), 
	.A2(n6399), 
	.A1(n5256));
   OAI22_X1 U1094 (.ZN(n3547), 
	.B2(n229), 
	.B1(n671), 
	.A2(n6404), 
	.A1(n5224));
   OAI22_X1 U1095 (.ZN(n3548), 
	.B2(n231), 
	.B1(n671), 
	.A2(n6398), 
	.A1(n5192));
   OAI22_X1 U1096 (.ZN(n3549), 
	.B2(n233), 
	.B1(n671), 
	.A2(n6396), 
	.A1(n5160));
   OAI22_X1 U1097 (.ZN(n3550), 
	.B2(n235), 
	.B1(n671), 
	.A2(n6393), 
	.A1(n5128));
   OAI22_X1 U1098 (.ZN(n3551), 
	.B2(n237), 
	.B1(n671), 
	.A2(n6391), 
	.A1(n5096));
   OAI22_X1 U1099 (.ZN(n3552), 
	.B2(n239), 
	.B1(n671), 
	.A2(n6390), 
	.A1(n5064));
   OAI22_X1 U1100 (.ZN(n3553), 
	.B2(n241), 
	.B1(n671), 
	.A2(n6388), 
	.A1(n5032));
   OAI22_X1 U1101 (.ZN(n3554), 
	.B2(n243), 
	.B1(n671), 
	.A2(n6385), 
	.A1(n5000));
   OAI22_X1 U1102 (.ZN(n3555), 
	.B2(n245), 
	.B1(n671), 
	.A2(n6383), 
	.A1(n4968));
   OAI22_X1 U1103 (.ZN(n3556), 
	.B2(n247), 
	.B1(n671), 
	.A2(n6382), 
	.A1(n4936));
   OAI22_X1 U1104 (.ZN(n3557), 
	.B2(n249), 
	.B1(n671), 
	.A2(n6380), 
	.A1(n4904));
   OAI22_X1 U1105 (.ZN(n3558), 
	.B2(n251), 
	.B1(n671), 
	.A2(n6384), 
	.A1(n4872));
   OAI22_X1 U1106 (.ZN(n3559), 
	.B2(n253), 
	.B1(n671), 
	.A2(n6381), 
	.A1(n4840));
   OAI22_X1 U1107 (.ZN(n3560), 
	.B2(n255), 
	.B1(n671), 
	.A2(n6387), 
	.A1(n4808));
   OAI22_X1 U1108 (.ZN(n3561), 
	.B2(n257), 
	.B1(n671), 
	.A2(n6386), 
	.A1(n4776));
   OAI22_X1 U1109 (.ZN(n3562), 
	.B2(n259), 
	.B1(n671), 
	.A2(n6392), 
	.A1(n4744));
   OAI22_X1 U1110 (.ZN(n3563), 
	.B2(n261), 
	.B1(n671), 
	.A2(n6394), 
	.A1(n4712));
   OAI22_X1 U1111 (.ZN(n3564), 
	.B2(n263), 
	.B1(n671), 
	.A2(n6389), 
	.A1(n4680));
   OAI22_X1 U1112 (.ZN(n3565), 
	.B2(n265), 
	.B1(n671), 
	.A2(n6395), 
	.A1(n4648));
   OAI22_X1 U1113 (.ZN(n3566), 
	.B2(n267), 
	.B1(n671), 
	.A2(n6400), 
	.A1(n4616));
   OAI22_X1 U1114 (.ZN(n3567), 
	.B2(n269), 
	.B1(n671), 
	.A2(n6402), 
	.A1(n4584));
   OAI22_X1 U1115 (.ZN(n3568), 
	.B2(n271), 
	.B1(n671), 
	.A2(n6397), 
	.A1(n4552));
   OAI22_X1 U1116 (.ZN(n3569), 
	.B2(n273), 
	.B1(n671), 
	.A2(n6403), 
	.A1(n4520));
   OAI22_X1 U1117 (.ZN(n3570), 
	.B2(n275), 
	.B1(n671), 
	.A2(n6408), 
	.A1(n4488));
   OAI22_X1 U1118 (.ZN(n3571), 
	.B2(n277), 
	.B1(n671), 
	.A2(n6405), 
	.A1(n4456));
   OAI22_X1 U1119 (.ZN(n3572), 
	.B2(n279), 
	.B1(n671), 
	.A2(n6411), 
	.A1(n4424));
   OAI211_X1 U1121 (.ZN(n680), 
	.C2(n5443), 
	.C1(n5710), 
	.B(n683), 
	.A(n682));
   AOI222_X1 U1122 (.ZN(n683), 
	.C2(n686), 
	.C1(n5774), 
	.B2(n513), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5769));
   INV_X1 U1123 (.ZN(n513), 
	.A(n5776));
   AOI22_X1 U1124 (.ZN(n682), 
	.B2(n688), 
	.B1(n5771), 
	.A2(n687), 
	.A1(n5775));
   OAI22_X1 U1125 (.ZN(n3573), 
	.B2(n670), 
	.B1(FE_OFN12_net54953), 
	.A2(net54881), 
	.A1(n5443));
   INV_X1 U1126 (.ZN(n670), 
	.A(n689));
   OAI211_X1 U1127 (.ZN(n689), 
	.C2(n321), 
	.C1(n5620), 
	.B(n691), 
	.A(n690));
   AOI222_X1 U1128 (.ZN(n691), 
	.C2(n693), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[6] ), 
	.A2(n692), 
	.A1(FE_OFN91_n285));
   INV_X1 U1129 (.ZN(n693), 
	.A(n5681));
   AOI22_X1 U1130 (.ZN(n690), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[6] ), 
	.A2(n6192), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1131 (.ZN(n3574), 
	.B2(n2685), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n694));
   OAI221_X1 U1132 (.ZN(n3575), 
	.C2(n71), 
	.C1(n88), 
	.B2(n69), 
	.B1(n695), 
	.A(n696));
   NAND2_X1 U1133 (.ZN(n696), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [5]));
   OAI222_X1 U1134 (.ZN(n3576), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N74 ), 
	.B2(n300), 
	.B1(n695), 
	.A2(n123), 
	.A1(n88));
   INV_X1 U1135 (.ZN(n695), 
	.A(\UUT/break_code[5] ));
   INV_X1 U1136 (.ZN(n88), 
	.A(n697));
   OAI222_X1 U1137 (.ZN(n697), 
	.C2(n132), 
	.C1(n5445), 
	.B2(n131), 
	.B1(n699), 
	.A2(n129), 
	.A1(n698));
   OAI221_X1 U1138 (.ZN(n3577), 
	.C2(n135), 
	.C1(n5682), 
	.B2(n700), 
	.B1(n133), 
	.A(n701));
   AOI22_X1 U1139 (.ZN(n701), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [37]), 
	.A2(n702), 
	.A1(n137));
   OAI221_X1 U1140 (.ZN(n3578), 
	.C2(n142), 
	.C1(n5622), 
	.B2(n703), 
	.B1(n140), 
	.A(n704));
   AOI22_X1 U1141 (.ZN(n704), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [5]), 
	.A2(n702), 
	.A1(n144));
   INV_X1 U1142 (.ZN(n702), 
	.A(n5623));
   OAI22_X1 U1143 (.ZN(n3579), 
	.B2(net54869), 
	.B1(n5623), 
	.A2(n705), 
	.A1(FE_OFN10_net54953));
   OAI221_X1 U1144 (.ZN(n3580), 
	.C2(n705), 
	.C1(n147), 
	.B2(n310), 
	.B1(n698), 
	.A(n706));
   AOI22_X1 U1145 (.ZN(n706), 
	.B2(n708), 
	.B1(FE_OFN6_n314), 
	.A2(n707), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1146 (.ZN(n705), 
	.A(FE_OFN156_UUT_Mpath_the_mult_x_operand1_5_));
   OAI221_X1 U1147 (.ZN(n3581), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N73 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n698), 
	.A(n709));
   AOI22_X1 U1148 (.ZN(n709), 
	.B2(n708), 
	.B1(FE_OFN4_n319), 
	.A2(n707), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1149 (.ZN(n3582), 
	.B2(n219), 
	.B1(n699), 
	.A2(n6407), 
	.A1(n5385));
   OAI22_X1 U1150 (.ZN(n3583), 
	.B2(n221), 
	.B1(n699), 
	.A2(n6410), 
	.A1(n5353));
   OAI22_X1 U1151 (.ZN(n3584), 
	.B2(n223), 
	.B1(n699), 
	.A2(n6401), 
	.A1(n5321));
   OAI22_X1 U1152 (.ZN(n3585), 
	.B2(n225), 
	.B1(n699), 
	.A2(n6406), 
	.A1(n5289));
   OAI22_X1 U1153 (.ZN(n3586), 
	.B2(n227), 
	.B1(n699), 
	.A2(n6399), 
	.A1(n5257));
   OAI22_X1 U1154 (.ZN(n3587), 
	.B2(n229), 
	.B1(n699), 
	.A2(n6404), 
	.A1(n5225));
   OAI22_X1 U1155 (.ZN(n3588), 
	.B2(n231), 
	.B1(n699), 
	.A2(n6398), 
	.A1(n5193));
   OAI22_X1 U1156 (.ZN(n3589), 
	.B2(n233), 
	.B1(n699), 
	.A2(n6396), 
	.A1(n5161));
   OAI22_X1 U1157 (.ZN(n3590), 
	.B2(n235), 
	.B1(n699), 
	.A2(n6393), 
	.A1(n5129));
   OAI22_X1 U1158 (.ZN(n3591), 
	.B2(n237), 
	.B1(n699), 
	.A2(n6391), 
	.A1(n5097));
   OAI22_X1 U1159 (.ZN(n3592), 
	.B2(n239), 
	.B1(n699), 
	.A2(n6390), 
	.A1(n5065));
   OAI22_X1 U1160 (.ZN(n3593), 
	.B2(n241), 
	.B1(n699), 
	.A2(n6388), 
	.A1(n5033));
   OAI22_X1 U1161 (.ZN(n3594), 
	.B2(n243), 
	.B1(n699), 
	.A2(n6385), 
	.A1(n5001));
   OAI22_X1 U1162 (.ZN(n3595), 
	.B2(n245), 
	.B1(n699), 
	.A2(n6383), 
	.A1(n4969));
   OAI22_X1 U1163 (.ZN(n3596), 
	.B2(n247), 
	.B1(n699), 
	.A2(n6382), 
	.A1(n4937));
   OAI22_X1 U1164 (.ZN(n3597), 
	.B2(n249), 
	.B1(n699), 
	.A2(n6380), 
	.A1(n4905));
   OAI22_X1 U1165 (.ZN(n3598), 
	.B2(n251), 
	.B1(n699), 
	.A2(n6384), 
	.A1(n4873));
   OAI22_X1 U1166 (.ZN(n3599), 
	.B2(n253), 
	.B1(n699), 
	.A2(n6381), 
	.A1(n4841));
   OAI22_X1 U1167 (.ZN(n3600), 
	.B2(n255), 
	.B1(n699), 
	.A2(n6387), 
	.A1(n4809));
   OAI22_X1 U1168 (.ZN(n3601), 
	.B2(n257), 
	.B1(n699), 
	.A2(n6386), 
	.A1(n4777));
   OAI22_X1 U1169 (.ZN(n3602), 
	.B2(n259), 
	.B1(n699), 
	.A2(n6392), 
	.A1(n4745));
   OAI22_X1 U1170 (.ZN(n3603), 
	.B2(n261), 
	.B1(n699), 
	.A2(n6394), 
	.A1(n4713));
   OAI22_X1 U1171 (.ZN(n3604), 
	.B2(n263), 
	.B1(n699), 
	.A2(n6389), 
	.A1(n4681));
   OAI22_X1 U1172 (.ZN(n3605), 
	.B2(n265), 
	.B1(n699), 
	.A2(n6395), 
	.A1(n4649));
   OAI22_X1 U1173 (.ZN(n3606), 
	.B2(n267), 
	.B1(n699), 
	.A2(n6400), 
	.A1(n4617));
   OAI22_X1 U1174 (.ZN(n3607), 
	.B2(n269), 
	.B1(n699), 
	.A2(n6402), 
	.A1(n4585));
   OAI22_X1 U1175 (.ZN(n3608), 
	.B2(n271), 
	.B1(n699), 
	.A2(n6397), 
	.A1(n4553));
   OAI22_X1 U1176 (.ZN(n3609), 
	.B2(n273), 
	.B1(n699), 
	.A2(n6403), 
	.A1(n4521));
   OAI22_X1 U1177 (.ZN(n3610), 
	.B2(n275), 
	.B1(n699), 
	.A2(n6408), 
	.A1(n4489));
   OAI22_X1 U1178 (.ZN(n3611), 
	.B2(n277), 
	.B1(n699), 
	.A2(n6405), 
	.A1(n4457));
   OAI22_X1 U1179 (.ZN(n3612), 
	.B2(n279), 
	.B1(n699), 
	.A2(n6411), 
	.A1(n4425));
   OAI211_X1 U1181 (.ZN(n708), 
	.C2(n5446), 
	.C1(n5710), 
	.B(n711), 
	.A(n710));
   AOI222_X1 U1182 (.ZN(n711), 
	.C2(n686), 
	.C1(n5791), 
	.B2(n538), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5786));
   INV_X1 U1183 (.ZN(n538), 
	.A(n5793));
   AOI22_X1 U1184 (.ZN(n710), 
	.B2(n688), 
	.B1(n5788), 
	.A2(n687), 
	.A1(n5792));
   OAI22_X1 U1185 (.ZN(n3613), 
	.B2(n698), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5446));
   INV_X1 U1186 (.ZN(n698), 
	.A(n712));
   OAI211_X1 U1187 (.ZN(n712), 
	.C2(n321), 
	.C1(n5622), 
	.B(n714), 
	.A(n713));
   AOI222_X1 U1188 (.ZN(n714), 
	.C2(n716), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[5] ), 
	.A2(n715), 
	.A1(FE_OFN91_n285));
   INV_X1 U1189 (.ZN(n716), 
	.A(n5682));
   AOI22_X1 U1190 (.ZN(n713), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[5] ), 
	.A2(n6193), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1191 (.ZN(n3614), 
	.B2(n2688), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n6463));
   OAI221_X1 U1192 (.ZN(n3615), 
	.C2(n71), 
	.C1(n87), 
	.B2(n69), 
	.B1(n718), 
	.A(n719));
   NAND2_X1 U1193 (.ZN(n719), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [4]));
   OAI222_X1 U1194 (.ZN(n3616), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N76 ), 
	.B2(n300), 
	.B1(n718), 
	.A2(n123), 
	.A1(n87));
   INV_X1 U1195 (.ZN(n87), 
	.A(n720));
   OAI222_X1 U1196 (.ZN(n720), 
	.C2(n132), 
	.C1(n5448), 
	.B2(n131), 
	.B1(n722), 
	.A2(n129), 
	.A1(n721));
   OAI221_X1 U1197 (.ZN(n3617), 
	.C2(n135), 
	.C1(n5683), 
	.B2(n723), 
	.B1(n133), 
	.A(n724));
   AOI22_X1 U1198 (.ZN(n724), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [36]), 
	.A2(n725), 
	.A1(n137));
   OAI221_X1 U1199 (.ZN(n3618), 
	.C2(n142), 
	.C1(n5624), 
	.B2(n726), 
	.B1(n140), 
	.A(n727));
   AOI22_X1 U1200 (.ZN(n727), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [4]), 
	.A2(n725), 
	.A1(n144));
   INV_X1 U1201 (.ZN(n725), 
	.A(n5625));
   OAI22_X1 U1202 (.ZN(n3619), 
	.B2(net54869), 
	.B1(n5625), 
	.A2(n728), 
	.A1(net54953));
   OAI221_X1 U1203 (.ZN(n3620), 
	.C2(n728), 
	.C1(n147), 
	.B2(n310), 
	.B1(n721), 
	.A(n729));
   AOI22_X1 U1204 (.ZN(n729), 
	.B2(n731), 
	.B1(FE_OFN6_n314), 
	.A2(n730), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1205 (.ZN(n728), 
	.A(\UUT/Mpath/the_mult/x_operand1[4] ));
   OAI221_X1 U1206 (.ZN(n3621), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N75 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n721), 
	.A(n732));
   AOI22_X1 U1207 (.ZN(n732), 
	.B2(n731), 
	.B1(FE_OFN4_n319), 
	.A2(n730), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1208 (.ZN(n3622), 
	.B2(n219), 
	.B1(n722), 
	.A2(n6407), 
	.A1(n5386));
   OAI22_X1 U1209 (.ZN(n3623), 
	.B2(n221), 
	.B1(n722), 
	.A2(n6410), 
	.A1(n5354));
   OAI22_X1 U1210 (.ZN(n3624), 
	.B2(n223), 
	.B1(n722), 
	.A2(n6401), 
	.A1(n5322));
   OAI22_X1 U1211 (.ZN(n3625), 
	.B2(n225), 
	.B1(n722), 
	.A2(n6406), 
	.A1(n5290));
   OAI22_X1 U1212 (.ZN(n3626), 
	.B2(n227), 
	.B1(n722), 
	.A2(n6399), 
	.A1(n5258));
   OAI22_X1 U1213 (.ZN(n3627), 
	.B2(n229), 
	.B1(n722), 
	.A2(n6404), 
	.A1(n5226));
   OAI22_X1 U1214 (.ZN(n3628), 
	.B2(n231), 
	.B1(n722), 
	.A2(n6398), 
	.A1(n5194));
   OAI22_X1 U1215 (.ZN(n3629), 
	.B2(n233), 
	.B1(n722), 
	.A2(n6396), 
	.A1(n5162));
   OAI22_X1 U1216 (.ZN(n3630), 
	.B2(n235), 
	.B1(n722), 
	.A2(n6393), 
	.A1(n5130));
   OAI22_X1 U1217 (.ZN(n3631), 
	.B2(n237), 
	.B1(n722), 
	.A2(n6391), 
	.A1(n5098));
   OAI22_X1 U1218 (.ZN(n3632), 
	.B2(n239), 
	.B1(n722), 
	.A2(n6390), 
	.A1(n5066));
   OAI22_X1 U1219 (.ZN(n3633), 
	.B2(n241), 
	.B1(n722), 
	.A2(n6388), 
	.A1(n5034));
   OAI22_X1 U1220 (.ZN(n3634), 
	.B2(n243), 
	.B1(n722), 
	.A2(n6385), 
	.A1(n5002));
   OAI22_X1 U1221 (.ZN(n3635), 
	.B2(n245), 
	.B1(n722), 
	.A2(n6383), 
	.A1(n4970));
   OAI22_X1 U1222 (.ZN(n3636), 
	.B2(n247), 
	.B1(n722), 
	.A2(n6382), 
	.A1(n4938));
   OAI22_X1 U1223 (.ZN(n3637), 
	.B2(n249), 
	.B1(n722), 
	.A2(n6380), 
	.A1(n4906));
   OAI22_X1 U1224 (.ZN(n3638), 
	.B2(n251), 
	.B1(n722), 
	.A2(n6384), 
	.A1(n4874));
   OAI22_X1 U1225 (.ZN(n3639), 
	.B2(n253), 
	.B1(n722), 
	.A2(n6381), 
	.A1(n4842));
   OAI22_X1 U1226 (.ZN(n3640), 
	.B2(n255), 
	.B1(n722), 
	.A2(n6387), 
	.A1(n4810));
   OAI22_X1 U1227 (.ZN(n3641), 
	.B2(n257), 
	.B1(n722), 
	.A2(n6386), 
	.A1(n4778));
   OAI22_X1 U1228 (.ZN(n3642), 
	.B2(n259), 
	.B1(n722), 
	.A2(n6392), 
	.A1(n4746));
   OAI22_X1 U1229 (.ZN(n3643), 
	.B2(n261), 
	.B1(n722), 
	.A2(n6394), 
	.A1(n4714));
   OAI22_X1 U1230 (.ZN(n3644), 
	.B2(n263), 
	.B1(n722), 
	.A2(n6389), 
	.A1(n4682));
   OAI22_X1 U1231 (.ZN(n3645), 
	.B2(n265), 
	.B1(n722), 
	.A2(n6395), 
	.A1(n4650));
   OAI22_X1 U1232 (.ZN(n3646), 
	.B2(n267), 
	.B1(n722), 
	.A2(n6400), 
	.A1(n4618));
   OAI22_X1 U1233 (.ZN(n3647), 
	.B2(n269), 
	.B1(n722), 
	.A2(n6402), 
	.A1(n4586));
   OAI22_X1 U1234 (.ZN(n3648), 
	.B2(n271), 
	.B1(n722), 
	.A2(n6397), 
	.A1(n4554));
   OAI22_X1 U1235 (.ZN(n3649), 
	.B2(n273), 
	.B1(n722), 
	.A2(n6403), 
	.A1(n4522));
   OAI22_X1 U1236 (.ZN(n3650), 
	.B2(n275), 
	.B1(n722), 
	.A2(n6408), 
	.A1(n4490));
   OAI22_X1 U1237 (.ZN(n3651), 
	.B2(n277), 
	.B1(n722), 
	.A2(n6405), 
	.A1(n4458));
   OAI22_X1 U1238 (.ZN(n3652), 
	.B2(n279), 
	.B1(n722), 
	.A2(n6411), 
	.A1(n4426));
   OAI211_X1 U1240 (.ZN(n731), 
	.C2(n5449), 
	.C1(n5710), 
	.B(n734), 
	.A(n733));
   AOI222_X1 U1241 (.ZN(n734), 
	.C2(n686), 
	.C1(n5804), 
	.B2(n564), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5799));
   INV_X1 U1242 (.ZN(n564), 
	.A(n5806));
   AOI22_X1 U1243 (.ZN(n733), 
	.B2(n688), 
	.B1(n5801), 
	.A2(n687), 
	.A1(n5805));
   OAI22_X1 U1244 (.ZN(n3653), 
	.B2(n721), 
	.B1(FE_OFN12_net54953), 
	.A2(net54881), 
	.A1(n5449));
   INV_X1 U1245 (.ZN(n721), 
	.A(n735));
   OAI211_X1 U1246 (.ZN(n735), 
	.C2(n321), 
	.C1(n5624), 
	.B(n737), 
	.A(n736));
   AOI222_X1 U1247 (.ZN(n737), 
	.C2(n739), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[4] ), 
	.A2(n738), 
	.A1(FE_OFN91_n285));
   INV_X1 U1248 (.ZN(n739), 
	.A(n5683));
   AOI22_X1 U1249 (.ZN(n736), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[4] ), 
	.A2(n6194), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1250 (.ZN(n3654), 
	.B2(n2691), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n740));
   OAI221_X1 U1251 (.ZN(n3655), 
	.C2(n71), 
	.C1(n86), 
	.B2(n69), 
	.B1(FE_OFN197_n741), 
	.A(n742));
   NAND2_X1 U1252 (.ZN(n742), 
	.A2(FE_OFN8_n73), 
	.A1(\UUT/Mpath/the_mult/x_operand2 [3]));
   OAI222_X1 U1253 (.ZN(n3656), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N78 ), 
	.B2(n300), 
	.B1(FE_OFN197_n741), 
	.A2(n123), 
	.A1(n86));
   INV_X1 U1254 (.ZN(n86), 
	.A(n743));
   OAI222_X1 U1255 (.ZN(n743), 
	.C2(n132), 
	.C1(n5451), 
	.B2(n131), 
	.B1(n745), 
	.A2(n129), 
	.A1(n744));
   OAI221_X1 U1256 (.ZN(n3657), 
	.C2(n135), 
	.C1(n5684), 
	.B2(n746), 
	.B1(n133), 
	.A(n747));
   AOI22_X1 U1257 (.ZN(n747), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [35]), 
	.A2(n748), 
	.A1(n137));
   OAI221_X1 U1258 (.ZN(n3658), 
	.C2(n142), 
	.C1(n5626), 
	.B2(n749), 
	.B1(n140), 
	.A(n750));
   AOI22_X1 U1259 (.ZN(n750), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [3]), 
	.A2(n748), 
	.A1(n144));
   INV_X1 U1260 (.ZN(n748), 
	.A(n5627));
   OAI22_X1 U1261 (.ZN(n3659), 
	.B2(net54871), 
	.B1(n5627), 
	.A2(n751), 
	.A1(net54953));
   OAI221_X1 U1262 (.ZN(n3660), 
	.C2(n751), 
	.C1(n147), 
	.B2(n310), 
	.B1(n744), 
	.A(n752));
   AOI22_X1 U1263 (.ZN(n752), 
	.B2(n754), 
	.B1(FE_OFN6_n314), 
	.A2(n753), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1264 (.ZN(n751), 
	.A(FE_OFN165_UUT_Mpath_the_mult_x_operand1_3_));
   OAI221_X1 U1265 (.ZN(n3661), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N77 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n744), 
	.A(n755));
   AOI22_X1 U1266 (.ZN(n755), 
	.B2(n754), 
	.B1(FE_OFN4_n319), 
	.A2(n753), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1267 (.ZN(n3662), 
	.B2(n219), 
	.B1(n745), 
	.A2(n6407), 
	.A1(n5387));
   OAI22_X1 U1268 (.ZN(n3663), 
	.B2(n221), 
	.B1(n745), 
	.A2(n6410), 
	.A1(n5355));
   OAI22_X1 U1269 (.ZN(n3664), 
	.B2(n223), 
	.B1(n745), 
	.A2(n6401), 
	.A1(n5323));
   OAI22_X1 U1270 (.ZN(n3665), 
	.B2(n225), 
	.B1(n745), 
	.A2(n6406), 
	.A1(n5291));
   OAI22_X1 U1271 (.ZN(n3666), 
	.B2(n227), 
	.B1(n745), 
	.A2(n6399), 
	.A1(n5259));
   OAI22_X1 U1272 (.ZN(n3667), 
	.B2(n229), 
	.B1(n745), 
	.A2(n6404), 
	.A1(n5227));
   OAI22_X1 U1273 (.ZN(n3668), 
	.B2(n231), 
	.B1(n745), 
	.A2(n6398), 
	.A1(n5195));
   OAI22_X1 U1274 (.ZN(n3669), 
	.B2(n233), 
	.B1(n745), 
	.A2(n6396), 
	.A1(n5163));
   OAI22_X1 U1275 (.ZN(n3670), 
	.B2(n235), 
	.B1(n745), 
	.A2(n6393), 
	.A1(n5131));
   OAI22_X1 U1276 (.ZN(n3671), 
	.B2(n237), 
	.B1(n745), 
	.A2(n6391), 
	.A1(n5099));
   OAI22_X1 U1277 (.ZN(n3672), 
	.B2(n239), 
	.B1(n745), 
	.A2(n6390), 
	.A1(n5067));
   OAI22_X1 U1278 (.ZN(n3673), 
	.B2(n241), 
	.B1(n745), 
	.A2(n6388), 
	.A1(n5035));
   OAI22_X1 U1279 (.ZN(n3674), 
	.B2(n243), 
	.B1(n745), 
	.A2(n6385), 
	.A1(n5003));
   OAI22_X1 U1280 (.ZN(n3675), 
	.B2(n245), 
	.B1(n745), 
	.A2(n6383), 
	.A1(n4971));
   OAI22_X1 U1281 (.ZN(n3676), 
	.B2(n247), 
	.B1(n745), 
	.A2(n6382), 
	.A1(n4939));
   OAI22_X1 U1282 (.ZN(n3677), 
	.B2(n249), 
	.B1(n745), 
	.A2(n6380), 
	.A1(n4907));
   OAI22_X1 U1283 (.ZN(n3678), 
	.B2(n251), 
	.B1(n745), 
	.A2(n6384), 
	.A1(n4875));
   OAI22_X1 U1284 (.ZN(n3679), 
	.B2(n253), 
	.B1(n745), 
	.A2(n6381), 
	.A1(n4843));
   OAI22_X1 U1285 (.ZN(n3680), 
	.B2(n255), 
	.B1(n745), 
	.A2(n6387), 
	.A1(n4811));
   OAI22_X1 U1286 (.ZN(n3681), 
	.B2(n257), 
	.B1(n745), 
	.A2(n6386), 
	.A1(n4779));
   OAI22_X1 U1287 (.ZN(n3682), 
	.B2(n259), 
	.B1(n745), 
	.A2(n6392), 
	.A1(n4747));
   OAI22_X1 U1288 (.ZN(n3683), 
	.B2(n261), 
	.B1(n745), 
	.A2(n6394), 
	.A1(n4715));
   OAI22_X1 U1289 (.ZN(n3684), 
	.B2(n263), 
	.B1(n745), 
	.A2(n6389), 
	.A1(n4683));
   OAI22_X1 U1290 (.ZN(n3685), 
	.B2(n265), 
	.B1(n745), 
	.A2(n6395), 
	.A1(n4651));
   OAI22_X1 U1291 (.ZN(n3686), 
	.B2(n267), 
	.B1(n745), 
	.A2(n6400), 
	.A1(n4619));
   OAI22_X1 U1292 (.ZN(n3687), 
	.B2(n269), 
	.B1(n745), 
	.A2(n6402), 
	.A1(n4587));
   OAI22_X1 U1293 (.ZN(n3688), 
	.B2(n271), 
	.B1(n745), 
	.A2(n6397), 
	.A1(n4555));
   OAI22_X1 U1294 (.ZN(n3689), 
	.B2(n273), 
	.B1(n745), 
	.A2(n6403), 
	.A1(n4523));
   OAI22_X1 U1295 (.ZN(n3690), 
	.B2(n275), 
	.B1(n745), 
	.A2(n6408), 
	.A1(n4491));
   OAI22_X1 U1296 (.ZN(n3691), 
	.B2(n277), 
	.B1(n745), 
	.A2(n6405), 
	.A1(n4459));
   OAI22_X1 U1297 (.ZN(n3692), 
	.B2(n279), 
	.B1(n745), 
	.A2(n6411), 
	.A1(n4427));
   OAI211_X1 U1299 (.ZN(n754), 
	.C2(n5452), 
	.C1(n5710), 
	.B(n757), 
	.A(n756));
   AOI222_X1 U1300 (.ZN(n757), 
	.C2(n686), 
	.C1(n5817), 
	.B2(n589), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5812));
   INV_X1 U1301 (.ZN(n589), 
	.A(n5819));
   AOI22_X1 U1302 (.ZN(n756), 
	.B2(n688), 
	.B1(n5814), 
	.A2(n687), 
	.A1(n5818));
   OAI22_X1 U1303 (.ZN(n3693), 
	.B2(n744), 
	.B1(FE_OFN12_net54953), 
	.A2(net54883), 
	.A1(n5452));
   INV_X1 U1304 (.ZN(n744), 
	.A(n758));
   OAI211_X1 U1305 (.ZN(n758), 
	.C2(n321), 
	.C1(n5626), 
	.B(n760), 
	.A(n759));
   AOI222_X1 U1306 (.ZN(n760), 
	.C2(n762), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[3] ), 
	.A2(n761), 
	.A1(FE_OFN91_n285));
   INV_X1 U1307 (.ZN(n762), 
	.A(n5684));
   AOI22_X1 U1308 (.ZN(n759), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[3] ), 
	.A2(n6195), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1309 (.ZN(n3694), 
	.B2(n2694), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n763));
   OAI221_X1 U1310 (.ZN(n3695), 
	.C2(n71), 
	.C1(n85), 
	.B2(n69), 
	.B1(FE_OFN196_n764), 
	.A(n765));
   NAND2_X1 U1311 (.ZN(n765), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN167_UUT_Mpath_the_mult_x_operand2_2_));
   OAI222_X1 U1312 (.ZN(n3696), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N80 ), 
	.B2(n300), 
	.B1(FE_OFN196_n764), 
	.A2(n123), 
	.A1(n85));
   INV_X1 U1313 (.ZN(n85), 
	.A(n766));
   OAI222_X1 U1314 (.ZN(n766), 
	.C2(n132), 
	.C1(n5460), 
	.B2(n131), 
	.B1(n768), 
	.A2(n129), 
	.A1(n767));
   OAI221_X1 U1315 (.ZN(n3697), 
	.C2(n135), 
	.C1(n5687), 
	.B2(n769), 
	.B1(n133), 
	.A(n770));
   AOI22_X1 U1316 (.ZN(n770), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [34]), 
	.A2(n771), 
	.A1(n137));
   OAI221_X1 U1317 (.ZN(n3698), 
	.C2(n142), 
	.C1(n5632), 
	.B2(n772), 
	.B1(n140), 
	.A(n773));
   AOI22_X1 U1318 (.ZN(n773), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [2]), 
	.A2(n771), 
	.A1(n144));
   INV_X1 U1319 (.ZN(n771), 
	.A(n5633));
   OAI22_X1 U1320 (.ZN(n3699), 
	.B2(net54871), 
	.B1(n5633), 
	.A2(n774), 
	.A1(net54953));
   OAI221_X1 U1321 (.ZN(n3700), 
	.C2(n774), 
	.C1(n147), 
	.B2(n310), 
	.B1(n767), 
	.A(n775));
   AOI22_X1 U1322 (.ZN(n775), 
	.B2(n777), 
	.B1(FE_OFN6_n314), 
	.A2(n776), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1323 (.ZN(n774), 
	.A(\UUT/Mpath/the_mult/x_operand1[2] ));
   OAI221_X1 U1324 (.ZN(n3701), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N79 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n767), 
	.A(n778));
   AOI22_X1 U1325 (.ZN(n778), 
	.B2(n777), 
	.B1(FE_OFN4_n319), 
	.A2(n776), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1326 (.ZN(n3702), 
	.B2(n219), 
	.B1(n768), 
	.A2(n6407), 
	.A1(n5390));
   OAI22_X1 U1327 (.ZN(n3703), 
	.B2(n221), 
	.B1(n768), 
	.A2(n6410), 
	.A1(n5358));
   OAI22_X1 U1328 (.ZN(n3704), 
	.B2(n223), 
	.B1(n768), 
	.A2(n6401), 
	.A1(n5326));
   OAI22_X1 U1329 (.ZN(n3705), 
	.B2(n225), 
	.B1(n768), 
	.A2(n6406), 
	.A1(n5294));
   OAI22_X1 U1330 (.ZN(n3706), 
	.B2(n227), 
	.B1(n768), 
	.A2(n6399), 
	.A1(n5262));
   OAI22_X1 U1331 (.ZN(n3707), 
	.B2(n229), 
	.B1(n768), 
	.A2(n6404), 
	.A1(n5230));
   OAI22_X1 U1332 (.ZN(n3708), 
	.B2(n231), 
	.B1(n768), 
	.A2(n6398), 
	.A1(n5198));
   OAI22_X1 U1333 (.ZN(n3709), 
	.B2(n233), 
	.B1(n768), 
	.A2(n6396), 
	.A1(n5166));
   OAI22_X1 U1334 (.ZN(n3710), 
	.B2(n235), 
	.B1(n768), 
	.A2(n6393), 
	.A1(n5134));
   OAI22_X1 U1335 (.ZN(n3711), 
	.B2(n237), 
	.B1(n768), 
	.A2(n6391), 
	.A1(n5102));
   OAI22_X1 U1336 (.ZN(n3712), 
	.B2(n239), 
	.B1(n768), 
	.A2(n6390), 
	.A1(n5070));
   OAI22_X1 U1337 (.ZN(n3713), 
	.B2(n241), 
	.B1(n768), 
	.A2(n6388), 
	.A1(n5038));
   OAI22_X1 U1338 (.ZN(n3714), 
	.B2(n243), 
	.B1(n768), 
	.A2(n6385), 
	.A1(n5006));
   OAI22_X1 U1339 (.ZN(n3715), 
	.B2(n245), 
	.B1(n768), 
	.A2(n6383), 
	.A1(n4974));
   OAI22_X1 U1340 (.ZN(n3716), 
	.B2(n247), 
	.B1(n768), 
	.A2(n6382), 
	.A1(n4942));
   OAI22_X1 U1341 (.ZN(n3717), 
	.B2(n249), 
	.B1(n768), 
	.A2(n6380), 
	.A1(n4910));
   OAI22_X1 U1342 (.ZN(n3718), 
	.B2(n251), 
	.B1(n768), 
	.A2(n6384), 
	.A1(n4878));
   OAI22_X1 U1343 (.ZN(n3719), 
	.B2(n253), 
	.B1(n768), 
	.A2(n6381), 
	.A1(n4846));
   OAI22_X1 U1344 (.ZN(n3720), 
	.B2(n255), 
	.B1(n768), 
	.A2(n6387), 
	.A1(n4814));
   OAI22_X1 U1345 (.ZN(n3721), 
	.B2(n257), 
	.B1(n768), 
	.A2(n6386), 
	.A1(n4782));
   OAI22_X1 U1346 (.ZN(n3722), 
	.B2(n259), 
	.B1(n768), 
	.A2(n6392), 
	.A1(n4750));
   OAI22_X1 U1347 (.ZN(n3723), 
	.B2(n261), 
	.B1(n768), 
	.A2(n6394), 
	.A1(n4718));
   OAI22_X1 U1348 (.ZN(n3724), 
	.B2(n263), 
	.B1(n768), 
	.A2(n6389), 
	.A1(n4686));
   OAI22_X1 U1349 (.ZN(n3725), 
	.B2(n265), 
	.B1(n768), 
	.A2(n6395), 
	.A1(n4654));
   OAI22_X1 U1350 (.ZN(n3726), 
	.B2(n267), 
	.B1(n768), 
	.A2(n6400), 
	.A1(n4622));
   OAI22_X1 U1351 (.ZN(n3727), 
	.B2(n269), 
	.B1(n768), 
	.A2(n6402), 
	.A1(n4590));
   OAI22_X1 U1352 (.ZN(n3728), 
	.B2(n271), 
	.B1(n768), 
	.A2(n6397), 
	.A1(n4558));
   OAI22_X1 U1353 (.ZN(n3729), 
	.B2(n273), 
	.B1(n768), 
	.A2(n6403), 
	.A1(n4526));
   OAI22_X1 U1354 (.ZN(n3730), 
	.B2(n275), 
	.B1(n768), 
	.A2(n6408), 
	.A1(n4494));
   OAI22_X1 U1355 (.ZN(n3731), 
	.B2(n277), 
	.B1(n768), 
	.A2(n6405), 
	.A1(n4462));
   OAI22_X1 U1356 (.ZN(n3732), 
	.B2(n279), 
	.B1(n768), 
	.A2(n6411), 
	.A1(n4430));
   OAI211_X1 U1358 (.ZN(n777), 
	.C2(n5461), 
	.C1(n5710), 
	.B(n780), 
	.A(n779));
   AOI222_X1 U1359 (.ZN(n780), 
	.C2(n686), 
	.C1(n5843), 
	.B2(n781), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5838));
   AOI22_X1 U1360 (.ZN(n779), 
	.B2(n688), 
	.B1(n5840), 
	.A2(n687), 
	.A1(n5844));
   OAI22_X1 U1361 (.ZN(n3733), 
	.B2(n767), 
	.B1(FE_OFN12_net54953), 
	.A2(net54885), 
	.A1(n5461));
   INV_X1 U1362 (.ZN(n767), 
	.A(n782));
   OAI211_X1 U1363 (.ZN(n782), 
	.C2(n321), 
	.C1(n5632), 
	.B(n784), 
	.A(n783));
   AOI222_X1 U1364 (.ZN(n784), 
	.C2(n786), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[2] ), 
	.A2(n785), 
	.A1(FE_OFN91_n285));
   INV_X1 U1365 (.ZN(n786), 
	.A(n5687));
   AOI22_X1 U1366 (.ZN(n783), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[2] ), 
	.A2(n6202), 
	.A1(FE_OFN89_n290));
   OAI221_X1 U1367 (.ZN(n3734), 
	.C2(n71), 
	.C1(n84), 
	.B2(n69), 
	.B1(n787), 
	.A(n788));
   NAND2_X1 U1368 (.ZN(n788), 
	.A2(FE_OFN8_n73), 
	.A1(FE_OFN170_UUT_Mpath_the_mult_x_operand2_1_));
   NAND2_X2 U1370 (.ZN(n69), 
	.A2(n789), 
	.A1(n147));
   OAI221_X1 U1373 (.ZN(n3736), 
	.C2(n135), 
	.C1(n5698), 
	.B2(n791), 
	.B1(n133), 
	.A(n792));
   AOI22_X1 U1374 (.ZN(n792), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [33]), 
	.A2(n793), 
	.A1(n137));
   OAI221_X1 U1375 (.ZN(n3737), 
	.C2(n142), 
	.C1(n5654), 
	.B2(n794), 
	.B1(n140), 
	.A(n795));
   AOI22_X1 U1376 (.ZN(n795), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [1]), 
	.A2(n793), 
	.A1(n144));
   INV_X1 U1377 (.ZN(n793), 
	.A(n5655));
   OAI22_X1 U1378 (.ZN(n3738), 
	.B2(net54871), 
	.B1(n5655), 
	.A2(n796), 
	.A1(net54953));
   OAI221_X1 U1379 (.ZN(n3739), 
	.C2(n796), 
	.C1(n147), 
	.B2(n310), 
	.B1(n797), 
	.A(n798));
   AOI22_X1 U1380 (.ZN(n798), 
	.B2(n800), 
	.B1(FE_OFN6_n314), 
	.A2(n799), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1381 (.ZN(n796), 
	.A(FE_OFN171_UUT_Mpath_the_mult_x_operand1_1_));
   OAI221_X1 U1382 (.ZN(n3740), 
	.C2(net54885), 
	.C1(\UUT/Mpath/the_alu/N81 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n797), 
	.A(n801));
   AOI22_X1 U1383 (.ZN(n801), 
	.B2(n800), 
	.B1(FE_OFN4_n319), 
	.A2(n799), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1384 (.ZN(n3741), 
	.B2(n219), 
	.B1(n802), 
	.A2(n6407), 
	.A1(n5401));
   OAI22_X1 U1385 (.ZN(n3742), 
	.B2(n221), 
	.B1(n802), 
	.A2(n6410), 
	.A1(n5369));
   OAI22_X1 U1386 (.ZN(n3743), 
	.B2(n223), 
	.B1(n802), 
	.A2(n6401), 
	.A1(n5337));
   OAI22_X1 U1387 (.ZN(n3744), 
	.B2(n225), 
	.B1(n802), 
	.A2(n6406), 
	.A1(n5305));
   OAI22_X1 U1388 (.ZN(n3745), 
	.B2(n227), 
	.B1(n802), 
	.A2(n6399), 
	.A1(n5273));
   OAI22_X1 U1389 (.ZN(n3746), 
	.B2(n229), 
	.B1(n802), 
	.A2(n6404), 
	.A1(n5241));
   OAI22_X1 U1390 (.ZN(n3747), 
	.B2(n231), 
	.B1(n802), 
	.A2(n6398), 
	.A1(n5209));
   OAI22_X1 U1391 (.ZN(n3748), 
	.B2(n233), 
	.B1(n802), 
	.A2(n6396), 
	.A1(n5177));
   OAI22_X1 U1392 (.ZN(n3749), 
	.B2(n235), 
	.B1(n802), 
	.A2(n6393), 
	.A1(n5145));
   OAI22_X1 U1393 (.ZN(n3750), 
	.B2(n237), 
	.B1(n802), 
	.A2(n6391), 
	.A1(n5113));
   OAI22_X1 U1394 (.ZN(n3751), 
	.B2(n239), 
	.B1(n802), 
	.A2(n6390), 
	.A1(n5081));
   OAI22_X1 U1395 (.ZN(n3752), 
	.B2(n241), 
	.B1(n802), 
	.A2(n6388), 
	.A1(n5049));
   OAI22_X1 U1396 (.ZN(n3753), 
	.B2(n243), 
	.B1(n802), 
	.A2(n6385), 
	.A1(n5017));
   OAI22_X1 U1397 (.ZN(n3754), 
	.B2(n245), 
	.B1(n802), 
	.A2(n6383), 
	.A1(n4985));
   OAI22_X1 U1398 (.ZN(n3755), 
	.B2(n247), 
	.B1(n802), 
	.A2(n6382), 
	.A1(n4953));
   OAI22_X1 U1399 (.ZN(n3756), 
	.B2(n249), 
	.B1(n802), 
	.A2(n6380), 
	.A1(n4921));
   OAI22_X1 U1400 (.ZN(n3757), 
	.B2(n251), 
	.B1(n802), 
	.A2(n6384), 
	.A1(n4889));
   OAI22_X1 U1401 (.ZN(n3758), 
	.B2(n253), 
	.B1(n802), 
	.A2(n6381), 
	.A1(n4857));
   OAI22_X1 U1402 (.ZN(n3759), 
	.B2(n255), 
	.B1(n802), 
	.A2(n6387), 
	.A1(n4825));
   OAI22_X1 U1403 (.ZN(n3760), 
	.B2(n257), 
	.B1(n802), 
	.A2(n6386), 
	.A1(n4793));
   OAI22_X1 U1404 (.ZN(n3761), 
	.B2(n259), 
	.B1(n802), 
	.A2(n6392), 
	.A1(n4761));
   OAI22_X1 U1405 (.ZN(n3762), 
	.B2(n261), 
	.B1(n802), 
	.A2(n6394), 
	.A1(n4729));
   OAI22_X1 U1406 (.ZN(n3763), 
	.B2(n263), 
	.B1(n802), 
	.A2(n6389), 
	.A1(n4697));
   OAI22_X1 U1407 (.ZN(n3764), 
	.B2(n265), 
	.B1(n802), 
	.A2(n6395), 
	.A1(n4665));
   OAI22_X1 U1408 (.ZN(n3765), 
	.B2(n267), 
	.B1(n802), 
	.A2(n6400), 
	.A1(n4633));
   OAI22_X1 U1409 (.ZN(n3766), 
	.B2(n269), 
	.B1(n802), 
	.A2(n6402), 
	.A1(n4601));
   OAI22_X1 U1410 (.ZN(n3767), 
	.B2(n271), 
	.B1(n802), 
	.A2(n6397), 
	.A1(n4569));
   OAI22_X1 U1411 (.ZN(n3768), 
	.B2(n273), 
	.B1(n802), 
	.A2(n6403), 
	.A1(n4537));
   OAI22_X1 U1412 (.ZN(n3769), 
	.B2(n275), 
	.B1(n802), 
	.A2(n6408), 
	.A1(n4505));
   OAI22_X1 U1413 (.ZN(n3770), 
	.B2(n277), 
	.B1(n802), 
	.A2(n6405), 
	.A1(n4473));
   OAI22_X1 U1414 (.ZN(n3771), 
	.B2(n279), 
	.B1(n802), 
	.A2(n6411), 
	.A1(n4441));
   OAI221_X1 U1415 (.ZN(n3772), 
	.C2(n135), 
	.C1(n5694), 
	.B2(n803), 
	.B1(n133), 
	.A(n804));
   AOI22_X1 U1416 (.ZN(n804), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [55]), 
	.A2(n805), 
	.A1(n137));
   OAI221_X1 U1417 (.ZN(n3773), 
	.C2(n142), 
	.C1(n5646), 
	.B2(n806), 
	.B1(n140), 
	.A(n807));
   AOI22_X1 U1418 (.ZN(n807), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [23]), 
	.A2(n805), 
	.A1(n144));
   INV_X1 U1419 (.ZN(n805), 
	.A(n5647));
   OAI22_X1 U1420 (.ZN(n3774), 
	.B2(net54871), 
	.B1(n5647), 
	.A2(n808), 
	.A1(FE_OFN11_net54953));
   OAI221_X1 U1421 (.ZN(n3775), 
	.C2(n808), 
	.C1(n147), 
	.B2(n310), 
	.B1(n809), 
	.A(n810));
   AOI22_X1 U1422 (.ZN(n810), 
	.B2(n812), 
	.B1(FE_OFN6_n314), 
	.A2(n811), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U1423 (.ZN(n808), 
	.A(FE_OFN173_UUT_Mpath_the_mult_x_operand1_23_));
   OAI221_X1 U1424 (.ZN(n3776), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N37 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n809), 
	.A(n813));
   AOI22_X1 U1425 (.ZN(n813), 
	.B2(n812), 
	.B1(FE_OFN4_n319), 
	.A2(n811), 
	.A1(FE_OFN5_n318));
   OAI22_X1 U1426 (.ZN(n3777), 
	.B2(n219), 
	.B1(n814), 
	.A2(n6407), 
	.A1(n5397));
   OAI22_X1 U1427 (.ZN(n3778), 
	.B2(n221), 
	.B1(n814), 
	.A2(n6410), 
	.A1(n5365));
   OAI22_X1 U1428 (.ZN(n3779), 
	.B2(n223), 
	.B1(n814), 
	.A2(n6401), 
	.A1(n5333));
   OAI22_X1 U1429 (.ZN(n3780), 
	.B2(n225), 
	.B1(n814), 
	.A2(n6406), 
	.A1(n5301));
   OAI22_X1 U1430 (.ZN(n3781), 
	.B2(n227), 
	.B1(n814), 
	.A2(n6399), 
	.A1(n5269));
   OAI22_X1 U1431 (.ZN(n3782), 
	.B2(n229), 
	.B1(n814), 
	.A2(n6404), 
	.A1(n5237));
   OAI22_X1 U1432 (.ZN(n3783), 
	.B2(n231), 
	.B1(n814), 
	.A2(n6398), 
	.A1(n5205));
   OAI22_X1 U1433 (.ZN(n3784), 
	.B2(n233), 
	.B1(n814), 
	.A2(n6396), 
	.A1(n5173));
   OAI22_X1 U1434 (.ZN(n3785), 
	.B2(n235), 
	.B1(n814), 
	.A2(n6393), 
	.A1(n5141));
   OAI22_X1 U1435 (.ZN(n3786), 
	.B2(n237), 
	.B1(n814), 
	.A2(n6391), 
	.A1(n5109));
   OAI22_X1 U1436 (.ZN(n3787), 
	.B2(n239), 
	.B1(n814), 
	.A2(n6390), 
	.A1(n5077));
   OAI22_X1 U1437 (.ZN(n3788), 
	.B2(n241), 
	.B1(n814), 
	.A2(n6388), 
	.A1(n5045));
   OAI22_X1 U1438 (.ZN(n3789), 
	.B2(n243), 
	.B1(n814), 
	.A2(n6385), 
	.A1(n5013));
   OAI22_X1 U1439 (.ZN(n3790), 
	.B2(n245), 
	.B1(n814), 
	.A2(n6383), 
	.A1(n4981));
   OAI22_X1 U1440 (.ZN(n3791), 
	.B2(n247), 
	.B1(n814), 
	.A2(n6382), 
	.A1(n4949));
   OAI22_X1 U1441 (.ZN(n3792), 
	.B2(n249), 
	.B1(n814), 
	.A2(n6380), 
	.A1(n4917));
   OAI22_X1 U1442 (.ZN(n3793), 
	.B2(n251), 
	.B1(n814), 
	.A2(n6384), 
	.A1(n4885));
   OAI22_X1 U1443 (.ZN(n3794), 
	.B2(n253), 
	.B1(n814), 
	.A2(n6381), 
	.A1(n4853));
   OAI22_X1 U1444 (.ZN(n3795), 
	.B2(n255), 
	.B1(n814), 
	.A2(n6387), 
	.A1(n4821));
   OAI22_X1 U1445 (.ZN(n3796), 
	.B2(n257), 
	.B1(n814), 
	.A2(n6386), 
	.A1(n4789));
   OAI22_X1 U1446 (.ZN(n3797), 
	.B2(n259), 
	.B1(n814), 
	.A2(n6392), 
	.A1(n4757));
   OAI22_X1 U1447 (.ZN(n3798), 
	.B2(n261), 
	.B1(n814), 
	.A2(n6394), 
	.A1(n4725));
   OAI22_X1 U1448 (.ZN(n3799), 
	.B2(n263), 
	.B1(n814), 
	.A2(n6389), 
	.A1(n4693));
   OAI22_X1 U1449 (.ZN(n3800), 
	.B2(n265), 
	.B1(n814), 
	.A2(n6395), 
	.A1(n4661));
   OAI22_X1 U1450 (.ZN(n3801), 
	.B2(n267), 
	.B1(n814), 
	.A2(n6400), 
	.A1(n4629));
   OAI22_X1 U1451 (.ZN(n3802), 
	.B2(n269), 
	.B1(n814), 
	.A2(n6402), 
	.A1(n4597));
   OAI22_X1 U1452 (.ZN(n3803), 
	.B2(n271), 
	.B1(n814), 
	.A2(n6397), 
	.A1(n4565));
   OAI22_X1 U1453 (.ZN(n3804), 
	.B2(n273), 
	.B1(n814), 
	.A2(n6403), 
	.A1(n4533));
   OAI22_X1 U1454 (.ZN(n3805), 
	.B2(n275), 
	.B1(n814), 
	.A2(n6408), 
	.A1(n4501));
   OAI22_X1 U1455 (.ZN(n3806), 
	.B2(n277), 
	.B1(n814), 
	.A2(n6405), 
	.A1(n4469));
   OAI22_X1 U1456 (.ZN(n3807), 
	.B2(n279), 
	.B1(n814), 
	.A2(n6411), 
	.A1(n4437));
   OAI22_X1 U1457 (.ZN(n3808), 
	.B2(\UUT/Mpath/the_memhandle/N239 ), 
	.B1(net54867), 
	.A2(n815), 
	.A1(FE_OFN11_net54953));
   INV_X1 U1458 (.ZN(n815), 
	.A(\UUT/daddr_out [1]));
   OAI222_X1 U1459 (.ZN(n3809), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N82 ), 
	.B2(n300), 
	.B1(n787), 
	.A2(n123), 
	.A1(n84));
   INV_X1 U1460 (.ZN(n787), 
	.A(\UUT/break_code[1] ));
   INV_X1 U1461 (.ZN(n84), 
	.A(n816));
   OAI222_X1 U1462 (.ZN(n816), 
	.C2(n132), 
	.C1(n5493), 
	.B2(n131), 
	.B1(n802), 
	.A2(n129), 
	.A1(n797));
   OAI211_X1 U1464 (.ZN(n800), 
	.C2(n5494), 
	.C1(n5710), 
	.B(n818), 
	.A(n817));
   AOI222_X1 U1465 (.ZN(n818), 
	.C2(n686), 
	.C1(n5922), 
	.B2(n624), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5712));
   INV_X1 U1466 (.ZN(n624), 
	.A(n5921));
   AOI22_X1 U1467 (.ZN(n817), 
	.B2(n688), 
	.B1(n5918), 
	.A2(n687), 
	.A1(n5923));
   OAI22_X1 U1468 (.ZN(n3810), 
	.B2(n797), 
	.B1(FE_OFN12_net54953), 
	.A2(net54877), 
	.A1(n5494));
   INV_X1 U1469 (.ZN(n797), 
	.A(n819));
   OAI211_X1 U1470 (.ZN(n819), 
	.C2(n321), 
	.C1(n5654), 
	.B(n821), 
	.A(n820));
   AOI222_X1 U1471 (.ZN(n821), 
	.C2(n823), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[1] ), 
	.A2(n822), 
	.A1(FE_OFN91_n285));
   INV_X1 U1472 (.ZN(n823), 
	.A(n5698));
   AOI22_X1 U1473 (.ZN(n820), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[1] ), 
	.A2(\UUT/daddr_out [1]), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U1474 (.ZN(n3811), 
	.B2(n201), 
	.B1(net54953), 
	.A2(net54877), 
	.A1(\UUT/Mpath/the_alu/N33 ));
   INV_X1 U1475 (.ZN(n201), 
	.A(n824));
   OAI222_X1 U1476 (.ZN(n824), 
	.C2(n5420), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN21_n193), 
	.B1(n5528), 
	.A2(n194), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1477 (.ZN(n3812), 
	.B2(n219), 
	.B1(n194), 
	.A2(n6407), 
	.A1(n5395));
   OAI22_X1 U1478 (.ZN(n3813), 
	.B2(n221), 
	.B1(n194), 
	.A2(n6410), 
	.A1(n5363));
   OAI22_X1 U1479 (.ZN(n3814), 
	.B2(n223), 
	.B1(n194), 
	.A2(n6401), 
	.A1(n5331));
   OAI22_X1 U1480 (.ZN(n3815), 
	.B2(n225), 
	.B1(n194), 
	.A2(n6406), 
	.A1(n5299));
   OAI22_X1 U1481 (.ZN(n3816), 
	.B2(n227), 
	.B1(n194), 
	.A2(n6399), 
	.A1(n5267));
   OAI22_X1 U1482 (.ZN(n3817), 
	.B2(n229), 
	.B1(n194), 
	.A2(n6404), 
	.A1(n5235));
   OAI22_X1 U1483 (.ZN(n3818), 
	.B2(n231), 
	.B1(n194), 
	.A2(n6398), 
	.A1(n5203));
   OAI22_X1 U1484 (.ZN(n3819), 
	.B2(n233), 
	.B1(n194), 
	.A2(n6396), 
	.A1(n5171));
   OAI22_X1 U1485 (.ZN(n3820), 
	.B2(n235), 
	.B1(n194), 
	.A2(n6393), 
	.A1(n5139));
   OAI22_X1 U1486 (.ZN(n3821), 
	.B2(n237), 
	.B1(n194), 
	.A2(n6391), 
	.A1(n5107));
   OAI22_X1 U1487 (.ZN(n3822), 
	.B2(n239), 
	.B1(n194), 
	.A2(n6390), 
	.A1(n5075));
   OAI22_X1 U1488 (.ZN(n3823), 
	.B2(n241), 
	.B1(n194), 
	.A2(n6388), 
	.A1(n5043));
   OAI22_X1 U1489 (.ZN(n3824), 
	.B2(n243), 
	.B1(n194), 
	.A2(n6385), 
	.A1(n5011));
   OAI22_X1 U1490 (.ZN(n3825), 
	.B2(n245), 
	.B1(n194), 
	.A2(n6383), 
	.A1(n4979));
   OAI22_X1 U1491 (.ZN(n3826), 
	.B2(n247), 
	.B1(n194), 
	.A2(n6382), 
	.A1(n4947));
   OAI22_X1 U1492 (.ZN(n3827), 
	.B2(n249), 
	.B1(n194), 
	.A2(n6380), 
	.A1(n4915));
   OAI22_X1 U1493 (.ZN(n3828), 
	.B2(n251), 
	.B1(n194), 
	.A2(n6384), 
	.A1(n4883));
   OAI22_X1 U1494 (.ZN(n3829), 
	.B2(n253), 
	.B1(n194), 
	.A2(n6381), 
	.A1(n4851));
   OAI22_X1 U1495 (.ZN(n3830), 
	.B2(n255), 
	.B1(n194), 
	.A2(n6387), 
	.A1(n4819));
   OAI22_X1 U1496 (.ZN(n3831), 
	.B2(n257), 
	.B1(n194), 
	.A2(n6386), 
	.A1(n4787));
   OAI22_X1 U1497 (.ZN(n3832), 
	.B2(n259), 
	.B1(n194), 
	.A2(n6392), 
	.A1(n4755));
   OAI22_X1 U1498 (.ZN(n3833), 
	.B2(n261), 
	.B1(n194), 
	.A2(n6394), 
	.A1(n4723));
   OAI22_X1 U1499 (.ZN(n3834), 
	.B2(n263), 
	.B1(n194), 
	.A2(n6389), 
	.A1(n4691));
   OAI22_X1 U1500 (.ZN(n3835), 
	.B2(n265), 
	.B1(n194), 
	.A2(n6395), 
	.A1(n4659));
   OAI22_X1 U1501 (.ZN(n3836), 
	.B2(n267), 
	.B1(n194), 
	.A2(n6400), 
	.A1(n4627));
   OAI22_X1 U1502 (.ZN(n3837), 
	.B2(n269), 
	.B1(n194), 
	.A2(n6402), 
	.A1(n4595));
   OAI22_X1 U1503 (.ZN(n3838), 
	.B2(n271), 
	.B1(n194), 
	.A2(n6397), 
	.A1(n4563));
   OAI22_X1 U1504 (.ZN(n3839), 
	.B2(n273), 
	.B1(n194), 
	.A2(n6403), 
	.A1(n4531));
   OAI22_X1 U1505 (.ZN(n3840), 
	.B2(n275), 
	.B1(n194), 
	.A2(n6408), 
	.A1(n4499));
   OAI22_X1 U1506 (.ZN(n3841), 
	.B2(n277), 
	.B1(n194), 
	.A2(n6405), 
	.A1(n4467));
   OAI22_X1 U1507 (.ZN(n3842), 
	.B2(n279), 
	.B1(n194), 
	.A2(n6411), 
	.A1(n4435));
   OAI22_X1 U1510 (.ZN(n3843), 
	.B2(FE_OFN21_n193), 
	.B1(FE_OFN11_net54953), 
	.A2(net54877), 
	.A1(n5476));
   AOI221_X1 U1511 (.ZN(n193), 
	.C2(FE_OFN91_n285), 
	.C1(n5598), 
	.B2(n284), 
	.B1(n826), 
	.A(n827));
   INV_X1 U1512 (.ZN(n827), 
	.A(n828));
   AOI222_X1 U1513 (.ZN(n828), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[25] ), 
	.B2(n5599), 
	.B1(FE_OFN89_n290), 
	.A2(n829), 
	.A1(n288));
   INV_X1 U1514 (.ZN(n829), 
	.A(n5642));
   INV_X1 U1515 (.ZN(n826), 
	.A(n5692));
   OAI22_X1 U1516 (.ZN(n3844), 
	.B2(n188), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N31 ));
   INV_X1 U1517 (.ZN(n188), 
	.A(n830));
   OAI222_X1 U1518 (.ZN(n830), 
	.C2(n5419), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN26_n180), 
	.B1(n5528), 
	.A2(n181), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1519 (.ZN(n3845), 
	.B2(n219), 
	.B1(n181), 
	.A2(n6407), 
	.A1(n5394));
   OAI22_X1 U1520 (.ZN(n3846), 
	.B2(n221), 
	.B1(n181), 
	.A2(n6410), 
	.A1(n5362));
   OAI22_X1 U1521 (.ZN(n3847), 
	.B2(n223), 
	.B1(n181), 
	.A2(n6401), 
	.A1(n5330));
   OAI22_X1 U1522 (.ZN(n3848), 
	.B2(n225), 
	.B1(n181), 
	.A2(n6406), 
	.A1(n5298));
   OAI22_X1 U1523 (.ZN(n3849), 
	.B2(n227), 
	.B1(n181), 
	.A2(n6399), 
	.A1(n5266));
   OAI22_X1 U1524 (.ZN(n3850), 
	.B2(n229), 
	.B1(n181), 
	.A2(n6404), 
	.A1(n5234));
   OAI22_X1 U1525 (.ZN(n3851), 
	.B2(n231), 
	.B1(n181), 
	.A2(n6398), 
	.A1(n5202));
   OAI22_X1 U1526 (.ZN(n3852), 
	.B2(n233), 
	.B1(n181), 
	.A2(n6396), 
	.A1(n5170));
   OAI22_X1 U1527 (.ZN(n3853), 
	.B2(n235), 
	.B1(n181), 
	.A2(n6393), 
	.A1(n5138));
   OAI22_X1 U1528 (.ZN(n3854), 
	.B2(n237), 
	.B1(n181), 
	.A2(n6391), 
	.A1(n5106));
   OAI22_X1 U1529 (.ZN(n3855), 
	.B2(n239), 
	.B1(n181), 
	.A2(n6390), 
	.A1(n5074));
   OAI22_X1 U1530 (.ZN(n3856), 
	.B2(n241), 
	.B1(n181), 
	.A2(n6388), 
	.A1(n5042));
   OAI22_X1 U1531 (.ZN(n3857), 
	.B2(n243), 
	.B1(n181), 
	.A2(n6385), 
	.A1(n5010));
   OAI22_X1 U1532 (.ZN(n3858), 
	.B2(n245), 
	.B1(n181), 
	.A2(n6383), 
	.A1(n4978));
   OAI22_X1 U1533 (.ZN(n3859), 
	.B2(n247), 
	.B1(n181), 
	.A2(n6382), 
	.A1(n4946));
   OAI22_X1 U1534 (.ZN(n3860), 
	.B2(n249), 
	.B1(n181), 
	.A2(n6380), 
	.A1(n4914));
   OAI22_X1 U1535 (.ZN(n3861), 
	.B2(n251), 
	.B1(n181), 
	.A2(n6384), 
	.A1(n4882));
   OAI22_X1 U1536 (.ZN(n3862), 
	.B2(n253), 
	.B1(n181), 
	.A2(n6381), 
	.A1(n4850));
   OAI22_X1 U1537 (.ZN(n3863), 
	.B2(n255), 
	.B1(n181), 
	.A2(n6387), 
	.A1(n4818));
   OAI22_X1 U1538 (.ZN(n3864), 
	.B2(n257), 
	.B1(n181), 
	.A2(n6386), 
	.A1(n4786));
   OAI22_X1 U1539 (.ZN(n3865), 
	.B2(n259), 
	.B1(n181), 
	.A2(n6392), 
	.A1(n4754));
   OAI22_X1 U1540 (.ZN(n3866), 
	.B2(n261), 
	.B1(n181), 
	.A2(n6394), 
	.A1(n4722));
   OAI22_X1 U1541 (.ZN(n3867), 
	.B2(n263), 
	.B1(n181), 
	.A2(n6389), 
	.A1(n4690));
   OAI22_X1 U1542 (.ZN(n3868), 
	.B2(n265), 
	.B1(n181), 
	.A2(n6395), 
	.A1(n4658));
   OAI22_X1 U1543 (.ZN(n3869), 
	.B2(n267), 
	.B1(n181), 
	.A2(n6400), 
	.A1(n4626));
   OAI22_X1 U1544 (.ZN(n3870), 
	.B2(n269), 
	.B1(n181), 
	.A2(n6402), 
	.A1(n4594));
   OAI22_X1 U1545 (.ZN(n3871), 
	.B2(n271), 
	.B1(n181), 
	.A2(n6397), 
	.A1(n4562));
   OAI22_X1 U1546 (.ZN(n3872), 
	.B2(n273), 
	.B1(n181), 
	.A2(n6403), 
	.A1(n4530));
   OAI22_X1 U1547 (.ZN(n3873), 
	.B2(n275), 
	.B1(n181), 
	.A2(n6408), 
	.A1(n4498));
   OAI22_X1 U1548 (.ZN(n3874), 
	.B2(n277), 
	.B1(n181), 
	.A2(n6405), 
	.A1(n4466));
   OAI22_X1 U1549 (.ZN(n3875), 
	.B2(n279), 
	.B1(n181), 
	.A2(n6411), 
	.A1(n4434));
   OAI22_X1 U1552 (.ZN(n3876), 
	.B2(FE_OFN26_n180), 
	.B1(FE_OFN11_net54953), 
	.A2(net54879), 
	.A1(n5473));
   AOI221_X1 U1553 (.ZN(n180), 
	.C2(FE_OFN91_n285), 
	.C1(n5591), 
	.B2(n284), 
	.B1(n832), 
	.A(n833));
   INV_X1 U1554 (.ZN(n833), 
	.A(n834));
   AOI222_X1 U1555 (.ZN(n834), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[26] ), 
	.B2(n5592), 
	.B1(FE_OFN89_n290), 
	.A2(n835), 
	.A1(n288));
   INV_X1 U1556 (.ZN(n835), 
	.A(n5640));
   INV_X1 U1557 (.ZN(n832), 
	.A(n5691));
   OAI22_X1 U1558 (.ZN(n3877), 
	.B2(n172), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N29 ));
   INV_X1 U1559 (.ZN(n172), 
	.A(n836));
   OAI222_X1 U1560 (.ZN(n836), 
	.C2(n5418), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN22_n164), 
	.B1(n5528), 
	.A2(n165), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1561 (.ZN(n3878), 
	.B2(n219), 
	.B1(n165), 
	.A2(n6407), 
	.A1(n5393));
   OAI22_X1 U1562 (.ZN(n3879), 
	.B2(n221), 
	.B1(n165), 
	.A2(n6410), 
	.A1(n5361));
   OAI22_X1 U1563 (.ZN(n3880), 
	.B2(n223), 
	.B1(n165), 
	.A2(n6401), 
	.A1(n5329));
   OAI22_X1 U1564 (.ZN(n3881), 
	.B2(n225), 
	.B1(n165), 
	.A2(n6406), 
	.A1(n5297));
   OAI22_X1 U1565 (.ZN(n3882), 
	.B2(n227), 
	.B1(n165), 
	.A2(n6399), 
	.A1(n5265));
   OAI22_X1 U1566 (.ZN(n3883), 
	.B2(n229), 
	.B1(n165), 
	.A2(n6404), 
	.A1(n5233));
   OAI22_X1 U1567 (.ZN(n3884), 
	.B2(n231), 
	.B1(n165), 
	.A2(n6398), 
	.A1(n5201));
   OAI22_X1 U1568 (.ZN(n3885), 
	.B2(n233), 
	.B1(n165), 
	.A2(n6396), 
	.A1(n5169));
   OAI22_X1 U1569 (.ZN(n3886), 
	.B2(n235), 
	.B1(n165), 
	.A2(n6393), 
	.A1(n5137));
   OAI22_X1 U1570 (.ZN(n3887), 
	.B2(n237), 
	.B1(n165), 
	.A2(n6391), 
	.A1(n5105));
   OAI22_X1 U1571 (.ZN(n3888), 
	.B2(n239), 
	.B1(n165), 
	.A2(n6390), 
	.A1(n5073));
   OAI22_X1 U1572 (.ZN(n3889), 
	.B2(n241), 
	.B1(n165), 
	.A2(n6388), 
	.A1(n5041));
   OAI22_X1 U1573 (.ZN(n3890), 
	.B2(n243), 
	.B1(n165), 
	.A2(n6385), 
	.A1(n5009));
   OAI22_X1 U1574 (.ZN(n3891), 
	.B2(n245), 
	.B1(n165), 
	.A2(n6383), 
	.A1(n4977));
   OAI22_X1 U1575 (.ZN(n3892), 
	.B2(n247), 
	.B1(n165), 
	.A2(n6382), 
	.A1(n4945));
   OAI22_X1 U1576 (.ZN(n3893), 
	.B2(n249), 
	.B1(n165), 
	.A2(n6380), 
	.A1(n4913));
   OAI22_X1 U1577 (.ZN(n3894), 
	.B2(n251), 
	.B1(n165), 
	.A2(n6384), 
	.A1(n4881));
   OAI22_X1 U1578 (.ZN(n3895), 
	.B2(n253), 
	.B1(n165), 
	.A2(n6381), 
	.A1(n4849));
   OAI22_X1 U1579 (.ZN(n3896), 
	.B2(n255), 
	.B1(n165), 
	.A2(n6387), 
	.A1(n4817));
   OAI22_X1 U1580 (.ZN(n3897), 
	.B2(n257), 
	.B1(n165), 
	.A2(n6386), 
	.A1(n4785));
   OAI22_X1 U1581 (.ZN(n3898), 
	.B2(n259), 
	.B1(n165), 
	.A2(n6392), 
	.A1(n4753));
   OAI22_X1 U1582 (.ZN(n3899), 
	.B2(n261), 
	.B1(n165), 
	.A2(n6394), 
	.A1(n4721));
   OAI22_X1 U1583 (.ZN(n3900), 
	.B2(n263), 
	.B1(n165), 
	.A2(n6389), 
	.A1(n4689));
   OAI22_X1 U1584 (.ZN(n3901), 
	.B2(n265), 
	.B1(n165), 
	.A2(n6395), 
	.A1(n4657));
   OAI22_X1 U1585 (.ZN(n3902), 
	.B2(n267), 
	.B1(n165), 
	.A2(n6400), 
	.A1(n4625));
   OAI22_X1 U1586 (.ZN(n3903), 
	.B2(n269), 
	.B1(n165), 
	.A2(n6402), 
	.A1(n4593));
   OAI22_X1 U1587 (.ZN(n3904), 
	.B2(n271), 
	.B1(n165), 
	.A2(n6397), 
	.A1(n4561));
   OAI22_X1 U1588 (.ZN(n3905), 
	.B2(n273), 
	.B1(n165), 
	.A2(n6403), 
	.A1(n4529));
   OAI22_X1 U1589 (.ZN(n3906), 
	.B2(n275), 
	.B1(n165), 
	.A2(n6408), 
	.A1(n4497));
   OAI22_X1 U1590 (.ZN(n3907), 
	.B2(n277), 
	.B1(n165), 
	.A2(n6405), 
	.A1(n4465));
   OAI22_X1 U1591 (.ZN(n3908), 
	.B2(n279), 
	.B1(n165), 
	.A2(n6411), 
	.A1(n4433));
   OAI22_X1 U1594 (.ZN(n3909), 
	.B2(FE_OFN22_n164), 
	.B1(FE_OFN11_net54953), 
	.A2(net54879), 
	.A1(n5470));
   AOI221_X1 U1595 (.ZN(n164), 
	.C2(FE_OFN91_n285), 
	.C1(n5584), 
	.B2(n284), 
	.B1(n838), 
	.A(n839));
   INV_X1 U1596 (.ZN(n839), 
	.A(n840));
   AOI222_X1 U1597 (.ZN(n840), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[27] ), 
	.B2(n5585), 
	.B1(FE_OFN89_n290), 
	.A2(n841), 
	.A1(n288));
   INV_X1 U1598 (.ZN(n841), 
	.A(n5638));
   INV_X1 U1599 (.ZN(n838), 
	.A(n5690));
   OAI22_X1 U1600 (.ZN(n3910), 
	.B2(n160), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N27 ));
   INV_X1 U1601 (.ZN(n160), 
	.A(n842));
   OAI222_X1 U1602 (.ZN(n842), 
	.C2(n5417), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN23_n152), 
	.B1(n5528), 
	.A2(n153), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1603 (.ZN(n3911), 
	.B2(n219), 
	.B1(n153), 
	.A2(n6407), 
	.A1(n5392));
   OAI22_X1 U1604 (.ZN(n3912), 
	.B2(n221), 
	.B1(n153), 
	.A2(n6410), 
	.A1(n5360));
   OAI22_X1 U1605 (.ZN(n3913), 
	.B2(n223), 
	.B1(n153), 
	.A2(n6401), 
	.A1(n5328));
   OAI22_X1 U1606 (.ZN(n3914), 
	.B2(n225), 
	.B1(n153), 
	.A2(n6406), 
	.A1(n5296));
   OAI22_X1 U1607 (.ZN(n3915), 
	.B2(n227), 
	.B1(n153), 
	.A2(n6399), 
	.A1(n5264));
   OAI22_X1 U1608 (.ZN(n3916), 
	.B2(n229), 
	.B1(n153), 
	.A2(n6404), 
	.A1(n5232));
   OAI22_X1 U1609 (.ZN(n3917), 
	.B2(n231), 
	.B1(n153), 
	.A2(n6398), 
	.A1(n5200));
   OAI22_X1 U1610 (.ZN(n3918), 
	.B2(n233), 
	.B1(n153), 
	.A2(n6396), 
	.A1(n5168));
   OAI22_X1 U1611 (.ZN(n3919), 
	.B2(n235), 
	.B1(n153), 
	.A2(n6393), 
	.A1(n5136));
   OAI22_X1 U1612 (.ZN(n3920), 
	.B2(n237), 
	.B1(n153), 
	.A2(n6391), 
	.A1(n5104));
   OAI22_X1 U1613 (.ZN(n3921), 
	.B2(n239), 
	.B1(n153), 
	.A2(n6390), 
	.A1(n5072));
   OAI22_X1 U1614 (.ZN(n3922), 
	.B2(n241), 
	.B1(n153), 
	.A2(n6388), 
	.A1(n5040));
   OAI22_X1 U1615 (.ZN(n3923), 
	.B2(n243), 
	.B1(n153), 
	.A2(n6385), 
	.A1(n5008));
   OAI22_X1 U1616 (.ZN(n3924), 
	.B2(n245), 
	.B1(n153), 
	.A2(n6383), 
	.A1(n4976));
   OAI22_X1 U1617 (.ZN(n3925), 
	.B2(n247), 
	.B1(n153), 
	.A2(n6382), 
	.A1(n4944));
   OAI22_X1 U1618 (.ZN(n3926), 
	.B2(n249), 
	.B1(n153), 
	.A2(n6380), 
	.A1(n4912));
   OAI22_X1 U1619 (.ZN(n3927), 
	.B2(n251), 
	.B1(n153), 
	.A2(n6384), 
	.A1(n4880));
   OAI22_X1 U1620 (.ZN(n3928), 
	.B2(n253), 
	.B1(n153), 
	.A2(n6381), 
	.A1(n4848));
   OAI22_X1 U1621 (.ZN(n3929), 
	.B2(n255), 
	.B1(n153), 
	.A2(n6387), 
	.A1(n4816));
   OAI22_X1 U1622 (.ZN(n3930), 
	.B2(n257), 
	.B1(n153), 
	.A2(n6386), 
	.A1(n4784));
   OAI22_X1 U1623 (.ZN(n3931), 
	.B2(n259), 
	.B1(n153), 
	.A2(n6392), 
	.A1(n4752));
   OAI22_X1 U1624 (.ZN(n3932), 
	.B2(n261), 
	.B1(n153), 
	.A2(n6394), 
	.A1(n4720));
   OAI22_X1 U1625 (.ZN(n3933), 
	.B2(n263), 
	.B1(n153), 
	.A2(n6389), 
	.A1(n4688));
   OAI22_X1 U1626 (.ZN(n3934), 
	.B2(n265), 
	.B1(n153), 
	.A2(n6395), 
	.A1(n4656));
   OAI22_X1 U1627 (.ZN(n3935), 
	.B2(n267), 
	.B1(n153), 
	.A2(n6400), 
	.A1(n4624));
   OAI22_X1 U1628 (.ZN(n3936), 
	.B2(n269), 
	.B1(n153), 
	.A2(n6402), 
	.A1(n4592));
   OAI22_X1 U1629 (.ZN(n3937), 
	.B2(n271), 
	.B1(n153), 
	.A2(n6397), 
	.A1(n4560));
   OAI22_X1 U1630 (.ZN(n3938), 
	.B2(n273), 
	.B1(n153), 
	.A2(n6403), 
	.A1(n4528));
   OAI22_X1 U1631 (.ZN(n3939), 
	.B2(n275), 
	.B1(n153), 
	.A2(n6408), 
	.A1(n4496));
   OAI22_X1 U1632 (.ZN(n3940), 
	.B2(n277), 
	.B1(n153), 
	.A2(n6405), 
	.A1(n4464));
   OAI22_X1 U1633 (.ZN(n3941), 
	.B2(n279), 
	.B1(n153), 
	.A2(n6411), 
	.A1(n4432));
   OAI22_X1 U1636 (.ZN(n3942), 
	.B2(FE_OFN23_n152), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5467));
   AOI221_X1 U1637 (.ZN(n152), 
	.C2(FE_OFN91_n285), 
	.C1(n5577), 
	.B2(n284), 
	.B1(n844), 
	.A(n845));
   INV_X1 U1638 (.ZN(n845), 
	.A(n846));
   AOI222_X1 U1639 (.ZN(n846), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[28] ), 
	.B2(n5578), 
	.B1(FE_OFN89_n290), 
	.A2(n847), 
	.A1(n288));
   INV_X1 U1640 (.ZN(n847), 
	.A(n5636));
   INV_X1 U1641 (.ZN(n844), 
	.A(n5689));
   OAI22_X1 U1642 (.ZN(n3943), 
	.B2(n148), 
	.B1(net54953), 
	.A2(net54881), 
	.A1(\UUT/Mpath/the_alu/N25 ));
   INV_X1 U1643 (.ZN(n148), 
	.A(n848));
   OAI222_X1 U1644 (.ZN(n848), 
	.C2(n5416), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN24_n128), 
	.B1(n5528), 
	.A2(n130), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1645 (.ZN(n3944), 
	.B2(n219), 
	.B1(n130), 
	.A2(n6407), 
	.A1(n5391));
   OAI22_X1 U1646 (.ZN(n3945), 
	.B2(n221), 
	.B1(n130), 
	.A2(n6410), 
	.A1(n5359));
   OAI22_X1 U1647 (.ZN(n3946), 
	.B2(n223), 
	.B1(n130), 
	.A2(n6401), 
	.A1(n5327));
   OAI22_X1 U1648 (.ZN(n3947), 
	.B2(n225), 
	.B1(n130), 
	.A2(n6406), 
	.A1(n5295));
   OAI22_X1 U1649 (.ZN(n3948), 
	.B2(n227), 
	.B1(n130), 
	.A2(n6399), 
	.A1(n5263));
   OAI22_X1 U1650 (.ZN(n3949), 
	.B2(n229), 
	.B1(n130), 
	.A2(n6404), 
	.A1(n5231));
   OAI22_X1 U1651 (.ZN(n3950), 
	.B2(n231), 
	.B1(n130), 
	.A2(n6398), 
	.A1(n5199));
   OAI22_X1 U1652 (.ZN(n3951), 
	.B2(n233), 
	.B1(n130), 
	.A2(n6396), 
	.A1(n5167));
   OAI22_X1 U1653 (.ZN(n3952), 
	.B2(n235), 
	.B1(n130), 
	.A2(n6393), 
	.A1(n5135));
   OAI22_X1 U1654 (.ZN(n3953), 
	.B2(n237), 
	.B1(n130), 
	.A2(n6391), 
	.A1(n5103));
   OAI22_X1 U1655 (.ZN(n3954), 
	.B2(n239), 
	.B1(n130), 
	.A2(n6390), 
	.A1(n5071));
   OAI22_X1 U1656 (.ZN(n3955), 
	.B2(n241), 
	.B1(n130), 
	.A2(n6388), 
	.A1(n5039));
   OAI22_X1 U1657 (.ZN(n3956), 
	.B2(n243), 
	.B1(n130), 
	.A2(n6385), 
	.A1(n5007));
   OAI22_X1 U1658 (.ZN(n3957), 
	.B2(n245), 
	.B1(n130), 
	.A2(n6383), 
	.A1(n4975));
   OAI22_X1 U1659 (.ZN(n3958), 
	.B2(n247), 
	.B1(n130), 
	.A2(n6382), 
	.A1(n4943));
   OAI22_X1 U1660 (.ZN(n3959), 
	.B2(n249), 
	.B1(n130), 
	.A2(n6380), 
	.A1(n4911));
   OAI22_X1 U1661 (.ZN(n3960), 
	.B2(n251), 
	.B1(n130), 
	.A2(n6384), 
	.A1(n4879));
   OAI22_X1 U1662 (.ZN(n3961), 
	.B2(n253), 
	.B1(n130), 
	.A2(n6381), 
	.A1(n4847));
   OAI22_X1 U1663 (.ZN(n3962), 
	.B2(n255), 
	.B1(n130), 
	.A2(n6387), 
	.A1(n4815));
   OAI22_X1 U1664 (.ZN(n3963), 
	.B2(n257), 
	.B1(n130), 
	.A2(n6386), 
	.A1(n4783));
   OAI22_X1 U1665 (.ZN(n3964), 
	.B2(n259), 
	.B1(n130), 
	.A2(n6392), 
	.A1(n4751));
   OAI22_X1 U1666 (.ZN(n3965), 
	.B2(n261), 
	.B1(n130), 
	.A2(n6394), 
	.A1(n4719));
   OAI22_X1 U1667 (.ZN(n3966), 
	.B2(n263), 
	.B1(n130), 
	.A2(n6389), 
	.A1(n4687));
   OAI22_X1 U1668 (.ZN(n3967), 
	.B2(n265), 
	.B1(n130), 
	.A2(n6395), 
	.A1(n4655));
   OAI22_X1 U1669 (.ZN(n3968), 
	.B2(n267), 
	.B1(n130), 
	.A2(n6400), 
	.A1(n4623));
   OAI22_X1 U1670 (.ZN(n3969), 
	.B2(n269), 
	.B1(n130), 
	.A2(n6402), 
	.A1(n4591));
   OAI22_X1 U1671 (.ZN(n3970), 
	.B2(n271), 
	.B1(n130), 
	.A2(n6397), 
	.A1(n4559));
   OAI22_X1 U1672 (.ZN(n3971), 
	.B2(n273), 
	.B1(n130), 
	.A2(n6403), 
	.A1(n4527));
   OAI22_X1 U1673 (.ZN(n3972), 
	.B2(n275), 
	.B1(n130), 
	.A2(n6408), 
	.A1(n4495));
   OAI22_X1 U1674 (.ZN(n3973), 
	.B2(n277), 
	.B1(n130), 
	.A2(n6405), 
	.A1(n4463));
   OAI22_X1 U1675 (.ZN(n3974), 
	.B2(n279), 
	.B1(n130), 
	.A2(n6411), 
	.A1(n4431));
   OAI22_X1 U1678 (.ZN(n3975), 
	.B2(FE_OFN24_n128), 
	.B1(FE_OFN11_net54953), 
	.A2(net54881), 
	.A1(n5464));
   AOI221_X1 U1679 (.ZN(n128), 
	.C2(FE_OFN91_n285), 
	.C1(n5570), 
	.B2(n284), 
	.B1(n850), 
	.A(n851));
   INV_X1 U1680 (.ZN(n851), 
	.A(n852));
   AOI222_X1 U1681 (.ZN(n852), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[29] ), 
	.B2(n5571), 
	.B1(FE_OFN89_n290), 
	.A2(n853), 
	.A1(n288));
   INV_X1 U1682 (.ZN(n853), 
	.A(n5634));
   INV_X1 U1683 (.ZN(n850), 
	.A(n5688));
   OAI222_X1 U1684 (.ZN(n3976), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N24 ), 
	.B2(n119), 
	.B1(net54953), 
	.A2(n123), 
	.A1(n114));
   AOI21_X1 U1685 (.ZN(n119), 
	.B2(n125), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [14]), 
	.A(n126));
   OR2_X1 U1686 (.ZN(n126), 
	.A2(n854), 
	.A1(n176));
   OAI21_X1 U1687 (.ZN(n176), 
	.B2(n855), 
	.B1(n450), 
	.A(n856));
   NOR2_X1 U1688 (.ZN(n125), 
	.A2(n450), 
	.A1(n857));
   INV_X1 U1689 (.ZN(n114), 
	.A(n858));
   OAI222_X1 U1690 (.ZN(n858), 
	.C2(n132), 
	.C1(n5457), 
	.B2(n131), 
	.B1(n860), 
	.A2(n129), 
	.A1(FE_OFN25_n859));
   OAI221_X1 U1693 (.ZN(n3978), 
	.C2(n142), 
	.C1(n5630), 
	.B2(n864), 
	.B1(n140), 
	.A(n865));
   AOI22_X1 U1694 (.ZN(n865), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [30]), 
	.A2(n863), 
	.A1(n144));
   INV_X1 U1695 (.ZN(n863), 
	.A(n5631));
   OAI22_X1 U1696 (.ZN(n3979), 
	.B2(net54873), 
	.B1(n5631), 
	.A2(n866), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U1697 (.ZN(n3980), 
	.B2(FE_OFN8_n73), 
	.B1(n867), 
	.A2(n866), 
	.A1(n147));
   INV_X1 U1698 (.ZN(n866), 
	.A(\UUT/Mpath/the_mult/x_operand1[30] ));
   OAI22_X1 U1699 (.ZN(n3981), 
	.B2(n867), 
	.B1(net54953), 
	.A2(net54883), 
	.A1(\UUT/Mpath/the_alu/N23 ));
   INV_X1 U1700 (.ZN(n867), 
	.A(n868));
   OAI222_X1 U1701 (.ZN(n868), 
	.C2(n5415), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN25_n859), 
	.B1(n5528), 
	.A2(n860), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1702 (.ZN(n3982), 
	.B2(n219), 
	.B1(n860), 
	.A2(n6407), 
	.A1(n5389));
   OAI22_X1 U1703 (.ZN(n3983), 
	.B2(n221), 
	.B1(n860), 
	.A2(n6410), 
	.A1(n5357));
   OAI22_X1 U1704 (.ZN(n3984), 
	.B2(n223), 
	.B1(n860), 
	.A2(n6401), 
	.A1(n5325));
   OAI22_X1 U1705 (.ZN(n3985), 
	.B2(n225), 
	.B1(n860), 
	.A2(n6406), 
	.A1(n5293));
   OAI22_X1 U1706 (.ZN(n3986), 
	.B2(n227), 
	.B1(n860), 
	.A2(n6399), 
	.A1(n5261));
   OAI22_X1 U1707 (.ZN(n3987), 
	.B2(n229), 
	.B1(n860), 
	.A2(n6404), 
	.A1(n5229));
   OAI22_X1 U1708 (.ZN(n3988), 
	.B2(n231), 
	.B1(n860), 
	.A2(n6398), 
	.A1(n5197));
   OAI22_X1 U1709 (.ZN(n3989), 
	.B2(n233), 
	.B1(n860), 
	.A2(n6396), 
	.A1(n5165));
   OAI22_X1 U1710 (.ZN(n3990), 
	.B2(n235), 
	.B1(n860), 
	.A2(n6393), 
	.A1(n5133));
   OAI22_X1 U1711 (.ZN(n3991), 
	.B2(n237), 
	.B1(n860), 
	.A2(n6391), 
	.A1(n5101));
   OAI22_X1 U1712 (.ZN(n3992), 
	.B2(n239), 
	.B1(n860), 
	.A2(n6390), 
	.A1(n5069));
   OAI22_X1 U1713 (.ZN(n3993), 
	.B2(n241), 
	.B1(n860), 
	.A2(n6388), 
	.A1(n5037));
   OAI22_X1 U1714 (.ZN(n3994), 
	.B2(n243), 
	.B1(n860), 
	.A2(n6385), 
	.A1(n5005));
   OAI22_X1 U1715 (.ZN(n3995), 
	.B2(n245), 
	.B1(n860), 
	.A2(n6383), 
	.A1(n4973));
   OAI22_X1 U1716 (.ZN(n3996), 
	.B2(n247), 
	.B1(n860), 
	.A2(n6382), 
	.A1(n4941));
   OAI22_X1 U1717 (.ZN(n3997), 
	.B2(n249), 
	.B1(n860), 
	.A2(n6380), 
	.A1(n4909));
   OAI22_X1 U1718 (.ZN(n3998), 
	.B2(n251), 
	.B1(n860), 
	.A2(n6384), 
	.A1(n4877));
   OAI22_X1 U1719 (.ZN(n3999), 
	.B2(n253), 
	.B1(n860), 
	.A2(n6381), 
	.A1(n4845));
   OAI22_X1 U1720 (.ZN(n4000), 
	.B2(n255), 
	.B1(n860), 
	.A2(n6387), 
	.A1(n4813));
   OAI22_X1 U1721 (.ZN(n4001), 
	.B2(n257), 
	.B1(n860), 
	.A2(n6386), 
	.A1(n4781));
   OAI22_X1 U1722 (.ZN(n4002), 
	.B2(n259), 
	.B1(n860), 
	.A2(n6392), 
	.A1(n4749));
   OAI22_X1 U1723 (.ZN(n4003), 
	.B2(n261), 
	.B1(n860), 
	.A2(n6394), 
	.A1(n4717));
   OAI22_X1 U1724 (.ZN(n4004), 
	.B2(n263), 
	.B1(n860), 
	.A2(n6389), 
	.A1(n4685));
   OAI22_X1 U1725 (.ZN(n4005), 
	.B2(n265), 
	.B1(n860), 
	.A2(n6395), 
	.A1(n4653));
   OAI22_X1 U1726 (.ZN(n4006), 
	.B2(n267), 
	.B1(n860), 
	.A2(n6400), 
	.A1(n4621));
   OAI22_X1 U1727 (.ZN(n4007), 
	.B2(n269), 
	.B1(n860), 
	.A2(n6402), 
	.A1(n4589));
   OAI22_X1 U1728 (.ZN(n4008), 
	.B2(n271), 
	.B1(n860), 
	.A2(n6397), 
	.A1(n4557));
   OAI22_X1 U1729 (.ZN(n4009), 
	.B2(n273), 
	.B1(n860), 
	.A2(n6403), 
	.A1(n4525));
   OAI22_X1 U1730 (.ZN(n4010), 
	.B2(n275), 
	.B1(n860), 
	.A2(n6408), 
	.A1(n4493));
   OAI22_X1 U1731 (.ZN(n4011), 
	.B2(n277), 
	.B1(n860), 
	.A2(n6405), 
	.A1(n4461));
   OAI22_X1 U1732 (.ZN(n4012), 
	.B2(n279), 
	.B1(n860), 
	.A2(n6411), 
	.A1(n4429));
   OAI22_X1 U1735 (.ZN(n4013), 
	.B2(FE_OFN25_n859), 
	.B1(FE_OFN11_net54953), 
	.A2(net54883), 
	.A1(n5458));
   AOI221_X1 U1736 (.ZN(n859), 
	.C2(FE_OFN91_n285), 
	.C1(n5562), 
	.B2(n284), 
	.B1(n870), 
	.A(n871));
   INV_X1 U1737 (.ZN(n871), 
	.A(n872));
   AOI222_X1 U1738 (.ZN(n872), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[30] ), 
	.B2(n5563), 
	.B1(FE_OFN89_n290), 
	.A2(n873), 
	.A1(n288));
   INV_X1 U1739 (.ZN(n873), 
	.A(n5630));
   INV_X1 U1740 (.ZN(n870), 
	.A(n5686));
   OAI222_X1 U1741 (.ZN(n4014), 
	.C2(net54891), 
	.C1(\UUT/Mpath/the_alu/N38 ), 
	.B2(n300), 
	.B1(FE_OFN102_n117), 
	.A2(n123), 
	.A1(n104));
   INV_X1 U1742 (.ZN(n104), 
	.A(n874));
   OAI222_X1 U1743 (.ZN(n874), 
	.C2(n132), 
	.C1(n5481), 
	.B2(n131), 
	.B1(n814), 
	.A2(n129), 
	.A1(n809));
   OAI221_X1 U1745 (.ZN(n812), 
	.C2(n5482), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5760), 
	.A(n282));
   OAI22_X1 U1746 (.ZN(n4015), 
	.B2(n809), 
	.B1(FE_OFN11_net54953), 
	.A2(net54885), 
	.A1(n5482));
   INV_X1 U1747 (.ZN(n809), 
	.A(n875));
   OAI211_X1 U1748 (.ZN(n875), 
	.C2(n321), 
	.C1(n5646), 
	.B(n877), 
	.A(n876));
   AOI222_X1 U1749 (.ZN(n877), 
	.C2(n879), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[23] ), 
	.A2(n878), 
	.A1(FE_OFN91_n285));
   INV_X1 U1750 (.ZN(n879), 
	.A(n5694));
   AOI22_X1 U1751 (.ZN(n876), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[23] ), 
	.A2(n6092), 
	.A1(FE_OFN89_n290));
   INV_X1 U1752 (.ZN(n4016), 
	.A(n880));
   AOI22_X1 U1753 (.ZN(n880), 
	.B2(\UUT/Mpath/out_jar[23] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [23]), 
	.A1(net54847));
   INV_X1 U1754 (.ZN(n4017), 
	.A(n881));
   AOI22_X1 U1755 (.ZN(n881), 
	.B2(\UUT/Mpath/out_jar[22] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [22]), 
	.A1(net54843));
   INV_X1 U1756 (.ZN(n4018), 
	.A(n882));
   AOI22_X1 U1757 (.ZN(n882), 
	.B2(\UUT/Mpath/out_jar[21] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [21]), 
	.A1(net54843));
   INV_X1 U1758 (.ZN(n4019), 
	.A(n883));
   AOI22_X1 U1759 (.ZN(n883), 
	.B2(\UUT/Mpath/out_jar[20] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [20]), 
	.A1(net54843));
   INV_X1 U1760 (.ZN(n4020), 
	.A(n884));
   AOI22_X1 U1761 (.ZN(n884), 
	.B2(\UUT/Mpath/out_jar[19] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [19]), 
	.A1(net54843));
   INV_X1 U1762 (.ZN(n4021), 
	.A(n885));
   AOI22_X1 U1763 (.ZN(n885), 
	.B2(\UUT/Mpath/out_jar[18] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [18]), 
	.A1(net54843));
   INV_X1 U1764 (.ZN(n4022), 
	.A(n886));
   AOI22_X1 U1765 (.ZN(n886), 
	.B2(\UUT/Mpath/out_jar[17] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [17]), 
	.A1(net54843));
   INV_X1 U1766 (.ZN(n4023), 
	.A(n887));
   AOI22_X1 U1767 (.ZN(n887), 
	.B2(\UUT/Mpath/out_jar[16] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [16]), 
	.A1(net54843));
   INV_X1 U1768 (.ZN(n4024), 
	.A(n888));
   AOI22_X1 U1769 (.ZN(n888), 
	.B2(\UUT/Mpath/out_jar[15] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [15]), 
	.A1(net54843));
   INV_X1 U1770 (.ZN(n4025), 
	.A(n889));
   AOI22_X1 U1771 (.ZN(n889), 
	.B2(\UUT/Mpath/out_jar[14] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [14]), 
	.A1(net54843));
   INV_X1 U1772 (.ZN(n4026), 
	.A(n890));
   AOI22_X1 U1773 (.ZN(n890), 
	.B2(\UUT/Mpath/out_jar[13] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [13]), 
	.A1(net54843));
   INV_X1 U1774 (.ZN(n4027), 
	.A(n891));
   AOI22_X1 U1775 (.ZN(n891), 
	.B2(\UUT/Mpath/out_jar[12] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [12]), 
	.A1(net54843));
   INV_X1 U1776 (.ZN(n4028), 
	.A(n892));
   AOI22_X1 U1777 (.ZN(n892), 
	.B2(\UUT/Mpath/out_jar[11] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [11]), 
	.A1(net54845));
   INV_X1 U1778 (.ZN(n4029), 
	.A(n893));
   AOI22_X1 U1779 (.ZN(n893), 
	.B2(\UUT/Mpath/out_jar[10] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [10]), 
	.A1(net54845));
   INV_X1 U1780 (.ZN(n4030), 
	.A(n894));
   AOI22_X1 U1781 (.ZN(n894), 
	.B2(\UUT/Mpath/out_jar[9] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [9]), 
	.A1(net54845));
   INV_X1 U1782 (.ZN(n4031), 
	.A(n895));
   AOI22_X1 U1783 (.ZN(n895), 
	.B2(\UUT/Mpath/out_jar[8] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [8]), 
	.A1(net54845));
   INV_X1 U1784 (.ZN(n4032), 
	.A(n896));
   AOI22_X1 U1785 (.ZN(n896), 
	.B2(\UUT/Mpath/out_jar[7] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [7]), 
	.A1(net54845));
   INV_X1 U1786 (.ZN(n4033), 
	.A(n897));
   AOI22_X1 U1787 (.ZN(n897), 
	.B2(\UUT/Mpath/out_jar[6] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [6]), 
	.A1(net54845));
   INV_X1 U1788 (.ZN(n4034), 
	.A(n898));
   AOI22_X1 U1789 (.ZN(n898), 
	.B2(\UUT/Mpath/out_jar[5] ), 
	.B1(FE_OFN10_net54953), 
	.A2(\UUT/jar_in [5]), 
	.A1(net54845));
   INV_X1 U1790 (.ZN(n4035), 
	.A(n899));
   AOI22_X1 U1791 (.ZN(n899), 
	.B2(\UUT/Mpath/out_jar[4] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [4]), 
	.A1(net54845));
   INV_X1 U1792 (.ZN(n4036), 
	.A(n900));
   AOI22_X1 U1793 (.ZN(n900), 
	.B2(\UUT/Mpath/out_jar[3] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [3]), 
	.A1(net54845));
   INV_X1 U1794 (.ZN(n4037), 
	.A(n901));
   AOI22_X1 U1795 (.ZN(n901), 
	.B2(\UUT/Mpath/out_jar[2] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [2]), 
	.A1(net54845));
   INV_X1 U1796 (.ZN(n4038), 
	.A(n902));
   AOI22_X1 U1797 (.ZN(n902), 
	.B2(\UUT/Mpath/out_jar[1] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [1]), 
	.A1(net54845));
   OAI221_X1 U1798 (.ZN(n4039), 
	.C2(n2725), 
	.C1(n295), 
	.B2(n294), 
	.B1(n68), 
	.A(n903));
   AOI22_X1 U1799 (.ZN(n903), 
	.B2(n6711), 
	.B1(\UUT/jar_in [0]), 
	.A2(n6511), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [0]));
   INV_X1 U1800 (.ZN(n4040), 
	.A(n904));
   AOI22_X1 U1801 (.ZN(n904), 
	.B2(\UUT/Mpath/out_jar[0] ), 
	.B1(net54953), 
	.A2(\UUT/jar_in [0]), 
	.A1(net54845));
   NOR2_X2 U1805 (.ZN(n298), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   NAND2_X1 U1807 (.ZN(n294), 
	.A2(n295), 
	.A1(n908));
   OAI22_X1 U1808 (.ZN(n4042), 
	.B2(n2728), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n6642));
   OAI221_X1 U1809 (.ZN(n4043), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N468 ), 
	.B2(n910), 
	.B1(n5428), 
	.A(n911));
   NAND3_X1 U1810 (.ZN(n911), 
	.A3(n913), 
	.A2(net54869), 
	.A1(n912));
   NAND3_X1 U1811 (.ZN(n912), 
	.A3(n916), 
	.A2(n915), 
	.A1(n914));
   OAI21_X1 U1812 (.ZN(n916), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N2071 ), 
	.A(n917));
   OAI21_X1 U1813 (.ZN(n917), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N2061 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2066 ));
   NAND3_X1 U1814 (.ZN(n914), 
	.A3(n6077), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2060 ), 
	.A1(n918));
   INV_X1 U1815 (.ZN(n918), 
	.A(n919));
   AOI21_X1 U1816 (.ZN(n919), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N2071 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N2047 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   OAI221_X1 U1817 (.ZN(n4044), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N467 ), 
	.B2(n910), 
	.B1(n5427), 
	.A(n920));
   NAND4_X1 U1818 (.ZN(n920), 
	.A4(net54859), 
	.A3(n922), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2054 ), 
	.A1(n921));
   NAND2_X1 U1819 (.ZN(n922), 
	.A2(n924), 
	.A1(n923));
   OAI221_X1 U1820 (.ZN(n4045), 
	.C2(n2729), 
	.C1(net54889), 
	.B2(n910), 
	.B1(n5426), 
	.A(n925));
   OAI221_X1 U1821 (.ZN(n4046), 
	.C2(n2730), 
	.C1(net54891), 
	.B2(n910), 
	.B1(n5425), 
	.A(n925));
   NAND3_X1 U1822 (.ZN(n925), 
	.A3(n927), 
	.A2(n926), 
	.A1(net54875));
   OAI221_X1 U1823 (.ZN(n4047), 
	.C2(net54887), 
	.C1(\UUT/Mpath/the_alu/N453 ), 
	.B2(n910), 
	.B1(n5424), 
	.A(n928));
   NAND4_X1 U1824 (.ZN(n928), 
	.A4(n6030), 
	.A3(net54859), 
	.A2(n930), 
	.A1(n929));
   NAND3_X1 U1825 (.ZN(n930), 
	.A3(n932), 
	.A2(n931), 
	.A1(n6074));
   NAND2_X1 U1826 (.ZN(n910), 
	.A2(n933), 
	.A1(net54877));
   OAI22_X1 U1827 (.ZN(n4048), 
	.B2(n934), 
	.B1(FE_OFN12_net54953), 
	.A2(net54881), 
	.A1(\UUT/Mpath/the_alu/N466 ));
   AOI22_X1 U1828 (.ZN(n934), 
	.B2(n933), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [5]), 
	.A2(n936), 
	.A1(n935));
   NAND2_X1 U1829 (.ZN(n936), 
	.A2(n937), 
	.A1(n923));
   INV_X1 U1830 (.ZN(n923), 
	.A(n926));
   OAI21_X1 U1831 (.ZN(n926), 
	.B2(n6074), 
	.B1(n6076), 
	.A(n931));
   NOR2_X1 U1832 (.ZN(n4049), 
	.A2(n939), 
	.A1(n938));
   AOI22_X1 U1833 (.ZN(n939), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [0]), 
	.B1(net54877), 
	.A2(FE_OFN12_net54953), 
	.A1(\UUT/shift_op [0]));
   NOR2_X1 U1834 (.ZN(n4050), 
	.A2(n940), 
	.A1(n938));
   AOI22_X1 U1835 (.ZN(n940), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [1]), 
	.B1(net54877), 
	.A2(FE_OFN12_net54953), 
	.A1(\UUT/shift_op [1]));
   NOR2_X1 U1836 (.ZN(n4051), 
	.A2(n941), 
	.A1(n938));
   AOI22_X1 U1837 (.ZN(n941), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [2]), 
	.B1(net54877), 
	.A2(FE_OFN12_net54953), 
	.A1(\UUT/shift_op [2]));
   AND2_X1 U1838 (.ZN(n938), 
	.A2(net54895), 
	.A1(n942));
   OAI211_X1 U1839 (.ZN(n942), 
	.C2(n943), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N2037 ), 
	.B(n927), 
	.A(n6028));
   OAI22_X1 U1840 (.ZN(n4052), 
	.B2(n945), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N1877 ), 
	.A2(n944), 
	.A1(net54847));
   INV_X1 U1841 (.ZN(n944), 
	.A(\UUT/exe_outsel [0]));
   OAI22_X1 U1842 (.ZN(n4053), 
	.B2(n945), 
	.B1(n6070), 
	.A2(\UUT/Mpath/N116 ), 
	.A1(net54847));
   OAI221_X1 U1843 (.ZN(n4054), 
	.C2(n142), 
	.C1(n5628), 
	.B2(n946), 
	.B1(n140), 
	.A(n947));
   AOI22_X1 U1844 (.ZN(n947), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [31]), 
	.A2(n948), 
	.A1(n144));
   OAI22_X1 U1845 (.ZN(n4055), 
	.B2(net54871), 
	.B1(n5629), 
	.A2(n949), 
	.A1(FE_OFN10_net54953));
   OAI22_X1 U1846 (.ZN(n4056), 
	.B2(FE_OFN8_n73), 
	.B1(n950), 
	.A2(n949), 
	.A1(n147));
   INV_X1 U1847 (.ZN(n949), 
	.A(FE_OFN177_UUT_Mpath_the_mult_x_operand1_31_));
   OAI22_X1 U1848 (.ZN(n4057), 
	.B2(n950), 
	.B1(net54953), 
	.A2(net54879), 
	.A1(\UUT/Mpath/the_alu/N21 ));
   INV_X1 U1849 (.ZN(n950), 
	.A(n951));
   OAI222_X1 U1850 (.ZN(n951), 
	.C2(n5414), 
	.C1(FE_OFN97_n5529), 
	.B2(FE_OFN13_n953), 
	.B1(n5528), 
	.A2(n952), 
	.A1(FE_OFN96_n5530));
   OAI22_X1 U1851 (.ZN(n4058), 
	.B2(\UUT/Mpath/the_memhandle/N236 ), 
	.B1(net54865), 
	.A2(\UUT/Mpath/the_memhandle/N234 ), 
	.A1(FE_OFN11_net54953));
   OAI22_X1 U1853 (.ZN(n4059), 
	.B2(\UUT/Mpath/the_memhandle/N238 ), 
	.B1(net54865), 
	.A2(\UUT/Mpath/the_memhandle/N237 ), 
	.A1(FE_OFN11_net54953));
   OAI22_X1 U1855 (.ZN(n4060), 
	.B2(net54871), 
	.B1(n5710), 
	.A2(\localbus/c1_op[OP][0] ), 
	.A1(FE_OFN12_net54953));
   OAI21_X1 U1857 (.ZN(n4063), 
	.B2(\UUT/Mpath/the_memhandle/N235 ), 
	.B1(net54847), 
	.A(n957));
   OAI21_X1 U1858 (.ZN(n957), 
	.B2(\UUT/x_we ), 
	.B1(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ), 
	.A(net54859));
   OAI22_X1 U1859 (.ZN(n4064), 
	.B2(n263), 
	.B1(n958), 
	.A2(n6389), 
	.A1(n4678));
   OAI22_X1 U1860 (.ZN(n4065), 
	.B2(n263), 
	.B1(n952), 
	.A2(n6389), 
	.A1(n4684));
   OAI22_X1 U1861 (.ZN(n4066), 
	.B2(n263), 
	.B1(n959), 
	.A2(n6389), 
	.A1(n4707));
   OAI22_X1 U1862 (.ZN(n4067), 
	.B2(n263), 
	.B1(n960), 
	.A2(n262), 
	.A1(n4708));
   NOR3_X1 U1864 (.ZN(n262), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N439 ));
   OAI22_X1 U1865 (.ZN(n4068), 
	.B2(n257), 
	.B1(n958), 
	.A2(n6386), 
	.A1(n4774));
   OAI22_X1 U1866 (.ZN(n4069), 
	.B2(n257), 
	.B1(n952), 
	.A2(n6386), 
	.A1(n4780));
   OAI22_X1 U1867 (.ZN(n4070), 
	.B2(n257), 
	.B1(n959), 
	.A2(n6386), 
	.A1(n4803));
   OAI22_X1 U1868 (.ZN(n4071), 
	.B2(n257), 
	.B1(n960), 
	.A2(n256), 
	.A1(n4804));
   NOR3_X1 U1870 (.ZN(n256), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N439 ));
   OAI22_X1 U1871 (.ZN(n4072), 
	.B2(n253), 
	.B1(n958), 
	.A2(n6381), 
	.A1(n4838));
   OAI22_X1 U1872 (.ZN(n4073), 
	.B2(n253), 
	.B1(n952), 
	.A2(n6381), 
	.A1(n4844));
   OAI22_X1 U1873 (.ZN(n4074), 
	.B2(n253), 
	.B1(n959), 
	.A2(n6381), 
	.A1(n4867));
   OAI22_X1 U1874 (.ZN(n4075), 
	.B2(n253), 
	.B1(n960), 
	.A2(n252), 
	.A1(n4868));
   NOR3_X1 U1876 (.ZN(n252), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N415 ));
   OAI22_X1 U1877 (.ZN(n4076), 
	.B2(n249), 
	.B1(n958), 
	.A2(n6380), 
	.A1(n4902));
   OAI22_X1 U1878 (.ZN(n4077), 
	.B2(n249), 
	.B1(n952), 
	.A2(n6380), 
	.A1(n4908));
   OAI22_X1 U1879 (.ZN(n4078), 
	.B2(n249), 
	.B1(n959), 
	.A2(n6380), 
	.A1(n4931));
   OAI22_X1 U1880 (.ZN(n4079), 
	.B2(n249), 
	.B1(n960), 
	.A2(n248), 
	.A1(n4932));
   NOR3_X1 U1882 (.ZN(n248), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N415 ));
   OAI22_X1 U1883 (.ZN(n4080), 
	.B2(n245), 
	.B1(n958), 
	.A2(n6383), 
	.A1(n4966));
   OAI22_X1 U1884 (.ZN(n4081), 
	.B2(n245), 
	.B1(n952), 
	.A2(n6383), 
	.A1(n4972));
   OAI22_X1 U1885 (.ZN(n4082), 
	.B2(n245), 
	.B1(n959), 
	.A2(n6383), 
	.A1(n4995));
   OAI22_X1 U1886 (.ZN(n4083), 
	.B2(n245), 
	.B1(n960), 
	.A2(n244), 
	.A1(n4996));
   NOR3_X1 U1888 (.ZN(n244), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N391 ));
   OAI22_X1 U1889 (.ZN(n4084), 
	.B2(n241), 
	.B1(n958), 
	.A2(n6388), 
	.A1(n5030));
   OAI22_X1 U1890 (.ZN(n4085), 
	.B2(n241), 
	.B1(n952), 
	.A2(n6388), 
	.A1(n5036));
   OAI22_X1 U1891 (.ZN(n4086), 
	.B2(n241), 
	.B1(n959), 
	.A2(n6388), 
	.A1(n5059));
   OAI22_X1 U1892 (.ZN(n4087), 
	.B2(n241), 
	.B1(n960), 
	.A2(n240), 
	.A1(n5060));
   NOR3_X1 U1894 (.ZN(n240), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N391 ));
   OAI22_X1 U1895 (.ZN(n4088), 
	.B2(n235), 
	.B1(n958), 
	.A2(n6393), 
	.A1(n5126));
   OAI22_X1 U1896 (.ZN(n4089), 
	.B2(n235), 
	.B1(n952), 
	.A2(n6393), 
	.A1(n5132));
   OAI22_X1 U1897 (.ZN(n4090), 
	.B2(n235), 
	.B1(n959), 
	.A2(n6393), 
	.A1(n5155));
   OAI22_X1 U1898 (.ZN(n4091), 
	.B2(n235), 
	.B1(n960), 
	.A2(n234), 
	.A1(n5156));
   NOR3_X1 U1900 (.ZN(n234), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N367 ));
   OAI22_X1 U1901 (.ZN(n4092), 
	.B2(n231), 
	.B1(n958), 
	.A2(n6398), 
	.A1(n5190));
   OAI22_X1 U1902 (.ZN(n4093), 
	.B2(n231), 
	.B1(n952), 
	.A2(n6398), 
	.A1(n5196));
   OAI22_X1 U1903 (.ZN(n4094), 
	.B2(n231), 
	.B1(n959), 
	.A2(n6398), 
	.A1(n5219));
   OAI22_X1 U1904 (.ZN(n4095), 
	.B2(n231), 
	.B1(n960), 
	.A2(n230), 
	.A1(n5220));
   NOR3_X1 U1906 (.ZN(n230), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N367 ));
   OAI22_X1 U1907 (.ZN(n4096), 
	.B2(n227), 
	.B1(n958), 
	.A2(n6399), 
	.A1(n5254));
   OAI22_X1 U1908 (.ZN(n4097), 
	.B2(n227), 
	.B1(n952), 
	.A2(n6399), 
	.A1(n5260));
   OAI22_X1 U1909 (.ZN(n4098), 
	.B2(n227), 
	.B1(n959), 
	.A2(n6399), 
	.A1(n5283));
   OAI22_X1 U1910 (.ZN(n4099), 
	.B2(n227), 
	.B1(n960), 
	.A2(n226), 
	.A1(n5284));
   NOR3_X1 U1912 (.ZN(n226), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N342 ));
   OAI22_X1 U1913 (.ZN(n4100), 
	.B2(n223), 
	.B1(n958), 
	.A2(n6401), 
	.A1(n5318));
   OAI22_X1 U1914 (.ZN(n4101), 
	.B2(n223), 
	.B1(n952), 
	.A2(n6401), 
	.A1(n5324));
   OAI22_X1 U1915 (.ZN(n4102), 
	.B2(n223), 
	.B1(n959), 
	.A2(n6401), 
	.A1(n5347));
   OAI22_X1 U1916 (.ZN(n4103), 
	.B2(n223), 
	.B1(n960), 
	.A2(n222), 
	.A1(n5348));
   NOR3_X1 U1918 (.ZN(n222), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N342 ));
   OAI22_X1 U1919 (.ZN(n4104), 
	.B2(n219), 
	.B1(n958), 
	.A2(n6407), 
	.A1(n5382));
   OAI22_X1 U1920 (.ZN(n4105), 
	.B2(n219), 
	.B1(n952), 
	.A2(n6407), 
	.A1(n5388));
   OAI22_X1 U1921 (.ZN(n4106), 
	.B2(n219), 
	.B1(n959), 
	.A2(n6407), 
	.A1(n5411));
   OAI22_X1 U1922 (.ZN(n4107), 
	.B2(n219), 
	.B1(n960), 
	.A2(n218), 
	.A1(n5412));
   NOR3_X1 U1924 (.ZN(n218), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N318 ));
   OAI22_X1 U1925 (.ZN(n4108), 
	.B2(n277), 
	.B1(n958), 
	.A2(n6405), 
	.A1(n4454));
   OAI22_X1 U1926 (.ZN(n4109), 
	.B2(n277), 
	.B1(n952), 
	.A2(n6405), 
	.A1(n4460));
   OAI22_X1 U1927 (.ZN(n4110), 
	.B2(n277), 
	.B1(n959), 
	.A2(n6405), 
	.A1(n4483));
   OAI22_X1 U1928 (.ZN(n4111), 
	.B2(n277), 
	.B1(n960), 
	.A2(n276), 
	.A1(n4484));
   NOR3_X1 U1930 (.ZN(n276), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N318 ));
   OAI22_X1 U1931 (.ZN(n4112), 
	.B2(n273), 
	.B1(n958), 
	.A2(n6403), 
	.A1(n4518));
   OAI22_X1 U1932 (.ZN(n4113), 
	.B2(n273), 
	.B1(n952), 
	.A2(n6403), 
	.A1(n4524));
   OAI22_X1 U1933 (.ZN(n4114), 
	.B2(n273), 
	.B1(n959), 
	.A2(n6403), 
	.A1(n4547));
   OAI22_X1 U1934 (.ZN(n4115), 
	.B2(n273), 
	.B1(n960), 
	.A2(n272), 
	.A1(n4548));
   NOR3_X1 U1936 (.ZN(n272), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N293 ));
   OAI22_X1 U1937 (.ZN(n4116), 
	.B2(n269), 
	.B1(n958), 
	.A2(n6402), 
	.A1(n4582));
   OAI22_X1 U1938 (.ZN(n4117), 
	.B2(n269), 
	.B1(n952), 
	.A2(n6402), 
	.A1(n4588));
   OAI22_X1 U1939 (.ZN(n4118), 
	.B2(n269), 
	.B1(n959), 
	.A2(n6402), 
	.A1(n4611));
   OAI22_X1 U1940 (.ZN(n4119), 
	.B2(n269), 
	.B1(n960), 
	.A2(n268), 
	.A1(n4612));
   NOR3_X1 U1942 (.ZN(n268), 
	.A3(n962), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N293 ));
   NAND2_X1 U1943 (.ZN(n962), 
	.A2(n964), 
	.A1(n963));
   OAI22_X1 U1944 (.ZN(n4120), 
	.B2(n261), 
	.B1(n958), 
	.A2(n6394), 
	.A1(n4710));
   OAI22_X1 U1945 (.ZN(n4121), 
	.B2(n261), 
	.B1(n952), 
	.A2(n6394), 
	.A1(n4716));
   OAI22_X1 U1946 (.ZN(n4122), 
	.B2(n261), 
	.B1(n959), 
	.A2(n6394), 
	.A1(n4739));
   OAI22_X1 U1947 (.ZN(n4123), 
	.B2(n261), 
	.B1(n960), 
	.A2(n260), 
	.A1(n4740));
   NOR3_X1 U1949 (.ZN(n260), 
	.A3(n961), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N273 ));
   NAND2_X1 U1950 (.ZN(n961), 
	.A2(n964), 
	.A1(\UUT/rd_addr [1]));
   OAI22_X1 U1951 (.ZN(n4124), 
	.B2(n265), 
	.B1(n958), 
	.A2(n6395), 
	.A1(n4646));
   OAI22_X1 U1952 (.ZN(n4125), 
	.B2(n265), 
	.B1(n952), 
	.A2(n6395), 
	.A1(n4652));
   OAI22_X1 U1953 (.ZN(n4126), 
	.B2(n265), 
	.B1(n959), 
	.A2(n6395), 
	.A1(n4675));
   OAI22_X1 U1954 (.ZN(n4127), 
	.B2(n265), 
	.B1(n960), 
	.A2(n264), 
	.A1(n4676));
   NOR3_X1 U1956 (.ZN(n264), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N439 ));
   OAI22_X1 U1957 (.ZN(n4128), 
	.B2(n259), 
	.B1(n958), 
	.A2(n6392), 
	.A1(n4742));
   OAI22_X1 U1958 (.ZN(n4129), 
	.B2(n259), 
	.B1(n952), 
	.A2(n6392), 
	.A1(n4748));
   OAI22_X1 U1959 (.ZN(n4130), 
	.B2(n259), 
	.B1(n959), 
	.A2(n6392), 
	.A1(n4771));
   OAI22_X1 U1960 (.ZN(n4131), 
	.B2(n259), 
	.B1(n960), 
	.A2(n258), 
	.A1(n4772));
   NOR3_X1 U1962 (.ZN(n258), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N439 ));
   OAI22_X1 U1963 (.ZN(n4132), 
	.B2(n255), 
	.B1(n958), 
	.A2(n6387), 
	.A1(n4806));
   OAI22_X1 U1964 (.ZN(n4133), 
	.B2(n255), 
	.B1(n952), 
	.A2(n6387), 
	.A1(n4812));
   OAI22_X1 U1965 (.ZN(n4134), 
	.B2(n255), 
	.B1(n959), 
	.A2(n6387), 
	.A1(n4835));
   OAI22_X1 U1966 (.ZN(n4135), 
	.B2(n255), 
	.B1(n960), 
	.A2(n254), 
	.A1(n4836));
   NOR3_X1 U1968 (.ZN(n254), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N415 ));
   OAI22_X1 U1969 (.ZN(n4136), 
	.B2(n251), 
	.B1(n958), 
	.A2(n6384), 
	.A1(n4870));
   OAI22_X1 U1970 (.ZN(n4137), 
	.B2(n251), 
	.B1(n952), 
	.A2(n6384), 
	.A1(n4876));
   OAI22_X1 U1971 (.ZN(n4138), 
	.B2(n251), 
	.B1(n959), 
	.A2(n6384), 
	.A1(n4899));
   OAI22_X1 U1972 (.ZN(n4139), 
	.B2(n251), 
	.B1(n960), 
	.A2(n250), 
	.A1(n4900));
   NOR3_X1 U1974 (.ZN(n250), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N415 ));
   OAI22_X1 U1975 (.ZN(n4140), 
	.B2(n247), 
	.B1(n958), 
	.A2(n6382), 
	.A1(n4934));
   OAI22_X1 U1976 (.ZN(n4141), 
	.B2(n247), 
	.B1(n952), 
	.A2(n6382), 
	.A1(n4940));
   OAI22_X1 U1977 (.ZN(n4142), 
	.B2(n247), 
	.B1(n959), 
	.A2(n6382), 
	.A1(n4963));
   OAI22_X1 U1978 (.ZN(n4143), 
	.B2(n247), 
	.B1(n960), 
	.A2(n246), 
	.A1(n4964));
   NOR3_X1 U1980 (.ZN(n246), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N391 ));
   OAI22_X1 U1981 (.ZN(n4144), 
	.B2(n243), 
	.B1(n958), 
	.A2(n6385), 
	.A1(n4998));
   OAI22_X1 U1982 (.ZN(n4145), 
	.B2(n243), 
	.B1(n952), 
	.A2(n6385), 
	.A1(n5004));
   OAI22_X1 U1983 (.ZN(n4146), 
	.B2(n243), 
	.B1(n959), 
	.A2(n6385), 
	.A1(n5027));
   OAI22_X1 U1984 (.ZN(n4147), 
	.B2(n243), 
	.B1(n960), 
	.A2(n242), 
	.A1(n5028));
   NOR3_X1 U1986 (.ZN(n242), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N391 ));
   OAI22_X1 U1987 (.ZN(n4148), 
	.B2(n237), 
	.B1(n958), 
	.A2(n6391), 
	.A1(n5094));
   OAI22_X1 U1988 (.ZN(n4149), 
	.B2(n237), 
	.B1(n952), 
	.A2(n6391), 
	.A1(n5100));
   OAI22_X1 U1989 (.ZN(n4150), 
	.B2(n237), 
	.B1(n959), 
	.A2(n6391), 
	.A1(n5123));
   OAI22_X1 U1990 (.ZN(n4151), 
	.B2(n237), 
	.B1(n960), 
	.A2(n236), 
	.A1(n5124));
   NOR3_X1 U1992 (.ZN(n236), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N367 ));
   OAI22_X1 U1993 (.ZN(n4152), 
	.B2(n233), 
	.B1(n958), 
	.A2(n6396), 
	.A1(n5158));
   OAI22_X1 U1994 (.ZN(n4153), 
	.B2(n233), 
	.B1(n952), 
	.A2(n6396), 
	.A1(n5164));
   OAI22_X1 U1995 (.ZN(n4154), 
	.B2(n233), 
	.B1(n959), 
	.A2(n6396), 
	.A1(n5187));
   OAI22_X1 U1996 (.ZN(n4155), 
	.B2(n233), 
	.B1(n960), 
	.A2(n232), 
	.A1(n5188));
   NOR3_X1 U1998 (.ZN(n232), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N367 ));
   OAI22_X1 U1999 (.ZN(n4156), 
	.B2(n229), 
	.B1(n958), 
	.A2(n6404), 
	.A1(n5222));
   OAI22_X1 U2000 (.ZN(n4157), 
	.B2(n229), 
	.B1(n952), 
	.A2(n6404), 
	.A1(n5228));
   OAI22_X1 U2001 (.ZN(n4158), 
	.B2(n229), 
	.B1(n959), 
	.A2(n6404), 
	.A1(n5251));
   OAI22_X1 U2002 (.ZN(n4159), 
	.B2(n229), 
	.B1(n960), 
	.A2(n228), 
	.A1(n5252));
   NOR3_X1 U2004 (.ZN(n228), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N342 ));
   OAI22_X1 U2005 (.ZN(n4160), 
	.B2(n225), 
	.B1(n958), 
	.A2(n6406), 
	.A1(n5286));
   OAI22_X1 U2006 (.ZN(n4161), 
	.B2(n225), 
	.B1(n952), 
	.A2(n6406), 
	.A1(n5292));
   OAI22_X1 U2007 (.ZN(n4162), 
	.B2(n225), 
	.B1(n959), 
	.A2(n6406), 
	.A1(n5315));
   OAI22_X1 U2008 (.ZN(n4163), 
	.B2(n225), 
	.B1(n960), 
	.A2(n224), 
	.A1(n5316));
   NOR3_X1 U2010 (.ZN(n224), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N342 ));
   OAI22_X1 U2011 (.ZN(n4164), 
	.B2(n221), 
	.B1(n958), 
	.A2(n6410), 
	.A1(n5350));
   OAI22_X1 U2012 (.ZN(n4165), 
	.B2(n221), 
	.B1(n952), 
	.A2(n6410), 
	.A1(n5356));
   OAI22_X1 U2013 (.ZN(n4166), 
	.B2(n221), 
	.B1(n959), 
	.A2(n6410), 
	.A1(n5379));
   OAI22_X1 U2014 (.ZN(n4167), 
	.B2(n221), 
	.B1(n960), 
	.A2(n220), 
	.A1(n5380));
   NOR3_X1 U2016 (.ZN(n220), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N318 ));
   OAI22_X1 U2017 (.ZN(n4168), 
	.B2(n279), 
	.B1(n958), 
	.A2(n6411), 
	.A1(n4422));
   OAI22_X1 U2018 (.ZN(n4169), 
	.B2(n279), 
	.B1(n952), 
	.A2(n6411), 
	.A1(n4428));
   OAI22_X1 U2019 (.ZN(n4170), 
	.B2(n279), 
	.B1(n959), 
	.A2(n6411), 
	.A1(n4451));
   OAI22_X1 U2020 (.ZN(n4171), 
	.B2(n279), 
	.B1(n960), 
	.A2(n278), 
	.A1(n4452));
   NOR3_X1 U2022 (.ZN(n278), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N318 ));
   OAI22_X1 U2023 (.ZN(n4172), 
	.B2(n275), 
	.B1(n958), 
	.A2(n6408), 
	.A1(n4486));
   OAI22_X1 U2024 (.ZN(n4173), 
	.B2(n275), 
	.B1(n952), 
	.A2(n6408), 
	.A1(n4492));
   OAI22_X1 U2025 (.ZN(n4174), 
	.B2(n275), 
	.B1(n959), 
	.A2(n6408), 
	.A1(n4515));
   OAI22_X1 U2026 (.ZN(n4175), 
	.B2(n275), 
	.B1(n960), 
	.A2(n274), 
	.A1(n4516));
   NOR3_X1 U2028 (.ZN(n274), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N293 ));
   OAI22_X1 U2029 (.ZN(n4176), 
	.B2(n271), 
	.B1(n958), 
	.A2(n6397), 
	.A1(n4550));
   OAI22_X1 U2030 (.ZN(n4177), 
	.B2(n271), 
	.B1(n952), 
	.A2(n6397), 
	.A1(n4556));
   OAI22_X1 U2031 (.ZN(n4178), 
	.B2(n271), 
	.B1(n959), 
	.A2(n6397), 
	.A1(n4579));
   OAI22_X1 U2032 (.ZN(n4179), 
	.B2(n271), 
	.B1(n960), 
	.A2(n270), 
	.A1(n4580));
   NOR3_X1 U2034 (.ZN(n270), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N293 ));
   OAI22_X1 U2035 (.ZN(n4180), 
	.B2(n267), 
	.B1(n958), 
	.A2(n6400), 
	.A1(n4614));
   OAI22_X1 U2036 (.ZN(n4181), 
	.B2(n267), 
	.B1(n952), 
	.A2(n6400), 
	.A1(n4620));
   OAI22_X1 U2037 (.ZN(n4182), 
	.B2(n267), 
	.B1(n959), 
	.A2(n6400), 
	.A1(n4643));
   OAI22_X1 U2038 (.ZN(n4183), 
	.B2(n267), 
	.B1(n960), 
	.A2(n266), 
	.A1(n4644));
   NOR3_X1 U2040 (.ZN(n266), 
	.A3(n965), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N273 ));
   NAND2_X1 U2041 (.ZN(n965), 
	.A2(\UUT/rd_addr [1]), 
	.A1(n967));
   OAI22_X1 U2042 (.ZN(n4184), 
	.B2(n239), 
	.B1(n958), 
	.A2(n6390), 
	.A1(n5062));
   OAI22_X1 U2043 (.ZN(n4185), 
	.B2(n239), 
	.B1(n952), 
	.A2(n6390), 
	.A1(n5068));
   OAI22_X1 U2044 (.ZN(n4186), 
	.B2(n239), 
	.B1(n959), 
	.A2(n6390), 
	.A1(n5091));
   OAI22_X1 U2045 (.ZN(n4187), 
	.B2(n239), 
	.B1(n960), 
	.A2(n238), 
	.A1(n5092));
   NOR3_X1 U2047 (.ZN(n238), 
	.A3(n966), 
	.A2(FE_OFN11_net54953), 
	.A1(\UUT/regfile/N273 ));
   NAND2_X1 U2048 (.ZN(n966), 
	.A2(n963), 
	.A1(n967));
   INV_X1 U2049 (.ZN(n963), 
	.A(\UUT/rd_addr [1]));
   INV_X1 U2050 (.ZN(n967), 
	.A(n964));
   NAND2_X1 U2051 (.ZN(n964), 
	.A2(n5413), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[0] ));
   OAI221_X1 U2052 (.ZN(n4188), 
	.C2(n142), 
	.C1(n5676), 
	.B2(n968), 
	.B1(n140), 
	.A(n969));
   AOI22_X1 U2053 (.ZN(n969), 
	.B2(n145), 
	.B1(\UUT/Mpath/the_mult/Mad_out [0]), 
	.A2(n970), 
	.A1(n144));
   NOR2_X1 U2055 (.ZN(n972), 
	.A2(n974), 
	.A1(n973));
   INV_X1 U2057 (.ZN(n973), 
	.A(\UUT/Mpath/the_mult/N255 ));
   NAND3_X1 U2059 (.ZN(n976), 
	.A3(\UUT/Mpath/the_mult/N255 ), 
	.A2(n974), 
	.A1(n971));
   INV_X1 U2060 (.ZN(n974), 
	.A(\UUT/Mpath/the_mult/N312 ));
   INV_X1 U2061 (.ZN(n971), 
	.A(\UUT/Mpath/the_mult/N311 ));
   OAI22_X1 U2063 (.ZN(n4189), 
	.B2(net54871), 
	.B1(n5413), 
	.A2(\UUT/Mcontrol/bp_logicA/N9 ), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2064 (.ZN(n4190), 
	.B2(\UUT/Mcontrol/bp_logicA/N9 ), 
	.B1(net54863), 
	.A2(n978), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2065 (.ZN(n4191), 
	.B2(n2732), 
	.B1(n295), 
	.A2(FE_OFCN206_FE_OFN186_n546), 
	.A1(n979));
   OAI22_X1 U2066 (.ZN(n4192), 
	.B2(n981), 
	.B1(net54863), 
	.A2(n980), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2067 (.ZN(n981), 
	.A(\UUT/Mcontrol/m_sampled_xrd[0] ));
   OAI221_X1 U2068 (.ZN(n4193), 
	.C2(n980), 
	.C1(net54889), 
	.B2(n982), 
	.B1(n6037), 
	.A(n983));
   AOI221_X1 U2069 (.ZN(n983), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [16]), 
	.C1(n985), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [11]), 
	.B1(n984), 
	.A(FE_OFN9_n986));
   INV_X1 U2070 (.ZN(n980), 
	.A(\UUT/Mcontrol/x_rd[0] ));
   OAI22_X1 U2071 (.ZN(n4194), 
	.B2(n2735), 
	.B1(net54863), 
	.A2(n987), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U2072 (.ZN(n4195), 
	.C2(n987), 
	.C1(net54891), 
	.B2(n982), 
	.B1(n5896), 
	.A(n988));
   AOI221_X1 U2073 (.ZN(n988), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [17]), 
	.C1(n985), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [12]), 
	.B1(n984), 
	.A(FE_OFN9_n986));
   INV_X1 U2074 (.ZN(n987), 
	.A(\UUT/Mcontrol/x_rd[1] ));
   OAI22_X1 U2075 (.ZN(n4196), 
	.B2(n2737), 
	.B1(net54863), 
	.A2(n989), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U2076 (.ZN(n4197), 
	.C2(n989), 
	.C1(net54889), 
	.B2(n982), 
	.B1(n5888), 
	.A(n990));
   AOI221_X1 U2077 (.ZN(n990), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [18]), 
	.C1(n985), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [13]), 
	.B1(n984), 
	.A(FE_OFN9_n986));
   INV_X1 U2078 (.ZN(n989), 
	.A(\UUT/Mcontrol/x_rd[2] ));
   OAI22_X1 U2079 (.ZN(n4198), 
	.B2(n2739), 
	.B1(net54863), 
	.A2(n991), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U2080 (.ZN(n4199), 
	.C2(n991), 
	.C1(net54889), 
	.B2(n982), 
	.B1(n5879), 
	.A(n992));
   AOI221_X1 U2081 (.ZN(n992), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [19]), 
	.C1(n985), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [14]), 
	.B1(n984), 
	.A(FE_OFN9_n986));
   INV_X1 U2082 (.ZN(n991), 
	.A(\UUT/Mcontrol/x_rd[3] ));
   OAI22_X1 U2083 (.ZN(n4200), 
	.B2(n2741), 
	.B1(net54861), 
	.A2(n993), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U2084 (.ZN(n4201), 
	.C2(n993), 
	.C1(net54889), 
	.B2(n982), 
	.B1(n5871), 
	.A(n994));
   AOI221_X1 U2085 (.ZN(n994), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [20]), 
	.C1(n985), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [15]), 
	.B1(n984), 
	.A(FE_OFN9_n986));
   NOR4_X1 U2086 (.ZN(n986), 
	.A4(\UUT/Mcontrol/Operation_decoding32/N1970 ), 
	.A3(n6038), 
	.A2(n6039), 
	.A1(n995));
   AND2_X1 U2087 (.ZN(n985), 
	.A2(net54895), 
	.A1(n996));
   OAI21_X1 U2088 (.ZN(n996), 
	.B2(n998), 
	.B1(n997), 
	.A(n999));
   INV_X1 U2089 (.ZN(n999), 
	.A(n1000));
   AOI21_X1 U2090 (.ZN(n1000), 
	.B2(n6075), 
	.B1(n929), 
	.A(n933));
   AOI221_X1 U2091 (.ZN(n997), 
	.C2(n1003), 
	.C1(n1002), 
	.B2(n931), 
	.B1(n1001), 
	.A(n1004));
   NAND3_X1 U2092 (.ZN(n1003), 
	.A3(n6043), 
	.A2(n6042), 
	.A1(n6041));
   NAND2_X1 U2093 (.ZN(n1001), 
	.A2(n857), 
	.A1(n6051));
   AOI21_X1 U2094 (.ZN(n984), 
	.B2(n6030), 
	.B1(n1005), 
	.A(FE_OFN12_net54953));
   OR3_X1 U2095 (.ZN(n1005), 
	.A3(n1004), 
	.A2(n931), 
	.A1(n998));
   INV_X1 U2096 (.ZN(n993), 
	.A(\UUT/Mcontrol/x_rd[4] ));
   NAND3_X1 U2097 (.ZN(n982), 
	.A3(n1007), 
	.A2(n1006), 
	.A1(n6044));
   NOR3_X1 U2098 (.ZN(n1007), 
	.A3(n6067), 
	.A2(n6079), 
	.A1(n1008));
   INV_X1 U2099 (.ZN(n1006), 
	.A(n995));
   NAND3_X1 U2100 (.ZN(n995), 
	.A3(n1002), 
	.A2(net54869), 
	.A1(n921));
   NOR3_X1 U2101 (.ZN(n1002), 
	.A3(n1004), 
	.A2(n6048), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2019 ));
   INV_X1 U2102 (.ZN(n921), 
	.A(n998));
   NAND3_X1 U2103 (.ZN(n998), 
	.A3(n6075), 
	.A2(n6030), 
	.A1(n929));
   OAI22_X1 U2104 (.ZN(n4202), 
	.B2(\UUT/Mpath/the_mult/N231 ), 
	.B1(net54861), 
	.A2(n1009), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2105 (.ZN(n4203), 
	.B2(n1009), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N223 ), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2106 (.ZN(n1009), 
	.A(\UUT/Mpath/the_mult/x_mul_command[0] ));
   OAI22_X1 U2107 (.ZN(n4204), 
	.B2(n295), 
	.B1(n5428), 
	.A2(n1011), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2108 (.ZN(n1011), 
	.A(I_DATA_INBUS[0]));
   OAI22_X1 U2109 (.ZN(n4205), 
	.B2(\UUT/Mpath/the_mult/N230 ), 
	.B1(net54861), 
	.A2(n1012), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2110 (.ZN(n4206), 
	.B2(n1012), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N222 ), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2111 (.ZN(n1012), 
	.A(\UUT/Mpath/the_mult/x_mul_command[1] ));
   OAI22_X1 U2112 (.ZN(n4207), 
	.B2(\UUT/Mcontrol/st_logic/N27 ), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N222 ), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2114 (.ZN(n4208), 
	.B2(n295), 
	.B1(n5427), 
	.A2(n1014), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2115 (.ZN(n1014), 
	.A(I_DATA_INBUS[1]));
   OAI22_X1 U2116 (.ZN(n4209), 
	.B2(\UUT/Mpath/the_mult/N244 ), 
	.B1(net54861), 
	.A2(n1015), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2117 (.ZN(n4210), 
	.B2(n1015), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N221 ), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2118 (.ZN(n1015), 
	.A(\UUT/Mpath/the_mult/x_mul_command[2] ));
   OAI22_X1 U2119 (.ZN(n4211), 
	.B2(\UUT/Mcontrol/st_logic/N26 ), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N221 ), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2121 (.ZN(n4212), 
	.B2(n295), 
	.B1(n5426), 
	.A2(n1017), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2122 (.ZN(n1017), 
	.A(I_DATA_INBUS[2]));
   OAI22_X1 U2123 (.ZN(n4213), 
	.B2(\UUT/Mpath/the_mult/N229 ), 
	.B1(net54861), 
	.A2(n1018), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2124 (.ZN(n4214), 
	.B2(n1018), 
	.B1(net54861), 
	.A2(\UUT/Mpath/the_mult/N220 ), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2125 (.ZN(n1018), 
	.A(\UUT/Mpath/the_mult/x_mul_command[3] ));
   OAI22_X1 U2126 (.ZN(n4215), 
	.B2(n2748), 
	.B1(net54859), 
	.A2(\UUT/Mpath/the_mult/N220 ), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2128 (.ZN(n4216), 
	.B2(n295), 
	.B1(n5425), 
	.A2(n1020), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2129 (.ZN(n1020), 
	.A(I_DATA_INBUS[3]));
   OAI22_X1 U2130 (.ZN(n4217), 
	.B2(n2750), 
	.B1(net54863), 
	.A2(n1021), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2131 (.ZN(n4218), 
	.B2(n1021), 
	.B1(net54859), 
	.A2(n1022), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2132 (.ZN(n1021), 
	.A(\UUT/Mpath/the_mult/x_mul_command[4] ));
   OAI22_X1 U2133 (.ZN(n4219), 
	.B2(n2752), 
	.B1(net54859), 
	.A2(n1022), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2134 (.ZN(n4220), 
	.B2(n295), 
	.B1(n5424), 
	.A2(n1023), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2135 (.ZN(n1023), 
	.A(I_DATA_INBUS[4]));
   OAI22_X1 U2136 (.ZN(n4221), 
	.B2(n2754), 
	.B1(net54859), 
	.A2(n1024), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2137 (.ZN(n4222), 
	.B2(n1024), 
	.B1(net54861), 
	.A2(n1025), 
	.A1(FE_OFN12_net54953));
   INV_X1 U2138 (.ZN(n1024), 
	.A(\UUT/Mpath/the_mult/x_mul_command[5] ));
   OAI22_X1 U2139 (.ZN(n4223), 
	.B2(n2756), 
	.B1(net54859), 
	.A2(n1025), 
	.A1(FE_OFN12_net54953));
   OAI22_X1 U2140 (.ZN(n4224), 
	.B2(n295), 
	.B1(n5423), 
	.A2(n1026), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2141 (.ZN(n1026), 
	.A(I_DATA_INBUS[5]));
   OAI22_X1 U2142 (.ZN(n4225), 
	.B2(n295), 
	.B1(n6143), 
	.A2(n1027), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2143 (.ZN(n1027), 
	.A(I_DATA_INBUS[6]));
   OAI22_X1 U2144 (.ZN(n4226), 
	.B2(n295), 
	.B1(n6094), 
	.A2(n1028), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2145 (.ZN(n1028), 
	.A(I_DATA_INBUS[7]));
   OAI22_X1 U2146 (.ZN(n4227), 
	.B2(n295), 
	.B1(n5897), 
	.A2(n1029), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2147 (.ZN(n1029), 
	.A(I_DATA_INBUS[8]));
   OAI22_X1 U2148 (.ZN(n4228), 
	.B2(n295), 
	.B1(n5889), 
	.A2(n1030), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2149 (.ZN(n1030), 
	.A(I_DATA_INBUS[9]));
   OAI22_X1 U2150 (.ZN(n4229), 
	.B2(n295), 
	.B1(n5881), 
	.A2(n1031), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2151 (.ZN(n1031), 
	.A(I_DATA_INBUS[10]));
   OAI22_X1 U2152 (.ZN(n4230), 
	.B2(n295), 
	.B1(n6036), 
	.A2(n1032), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2153 (.ZN(n1032), 
	.A(I_DATA_INBUS[11]));
   OAI22_X1 U2154 (.ZN(n4231), 
	.B2(n295), 
	.B1(n6035), 
	.A2(n1033), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2155 (.ZN(n1033), 
	.A(I_DATA_INBUS[12]));
   OAI22_X1 U2156 (.ZN(n4232), 
	.B2(n295), 
	.B1(n6033), 
	.A2(n1034), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2157 (.ZN(n1034), 
	.A(I_DATA_INBUS[13]));
   OAI22_X1 U2158 (.ZN(n4233), 
	.B2(n295), 
	.B1(n6032), 
	.A2(n1035), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2159 (.ZN(n1035), 
	.A(I_DATA_INBUS[14]));
   OAI22_X1 U2160 (.ZN(n4234), 
	.B2(n295), 
	.B1(n5831), 
	.A2(n1036), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2161 (.ZN(n1036), 
	.A(I_DATA_INBUS[15]));
   OAI22_X1 U2162 (.ZN(n4235), 
	.B2(n295), 
	.B1(n6027), 
	.A2(n1037), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2163 (.ZN(n1037), 
	.A(I_DATA_INBUS[16]));
   OAI22_X1 U2164 (.ZN(n4236), 
	.B2(n295), 
	.B1(n6034), 
	.A2(n1038), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2165 (.ZN(n1038), 
	.A(I_DATA_INBUS[17]));
   OAI22_X1 U2166 (.ZN(n4237), 
	.B2(n295), 
	.B1(n6026), 
	.A2(n1039), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2167 (.ZN(n1039), 
	.A(I_DATA_INBUS[18]));
   OAI22_X1 U2168 (.ZN(n4238), 
	.B2(n295), 
	.B1(n6031), 
	.A2(n1040), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2169 (.ZN(n1040), 
	.A(I_DATA_INBUS[19]));
   OAI22_X1 U2170 (.ZN(n4239), 
	.B2(n295), 
	.B1(n6029), 
	.A2(n1041), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2171 (.ZN(n1041), 
	.A(I_DATA_INBUS[20]));
   OAI22_X1 U2172 (.ZN(n4240), 
	.B2(n295), 
	.B1(n6037), 
	.A2(n1042), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2173 (.ZN(n1042), 
	.A(I_DATA_INBUS[21]));
   OAI22_X1 U2174 (.ZN(n4241), 
	.B2(n295), 
	.B1(n5896), 
	.A2(n1043), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2175 (.ZN(n1043), 
	.A(I_DATA_INBUS[22]));
   OAI22_X1 U2176 (.ZN(n4242), 
	.B2(n295), 
	.B1(n5888), 
	.A2(n1044), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2177 (.ZN(n1044), 
	.A(I_DATA_INBUS[23]));
   OAI22_X1 U2178 (.ZN(n4243), 
	.B2(n295), 
	.B1(n5879), 
	.A2(n1045), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2179 (.ZN(n1045), 
	.A(I_DATA_INBUS[24]));
   OAI22_X1 U2180 (.ZN(n4244), 
	.B2(n295), 
	.B1(n5871), 
	.A2(n1046), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2181 (.ZN(n1046), 
	.A(I_DATA_INBUS[25]));
   OAI21_X1 U2182 (.ZN(n4245), 
	.B2(n1047), 
	.B1(net54847), 
	.A(n1048));
   OAI21_X1 U2183 (.ZN(n1048), 
	.B2(n1050), 
	.B1(n1049), 
	.A(net54859));
   INV_X1 U2184 (.ZN(n1050), 
	.A(n1051));
   NOR3_X1 U2185 (.ZN(n1049), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1995 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2007 ), 
	.A1(n1052));
   OAI221_X1 U2186 (.ZN(n4246), 
	.C2(n1054), 
	.C1(net54891), 
	.B2(n1053), 
	.B1(FE_OFN12_net54953), 
	.A(n1055));
   AOI21_X1 U2187 (.ZN(n1053), 
	.B2(n6042), 
	.B1(n1056), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2019 ));
   OAI21_X1 U2188 (.ZN(n1056), 
	.B2(n1057), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N2001 ), 
	.A(n1058));
   NOR3_X1 U2189 (.ZN(n1057), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1995 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A1(n1052));
   INV_X1 U2190 (.ZN(n1052), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1987 ));
   OAI211_X1 U2191 (.ZN(n4247), 
	.C2(n1059), 
	.C1(net54877), 
	.B(n1055), 
	.A(n1060));
   NAND4_X1 U2192 (.ZN(n1060), 
	.A4(\UUT/Mcontrol/Operation_decoding32/N1994 ), 
	.A3(n6042), 
	.A2(net54869), 
	.A1(n1061));
   OAI22_X1 U2193 (.ZN(n4248), 
	.B2(n116), 
	.B1(FE_OFN12_net54953), 
	.A2(n2781), 
	.A1(net54847));
   AND4_X1 U2194 (.ZN(n116), 
	.A4(n1058), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1994 ), 
	.A2(n1062), 
	.A1(n1051));
   INV_X1 U2195 (.ZN(n1058), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2007 ));
   NAND3_X1 U2196 (.ZN(n1062), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1987 ));
   NOR4_X1 U2197 (.ZN(n1051), 
	.A4(\UUT/Mcontrol/Operation_decoding32/N2001 ), 
	.A3(n1064), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
	.A1(n1063));
   OAI221_X1 U2198 (.ZN(n4249), 
	.C2(n1067), 
	.C1(net54889), 
	.B2(n1066), 
	.B1(n1065), 
	.A(n1055));
   NAND2_X1 U2199 (.ZN(n1055), 
	.A2(n1063), 
	.A1(net54877));
   INV_X1 U2200 (.ZN(n1063), 
	.A(n6050));
   INV_X1 U2201 (.ZN(n1067), 
	.A(\UUT/Mcontrol/x_sampled_dmem_command[SIGN] ));
   NAND2_X1 U2202 (.ZN(n1066), 
	.A2(n6042), 
	.A1(net54875));
   AOI21_X1 U2203 (.ZN(n1065), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N2005 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N1993 ), 
	.A(\UUT/Mcontrol/d_instr [26]));
   OAI21_X1 U2204 (.ZN(n4250), 
	.B2(n2783), 
	.B1(n295), 
	.A(n1068));
   NAND2_X1 U2205 (.ZN(n1068), 
	.A2(n295), 
	.A1(I_DATA_INBUS[26]));
   OAI21_X1 U2206 (.ZN(n4251), 
	.B2(n2784), 
	.B1(n295), 
	.A(n1069));
   NAND2_X1 U2207 (.ZN(n1069), 
	.A2(n295), 
	.A1(I_DATA_INBUS[27]));
   OAI21_X1 U2208 (.ZN(n4252), 
	.B2(n2785), 
	.B1(n295), 
	.A(n1070));
   NAND2_X1 U2209 (.ZN(n1070), 
	.A2(n295), 
	.A1(I_DATA_INBUS[28]));
   OAI22_X1 U2210 (.ZN(n4253), 
	.B2(n295), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N1877 ), 
	.A2(n1071), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2211 (.ZN(n1071), 
	.A(I_DATA_INBUS[29]));
   OAI22_X1 U2212 (.ZN(n4254), 
	.B2(n295), 
	.B1(n6070), 
	.A2(n1072), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2213 (.ZN(n1072), 
	.A(I_DATA_INBUS[30]));
   OAI22_X1 U2214 (.ZN(n4255), 
	.B2(\UUT/Mcontrol/st_logic/N34 ), 
	.B1(net54863), 
	.A2(\UUT/Mpath/the_mult/N223 ), 
	.A1(FE_OFN12_net54953));
   OAI221_X1 U2216 (.ZN(n4256), 
	.C2(net54889), 
	.C1(\UUT/Mpath/the_alu/N83 ), 
	.B2(FE_OFCN207_n316), 
	.B1(n1073), 
	.A(n1074));
   AOI22_X1 U2217 (.ZN(n1074), 
	.B2(n1076), 
	.B1(FE_OFN4_n319), 
	.A2(n1075), 
	.A1(FE_OFN5_n318));
   NAND2_X1 U2220 (.ZN(n316), 
	.A2(n1077), 
	.A1(net54875));
   OAI22_X1 U2221 (.ZN(n4257), 
	.B2(n968), 
	.B1(net54863), 
	.A2(n1078), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2222 (.ZN(n968), 
	.A(\UUT/Mpath/the_mult/Mult_out[0] ));
   INV_X1 U2223 (.ZN(n1078), 
	.A(\UUT/Mpath/the_mult/x_mult_out[0] ));
   OAI22_X1 U2224 (.ZN(n4258), 
	.B2(n794), 
	.B1(net54863), 
	.A2(n1079), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2225 (.ZN(n794), 
	.A(\UUT/Mpath/the_mult/Mult_out[1] ));
   INV_X1 U2226 (.ZN(n1079), 
	.A(\UUT/Mpath/the_mult/x_mult_out[1] ));
   OAI22_X1 U2227 (.ZN(n4259), 
	.B2(n772), 
	.B1(net54863), 
	.A2(n1080), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2228 (.ZN(n772), 
	.A(\UUT/Mpath/the_mult/Mult_out[2] ));
   INV_X1 U2229 (.ZN(n1080), 
	.A(\UUT/Mpath/the_mult/x_mult_out[2] ));
   OAI22_X1 U2230 (.ZN(n4260), 
	.B2(n749), 
	.B1(net54867), 
	.A2(n1081), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2231 (.ZN(n749), 
	.A(\UUT/Mpath/the_mult/Mult_out[3] ));
   INV_X1 U2232 (.ZN(n1081), 
	.A(\UUT/Mpath/the_mult/x_mult_out[3] ));
   OAI22_X1 U2233 (.ZN(n4261), 
	.B2(n726), 
	.B1(net54863), 
	.A2(n1082), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2234 (.ZN(n726), 
	.A(\UUT/Mpath/the_mult/Mult_out[4] ));
   INV_X1 U2235 (.ZN(n1082), 
	.A(\UUT/Mpath/the_mult/x_mult_out[4] ));
   OAI22_X1 U2236 (.ZN(n4262), 
	.B2(n703), 
	.B1(net54865), 
	.A2(n1083), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2237 (.ZN(n703), 
	.A(\UUT/Mpath/the_mult/Mult_out[5] ));
   INV_X1 U2238 (.ZN(n1083), 
	.A(\UUT/Mpath/the_mult/x_mult_out[5] ));
   OAI22_X1 U2239 (.ZN(n4263), 
	.B2(n675), 
	.B1(net54863), 
	.A2(n1084), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2240 (.ZN(n675), 
	.A(\UUT/Mpath/the_mult/Mult_out[6] ));
   INV_X1 U2241 (.ZN(n1084), 
	.A(\UUT/Mpath/the_mult/x_mult_out[6] ));
   OAI22_X1 U2242 (.ZN(n4264), 
	.B2(n652), 
	.B1(net54865), 
	.A2(n1085), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2243 (.ZN(n652), 
	.A(\UUT/Mpath/the_mult/Mult_out[7] ));
   INV_X1 U2244 (.ZN(n1085), 
	.A(\UUT/Mpath/the_mult/x_mult_out[7] ));
   OAI22_X1 U2245 (.ZN(n4265), 
	.B2(n635), 
	.B1(net54865), 
	.A2(n1086), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2246 (.ZN(n635), 
	.A(\UUT/Mpath/the_mult/Mult_out[8] ));
   INV_X1 U2247 (.ZN(n1086), 
	.A(\UUT/Mpath/the_mult/x_mult_out[8] ));
   OAI22_X1 U2248 (.ZN(n4266), 
	.B2(n615), 
	.B1(net54865), 
	.A2(n1087), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2249 (.ZN(n615), 
	.A(\UUT/Mpath/the_mult/Mult_out[9] ));
   INV_X1 U2250 (.ZN(n1087), 
	.A(\UUT/Mpath/the_mult/x_mult_out[9] ));
   OAI22_X1 U2251 (.ZN(n4267), 
	.B2(n599), 
	.B1(net54865), 
	.A2(n1088), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2252 (.ZN(n599), 
	.A(\UUT/Mpath/the_mult/Mult_out[10] ));
   INV_X1 U2253 (.ZN(n1088), 
	.A(\UUT/Mpath/the_mult/x_mult_out[10] ));
   OAI22_X1 U2254 (.ZN(n4268), 
	.B2(n580), 
	.B1(net54865), 
	.A2(n1089), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2255 (.ZN(n580), 
	.A(\UUT/Mpath/the_mult/Mult_out[11] ));
   INV_X1 U2256 (.ZN(n1089), 
	.A(\UUT/Mpath/the_mult/x_mult_out[11] ));
   OAI22_X1 U2257 (.ZN(n4269), 
	.B2(n555), 
	.B1(net54865), 
	.A2(n1090), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2258 (.ZN(n555), 
	.A(\UUT/Mpath/the_mult/Mult_out[12] ));
   INV_X1 U2259 (.ZN(n1090), 
	.A(\UUT/Mpath/the_mult/x_mult_out[12] ));
   OAI22_X1 U2260 (.ZN(n4270), 
	.B2(n529), 
	.B1(net54865), 
	.A2(n1091), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2261 (.ZN(n529), 
	.A(\UUT/Mpath/the_mult/Mult_out[13] ));
   INV_X1 U2262 (.ZN(n1091), 
	.A(\UUT/Mpath/the_mult/x_mult_out[13] ));
   OAI22_X1 U2263 (.ZN(n4271), 
	.B2(n504), 
	.B1(net54865), 
	.A2(n1092), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2264 (.ZN(n504), 
	.A(\UUT/Mpath/the_mult/Mult_out[14] ));
   INV_X1 U2265 (.ZN(n1092), 
	.A(\UUT/Mpath/the_mult/x_mult_out[14] ));
   OAI22_X1 U2266 (.ZN(n4272), 
	.B2(n475), 
	.B1(net54865), 
	.A2(n1093), 
	.A1(net54953));
   INV_X1 U2267 (.ZN(n475), 
	.A(\UUT/Mpath/the_mult/Mult_out[15] ));
   INV_X1 U2268 (.ZN(n1093), 
	.A(\UUT/Mpath/the_mult/x_mult_out[15] ));
   OAI22_X1 U2269 (.ZN(n4273), 
	.B2(n454), 
	.B1(net54867), 
	.A2(n1094), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2270 (.ZN(n454), 
	.A(\UUT/Mpath/the_mult/Mult_out[16] ));
   INV_X1 U2271 (.ZN(n1094), 
	.A(\UUT/Mpath/the_mult/x_mult_out[16] ));
   OAI22_X1 U2272 (.ZN(n4274), 
	.B2(n427), 
	.B1(net54867), 
	.A2(n1095), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2273 (.ZN(n427), 
	.A(\UUT/Mpath/the_mult/Mult_out[17] ));
   INV_X1 U2274 (.ZN(n1095), 
	.A(\UUT/Mpath/the_mult/x_mult_out[17] ));
   OAI22_X1 U2275 (.ZN(n4275), 
	.B2(n405), 
	.B1(net54867), 
	.A2(n1096), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2276 (.ZN(n405), 
	.A(\UUT/Mpath/the_mult/Mult_out[18] ));
   INV_X1 U2277 (.ZN(n1096), 
	.A(\UUT/Mpath/the_mult/x_mult_out[18] ));
   OAI22_X1 U2278 (.ZN(n4276), 
	.B2(n383), 
	.B1(net54867), 
	.A2(n1097), 
	.A1(net54953));
   INV_X1 U2279 (.ZN(n383), 
	.A(\UUT/Mpath/the_mult/Mult_out[19] ));
   INV_X1 U2280 (.ZN(n1097), 
	.A(\UUT/Mpath/the_mult/x_mult_out[19] ));
   OAI22_X1 U2281 (.ZN(n4277), 
	.B2(n357), 
	.B1(net54867), 
	.A2(n1098), 
	.A1(net54953));
   INV_X1 U2282 (.ZN(n357), 
	.A(\UUT/Mpath/the_mult/Mult_out[20] ));
   INV_X1 U2283 (.ZN(n1098), 
	.A(\UUT/Mpath/the_mult/x_mult_out[20] ));
   OAI22_X1 U2284 (.ZN(n4278), 
	.B2(n336), 
	.B1(net54867), 
	.A2(n1099), 
	.A1(net54953));
   INV_X1 U2285 (.ZN(n336), 
	.A(\UUT/Mpath/the_mult/Mult_out[21] ));
   INV_X1 U2286 (.ZN(n1099), 
	.A(\UUT/Mpath/the_mult/x_mult_out[21] ));
   OAI22_X1 U2287 (.ZN(n4279), 
	.B2(n307), 
	.B1(net54867), 
	.A2(n1100), 
	.A1(net54953));
   INV_X1 U2288 (.ZN(n307), 
	.A(\UUT/Mpath/the_mult/Mult_out[22] ));
   INV_X1 U2289 (.ZN(n1100), 
	.A(\UUT/Mpath/the_mult/x_mult_out[22] ));
   OAI22_X1 U2290 (.ZN(n4280), 
	.B2(n806), 
	.B1(net54867), 
	.A2(n1101), 
	.A1(net54953));
   INV_X1 U2291 (.ZN(n806), 
	.A(\UUT/Mpath/the_mult/Mult_out[23] ));
   INV_X1 U2292 (.ZN(n1101), 
	.A(\UUT/Mpath/the_mult/x_mult_out[23] ));
   OAI22_X1 U2293 (.ZN(n4281), 
	.B2(n213), 
	.B1(net54867), 
	.A2(n1102), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2294 (.ZN(n213), 
	.A(\UUT/Mpath/the_mult/Mult_out[24] ));
   INV_X1 U2295 (.ZN(n1102), 
	.A(\UUT/Mpath/the_mult/x_mult_out[24] ));
   OAI22_X1 U2296 (.ZN(n4282), 
	.B2(n198), 
	.B1(net54867), 
	.A2(n1103), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2297 (.ZN(n198), 
	.A(\UUT/Mpath/the_mult/Mult_out[25] ));
   INV_X1 U2298 (.ZN(n1103), 
	.A(\UUT/Mpath/the_mult/x_mult_out[25] ));
   OAI22_X1 U2299 (.ZN(n4283), 
	.B2(n185), 
	.B1(net54869), 
	.A2(n1104), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2300 (.ZN(n185), 
	.A(\UUT/Mpath/the_mult/Mult_out[26] ));
   INV_X1 U2301 (.ZN(n1104), 
	.A(\UUT/Mpath/the_mult/x_mult_out[26] ));
   OAI22_X1 U2302 (.ZN(n4284), 
	.B2(n169), 
	.B1(net54869), 
	.A2(n1105), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2303 (.ZN(n169), 
	.A(\UUT/Mpath/the_mult/Mult_out[27] ));
   INV_X1 U2304 (.ZN(n1105), 
	.A(\UUT/Mpath/the_mult/x_mult_out[27] ));
   OAI22_X1 U2305 (.ZN(n4285), 
	.B2(n157), 
	.B1(net54869), 
	.A2(n1106), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2306 (.ZN(n157), 
	.A(\UUT/Mpath/the_mult/Mult_out[28] ));
   INV_X1 U2307 (.ZN(n1106), 
	.A(\UUT/Mpath/the_mult/x_mult_out[28] ));
   OAI22_X1 U2308 (.ZN(n4286), 
	.B2(n141), 
	.B1(net54869), 
	.A2(n1107), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2309 (.ZN(n141), 
	.A(\UUT/Mpath/the_mult/Mult_out[29] ));
   INV_X1 U2310 (.ZN(n1107), 
	.A(\UUT/Mpath/the_mult/x_mult_out[29] ));
   OAI22_X1 U2311 (.ZN(n4287), 
	.B2(n864), 
	.B1(net54869), 
	.A2(n1108), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2312 (.ZN(n864), 
	.A(\UUT/Mpath/the_mult/Mult_out[30] ));
   INV_X1 U2313 (.ZN(n1108), 
	.A(\UUT/Mpath/the_mult/x_mult_out[30] ));
   OAI22_X1 U2314 (.ZN(n4288), 
	.B2(n946), 
	.B1(net54869), 
	.A2(n1109), 
	.A1(FE_OFN10_net54953));
   INV_X1 U2315 (.ZN(n946), 
	.A(\UUT/Mpath/the_mult/Mult_out[31] ));
   INV_X1 U2316 (.ZN(n1109), 
	.A(\UUT/Mpath/the_mult/x_mult_out[31] ));
   OAI21_X1 U2317 (.ZN(n4289), 
	.B2(n1110), 
	.B1(net54847), 
	.A(n1111));
   NAND2_X1 U2318 (.ZN(n1111), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[32] ));
   OAI21_X1 U2319 (.ZN(n4290), 
	.B2(n791), 
	.B1(net54847), 
	.A(n1112));
   NAND2_X1 U2320 (.ZN(n1112), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[33] ));
   INV_X1 U2321 (.ZN(n791), 
	.A(\UUT/Mpath/the_mult/Mult_out[33] ));
   OAI21_X1 U2322 (.ZN(n4291), 
	.B2(n769), 
	.B1(net54847), 
	.A(n1113));
   NAND2_X1 U2323 (.ZN(n1113), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[34] ));
   INV_X1 U2324 (.ZN(n769), 
	.A(\UUT/Mpath/the_mult/Mult_out[34] ));
   OAI21_X1 U2325 (.ZN(n4292), 
	.B2(n746), 
	.B1(net54847), 
	.A(n1114));
   NAND2_X1 U2326 (.ZN(n1114), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[35] ));
   INV_X1 U2327 (.ZN(n746), 
	.A(\UUT/Mpath/the_mult/Mult_out[35] ));
   OAI21_X1 U2328 (.ZN(n4293), 
	.B2(n723), 
	.B1(net54847), 
	.A(n1115));
   NAND2_X1 U2329 (.ZN(n1115), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[36] ));
   INV_X1 U2330 (.ZN(n723), 
	.A(\UUT/Mpath/the_mult/Mult_out[36] ));
   OAI21_X1 U2331 (.ZN(n4294), 
	.B2(n700), 
	.B1(net54849), 
	.A(n1116));
   NAND2_X1 U2332 (.ZN(n1116), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[37] ));
   INV_X1 U2333 (.ZN(n700), 
	.A(\UUT/Mpath/the_mult/Mult_out[37] ));
   OAI21_X1 U2334 (.ZN(n4295), 
	.B2(n672), 
	.B1(net54849), 
	.A(n1117));
   NAND2_X1 U2335 (.ZN(n1117), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[38] ));
   INV_X1 U2336 (.ZN(n672), 
	.A(\UUT/Mpath/the_mult/Mult_out[38] ));
   OAI21_X1 U2337 (.ZN(n4296), 
	.B2(n649), 
	.B1(net54849), 
	.A(n1118));
   NAND2_X1 U2338 (.ZN(n1118), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[39] ));
   INV_X1 U2339 (.ZN(n649), 
	.A(\UUT/Mpath/the_mult/Mult_out[39] ));
   OAI21_X1 U2340 (.ZN(n4297), 
	.B2(n632), 
	.B1(net54849), 
	.A(n1119));
   NAND2_X1 U2341 (.ZN(n1119), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[40] ));
   INV_X1 U2342 (.ZN(n632), 
	.A(\UUT/Mpath/the_mult/Mult_out[40] ));
   OAI21_X1 U2343 (.ZN(n4298), 
	.B2(n612), 
	.B1(net54849), 
	.A(n1120));
   NAND2_X1 U2344 (.ZN(n1120), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[41] ));
   INV_X1 U2345 (.ZN(n612), 
	.A(\UUT/Mpath/the_mult/Mult_out[41] ));
   OAI21_X1 U2346 (.ZN(n4299), 
	.B2(n596), 
	.B1(net54849), 
	.A(n1121));
   NAND2_X1 U2347 (.ZN(n1121), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[42] ));
   INV_X1 U2348 (.ZN(n596), 
	.A(\UUT/Mpath/the_mult/Mult_out[42] ));
   OAI21_X1 U2349 (.ZN(n4300), 
	.B2(n577), 
	.B1(net54849), 
	.A(n1122));
   NAND2_X1 U2350 (.ZN(n1122), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[43] ));
   INV_X1 U2351 (.ZN(n577), 
	.A(\UUT/Mpath/the_mult/Mult_out[43] ));
   OAI21_X1 U2352 (.ZN(n4301), 
	.B2(n552), 
	.B1(net54849), 
	.A(n1123));
   NAND2_X1 U2353 (.ZN(n1123), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[44] ));
   INV_X1 U2354 (.ZN(n552), 
	.A(\UUT/Mpath/the_mult/Mult_out[44] ));
   OAI21_X1 U2355 (.ZN(n4302), 
	.B2(n526), 
	.B1(net54849), 
	.A(n1124));
   NAND2_X1 U2356 (.ZN(n1124), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[45] ));
   INV_X1 U2357 (.ZN(n526), 
	.A(\UUT/Mpath/the_mult/Mult_out[45] ));
   OAI21_X1 U2358 (.ZN(n4303), 
	.B2(n501), 
	.B1(net54851), 
	.A(n1125));
   NAND2_X1 U2359 (.ZN(n1125), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[46] ));
   INV_X1 U2360 (.ZN(n501), 
	.A(\UUT/Mpath/the_mult/Mult_out[46] ));
   OAI21_X1 U2361 (.ZN(n4304), 
	.B2(n472), 
	.B1(net54851), 
	.A(n1126));
   NAND2_X1 U2362 (.ZN(n1126), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[47] ));
   INV_X1 U2363 (.ZN(n472), 
	.A(\UUT/Mpath/the_mult/Mult_out[47] ));
   OAI21_X1 U2364 (.ZN(n4305), 
	.B2(n451), 
	.B1(net54851), 
	.A(n1127));
   NAND2_X1 U2365 (.ZN(n1127), 
	.A2(net54853), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[48] ));
   INV_X1 U2366 (.ZN(n451), 
	.A(\UUT/Mpath/the_mult/Mult_out[48] ));
   OAI21_X1 U2367 (.ZN(n4306), 
	.B2(n424), 
	.B1(net54849), 
	.A(n1128));
   NAND2_X1 U2368 (.ZN(n1128), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[49] ));
   INV_X1 U2369 (.ZN(n424), 
	.A(\UUT/Mpath/the_mult/Mult_out[49] ));
   OAI21_X1 U2370 (.ZN(n4307), 
	.B2(n402), 
	.B1(net54851), 
	.A(n1129));
   NAND2_X1 U2371 (.ZN(n1129), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[50] ));
   INV_X1 U2372 (.ZN(n402), 
	.A(\UUT/Mpath/the_mult/Mult_out[50] ));
   OAI21_X1 U2373 (.ZN(n4308), 
	.B2(n380), 
	.B1(net54851), 
	.A(n1130));
   NAND2_X1 U2374 (.ZN(n1130), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[51] ));
   INV_X1 U2375 (.ZN(n380), 
	.A(\UUT/Mpath/the_mult/Mult_out[51] ));
   OAI21_X1 U2376 (.ZN(n4309), 
	.B2(n354), 
	.B1(net54851), 
	.A(n1131));
   NAND2_X1 U2377 (.ZN(n1131), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[52] ));
   INV_X1 U2378 (.ZN(n354), 
	.A(\UUT/Mpath/the_mult/Mult_out[52] ));
   OAI21_X1 U2379 (.ZN(n4310), 
	.B2(n333), 
	.B1(net54851), 
	.A(n1132));
   NAND2_X1 U2380 (.ZN(n1132), 
	.A2(net54855), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[53] ));
   INV_X1 U2381 (.ZN(n333), 
	.A(\UUT/Mpath/the_mult/Mult_out[53] ));
   OAI21_X1 U2382 (.ZN(n4311), 
	.B2(n304), 
	.B1(net54849), 
	.A(n1133));
   NAND2_X1 U2383 (.ZN(n1133), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[54] ));
   INV_X1 U2384 (.ZN(n304), 
	.A(\UUT/Mpath/the_mult/Mult_out[54] ));
   OAI21_X1 U2385 (.ZN(n4312), 
	.B2(n803), 
	.B1(net54851), 
	.A(n1134));
   NAND2_X1 U2386 (.ZN(n1134), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[55] ));
   INV_X1 U2387 (.ZN(n803), 
	.A(\UUT/Mpath/the_mult/Mult_out[55] ));
   OAI21_X1 U2388 (.ZN(n4313), 
	.B2(n210), 
	.B1(net54851), 
	.A(n1135));
   NAND2_X1 U2389 (.ZN(n1135), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[56] ));
   INV_X1 U2390 (.ZN(n210), 
	.A(\UUT/Mpath/the_mult/Mult_out[56] ));
   OAI21_X1 U2391 (.ZN(n4314), 
	.B2(n195), 
	.B1(net54851), 
	.A(n1136));
   NAND2_X1 U2392 (.ZN(n1136), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[57] ));
   INV_X1 U2393 (.ZN(n195), 
	.A(\UUT/Mpath/the_mult/Mult_out[57] ));
   OAI21_X1 U2394 (.ZN(n4315), 
	.B2(n182), 
	.B1(net54851), 
	.A(n1137));
   NAND2_X1 U2395 (.ZN(n1137), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[58] ));
   INV_X1 U2396 (.ZN(n182), 
	.A(\UUT/Mpath/the_mult/Mult_out[58] ));
   OAI21_X1 U2397 (.ZN(n4316), 
	.B2(n166), 
	.B1(net54853), 
	.A(n1138));
   NAND2_X1 U2398 (.ZN(n1138), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[59] ));
   INV_X1 U2399 (.ZN(n166), 
	.A(\UUT/Mpath/the_mult/Mult_out[59] ));
   OAI21_X1 U2400 (.ZN(n4317), 
	.B2(n154), 
	.B1(net54849), 
	.A(n1139));
   NAND2_X1 U2401 (.ZN(n1139), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[60] ));
   INV_X1 U2402 (.ZN(n154), 
	.A(\UUT/Mpath/the_mult/Mult_out[60] ));
   OAI21_X1 U2403 (.ZN(n4318), 
	.B2(n134), 
	.B1(net54853), 
	.A(n1140));
   NAND2_X1 U2404 (.ZN(n1140), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[61] ));
   INV_X1 U2405 (.ZN(n134), 
	.A(\UUT/Mpath/the_mult/Mult_out[61] ));
   OAI21_X1 U2406 (.ZN(n4319), 
	.B2(n861), 
	.B1(net54853), 
	.A(n1141));
   NAND2_X1 U2407 (.ZN(n1141), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[62] ));
   INV_X1 U2408 (.ZN(n861), 
	.A(\UUT/Mpath/the_mult/Mult_out[62] ));
   OAI21_X1 U2409 (.ZN(n4320), 
	.B2(n1142), 
	.B1(net54851), 
	.A(n1143));
   NAND2_X1 U2410 (.ZN(n1143), 
	.A2(net54857), 
	.A1(\UUT/Mpath/the_mult/x_mult_out[63] ));
   OAI22_X1 U2411 (.ZN(n4321), 
	.B2(FE_OFN12_net54953), 
	.B1(n1073), 
	.A2(net54879), 
	.A1(n5527));
   OAI22_X1 U2412 (.ZN(n4322), 
	.B2(net54875), 
	.B1(\UUT/Mpath/the_memhandle/N240 ), 
	.A2(FE_OFN11_net54953), 
	.A1(n1144));
   INV_X1 U2413 (.ZN(n1144), 
	.A(\UUT/daddr_out [0]));
   OAI222_X1 U2414 (.ZN(n4324), 
	.C2(net54893), 
	.C1(\UUT/Mpath/the_alu/N68 ), 
	.B2(n300), 
	.B1(n79), 
	.A2(n123), 
	.A1(n80));
   INV_X1 U2415 (.ZN(n79), 
	.A(\UUT/break_code[8] ));
   INV_X1 U2416 (.ZN(n80), 
	.A(n1145));
   OAI222_X1 U2417 (.ZN(n1145), 
	.C2(n132), 
	.C1(n5436), 
	.B2(n131), 
	.B1(n958), 
	.A2(n129), 
	.A1(n638));
   OAI211_X1 U2419 (.ZN(n641), 
	.C2(n482), 
	.C1(n1146), 
	.B(n1147), 
	.A(n484));
   AOI22_X1 U2420 (.ZN(n1147), 
	.B2(n489), 
	.B1(n1149), 
	.A2(n1148), 
	.A1(n486));
   INV_X1 U2421 (.ZN(n1149), 
	.A(n5437));
   INV_X1 U2422 (.ZN(n1146), 
	.A(n5747));
   INV_X1 U2423 (.ZN(n638), 
	.A(n1150));
   OAI211_X1 U2424 (.ZN(n1150), 
	.C2(n321), 
	.C1(n5616), 
	.B(n1152), 
	.A(n1151));
   AOI222_X1 U2425 (.ZN(n1152), 
	.C2(n1154), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[8] ), 
	.A2(n1153), 
	.A1(FE_OFN91_n285));
   INV_X1 U2426 (.ZN(n1154), 
	.A(n5679));
   AOI22_X1 U2427 (.ZN(n1151), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[8] ), 
	.A2(n6190), 
	.A1(FE_OFN89_n290));
   OAI222_X1 U2428 (.ZN(n4325), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N64 ), 
	.B2(n300), 
	.B1(n76), 
	.A2(n123), 
	.A1(n77));
   INV_X1 U2429 (.ZN(n76), 
	.A(\UUT/break_code[10] ));
   INV_X1 U2430 (.ZN(n77), 
	.A(n1155));
   OAI222_X1 U2431 (.ZN(n1155), 
	.C2(n132), 
	.C1(n5523), 
	.B2(n131), 
	.B1(n959), 
	.A2(n129), 
	.A1(n602));
   OAI211_X1 U2433 (.ZN(n605), 
	.C2(n1156), 
	.C1(n482), 
	.B(n1157), 
	.A(n484));
   AOI22_X1 U2434 (.ZN(n1157), 
	.B2(n489), 
	.B1(n1158), 
	.A2(n781), 
	.A1(n486));
   INV_X1 U2435 (.ZN(n1158), 
	.A(n5524));
   INV_X1 U2436 (.ZN(n781), 
	.A(n5845));
   AND2_X1 U2437 (.ZN(n486), 
	.A2(n5710), 
	.A1(n5713));
   INV_X1 U2438 (.ZN(n1156), 
	.A(n5838));
   NAND2_X1 U2439 (.ZN(n482), 
	.A2(n5710), 
	.A1(n5711));
   INV_X1 U2440 (.ZN(n602), 
	.A(n1159));
   OAI211_X1 U2441 (.ZN(n1159), 
	.C2(n321), 
	.C1(n5674), 
	.B(n1161), 
	.A(n1160));
   AOI222_X1 U2442 (.ZN(n1161), 
	.C2(n1163), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[10] ), 
	.A2(n1162), 
	.A1(FE_OFN91_n285));
   INV_X1 U2443 (.ZN(n1163), 
	.A(n5708));
   AOI22_X1 U2444 (.ZN(n1160), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[10] ), 
	.A2(n6205), 
	.A1(FE_OFN89_n290));
   OAI22_X1 U2445 (.ZN(n4327), 
	.B2(n74), 
	.B1(net54953), 
	.A2(net54877), 
	.A1(\UUT/Mpath/the_alu/N22 ));
   INV_X1 U2446 (.ZN(n74), 
	.A(n1164));
   OAI211_X1 U2447 (.ZN(n1164), 
	.C2(n115), 
	.C1(n789), 
	.B(n1165), 
	.A(n856));
   NOR2_X1 U2448 (.ZN(n1165), 
	.A2(n1166), 
	.A1(n854));
   NOR3_X1 U2449 (.ZN(n1166), 
	.A3(n1167), 
	.A2(n5831), 
	.A1(n450));
   AND2_X1 U2450 (.ZN(n854), 
	.A2(n207), 
	.A1(n5869));
   AOI21_X1 U2451 (.ZN(n856), 
	.B2(n207), 
	.B1(n5870), 
	.A(n448));
   NOR2_X1 U2452 (.ZN(n207), 
	.A2(n1168), 
	.A1(n450));
   OR2_X1 U2453 (.ZN(n450), 
	.A2(n175), 
	.A1(n1169));
   INV_X1 U2454 (.ZN(n115), 
	.A(n1170));
   OAI222_X1 U2455 (.ZN(n1170), 
	.C2(n132), 
	.C1(n5454), 
	.B2(n131), 
	.B1(n952), 
	.A2(n129), 
	.A1(FE_OFN13_n953));
   AND2_X1 U2458 (.ZN(n282), 
	.A2(n1172), 
	.A1(n484));
   NAND2_X1 U2459 (.ZN(n1172), 
	.A2(n5710), 
	.A1(n5945));
   NAND2_X1 U2460 (.ZN(n484), 
	.A2(n5710), 
	.A1(n5715));
   NAND3_X1 U2461 (.ZN(n281), 
	.A3(n5951), 
	.A2(n5710), 
	.A1(n5950));
   INV_X1 U2462 (.ZN(n789), 
	.A(n175));
   OAI22_X1 U2463 (.ZN(n4328), 
	.B2(FE_OFN13_n953), 
	.B1(FE_OFN12_net54953), 
	.A2(net54877), 
	.A1(n5455));
   AOI221_X1 U2464 (.ZN(n953), 
	.C2(FE_OFN91_n285), 
	.C1(n6197), 
	.B2(n284), 
	.B1(n1173), 
	.A(n1174));
   INV_X1 U2465 (.ZN(n1174), 
	.A(n1175));
   AOI222_X1 U2466 (.ZN(n1175), 
	.C2(n291), 
	.C1(\UUT/Mpath/the_mult/x_mult_out[31] ), 
	.B2(n6644), 
	.B1(FE_OFN89_n290), 
	.A2(n1176), 
	.A1(n288));
   INV_X1 U2467 (.ZN(n1176), 
	.A(n5628));
   INV_X1 U2468 (.ZN(n288), 
	.A(n321));
   INV_X1 U2469 (.ZN(n1173), 
	.A(n5685));
   INV_X1 U2472 (.ZN(n948), 
	.A(n5629));
   INV_X1 U2473 (.ZN(n1142), 
	.A(\UUT/Mpath/the_mult/Mult_out[63] ));
   OAI221_X1 U2474 (.ZN(n4330), 
	.C2(n135), 
	.C1(n5709), 
	.B2(n1110), 
	.B1(n133), 
	.A(n1178));
   AOI22_X1 U2475 (.ZN(n1178), 
	.B2(n139), 
	.B1(\UUT/Mpath/the_mult/Mad_out [32]), 
	.A2(n970), 
	.A1(n137));
   INV_X1 U2478 (.ZN(n970), 
	.A(n5677));
   INV_X1 U2485 (.ZN(n1110), 
	.A(\UUT/Mpath/the_mult/Mult_out[32] ));
   AND2_X1 U2487 (.ZN(n975), 
	.A2(net54895), 
	.A1(n5413));
   OAI22_X1 U2488 (.ZN(n4331), 
	.B2(net54875), 
	.B1(n5677), 
	.A2(n1184), 
	.A1(FE_OFN10_net54953));
   OAI221_X1 U2489 (.ZN(n4332), 
	.C2(n1184), 
	.C1(n147), 
	.B2(n310), 
	.B1(n1073), 
	.A(n1185));
   AOI22_X1 U2490 (.ZN(n1185), 
	.B2(n1076), 
	.B1(FE_OFN6_n314), 
	.A2(n1075), 
	.A1(FE_OFCN208_FE_OFN7_n312));
   INV_X1 U2493 (.ZN(n1184), 
	.A(\UUT/Mpath/the_mult/x_operand1[0] ));
   NAND2_X2 U2494 (.ZN(n310), 
	.A2(n1077), 
	.A1(n147));
   INV_X1 U2495 (.ZN(n1077), 
	.A(n5528));
   OAI21_X1 U2497 (.ZN(n73), 
	.B2(\UUT/Mpath/the_mult/N223 ), 
	.B1(\UUT/Mpath/the_mult/N227 ), 
	.A(net54859));
   OAI22_X1 U2498 (.ZN(n4333), 
	.B2(n945), 
	.B1(n6069), 
	.A2(\UUT/Mpath/N111 ), 
	.A1(net54847));
   NAND2_X1 U2499 (.ZN(n945), 
	.A2(net54857), 
	.A1(n1186));
   NAND4_X1 U2500 (.ZN(n1186), 
	.A4(n937), 
	.A3(n931), 
	.A2(n935), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2025 ));
   OAI22_X1 U2501 (.ZN(n4334), 
	.B2(n295), 
	.B1(n6069), 
	.A2(n1187), 
	.A1(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U2503 (.ZN(n1187), 
	.A(I_DATA_INBUS[31]));
   INV_X1 U2505 (.ZN(n978), 
	.A(\UUT/Mcontrol/st_logic/N10 ));
   OAI222_X1 U2506 (.ZN(n4335), 
	.C2(net54895), 
	.C1(\UUT/Mpath/the_alu/N84 ), 
	.B2(n300), 
	.B1(n68), 
	.A2(n123), 
	.A1(n70));
   INV_X1 U2507 (.ZN(n300), 
	.A(n449));
   NOR2_X1 U2508 (.ZN(n449), 
	.A2(FE_OFN12_net54953), 
	.A1(n175));
   INV_X1 U2510 (.ZN(n68), 
	.A(\UUT/break_code[0] ));
   NAND2_X2 U2511 (.ZN(n123), 
	.A2(net54859), 
	.A1(n175));
   OAI21_X2 U2512 (.ZN(n175), 
	.B2(n6170), 
	.B1(n6206), 
	.A(n6030));
   INV_X1 U2513 (.ZN(n70), 
	.A(n1188));
   OAI222_X1 U2514 (.ZN(n1188), 
	.C2(n129), 
	.C1(n1073), 
	.B2(n131), 
	.B1(n960), 
	.A2(n132), 
	.A1(n5526));
   INV_X1 U2516 (.ZN(n1073), 
	.A(n1189));
   OAI211_X1 U2517 (.ZN(n1189), 
	.C2(n321), 
	.C1(n5676), 
	.B(n1191), 
	.A(n1190));
   AOI222_X1 U2518 (.ZN(n1191), 
	.C2(n1192), 
	.C1(n284), 
	.B2(FE_OFN90_n325), 
	.B1(\UUT/Mpath/out_jar[0] ), 
	.A2(n5613), 
	.A1(FE_OFN91_n285));
   INV_X1 U2519 (.ZN(n1192), 
	.A(n5709));
   INV_X1 U2521 (.ZN(n1193), 
	.A(n1194));
   AOI22_X1 U2523 (.ZN(n1190), 
	.B2(n291), 
	.B1(\UUT/Mpath/the_mult/x_mult_out[0] ), 
	.A2(\UUT/daddr_out [0]), 
	.A1(FE_OFN89_n290));
   NOR3_X1 U2525 (.ZN(n290), 
	.A3(\UUT/Mpath/N115 ), 
	.A2(FE_OFN91_n285), 
	.A1(n1195));
   INV_X1 U2527 (.ZN(n1195), 
	.A(\UUT/Mpath/N125 ));
   NAND3_X2 U2528 (.ZN(n321), 
	.A3(\UUT/Mpath/the_mult/N216 ), 
	.A2(n1197), 
	.A1(n1194));
   INV_X1 U2529 (.ZN(n1197), 
	.A(\UUT/Mpath/the_mult/N198 ));
   NOR2_X1 U2530 (.ZN(n1194), 
	.A2(\UUT/Mpath/N125 ), 
	.A1(FE_OFN91_n285));
   OAI211_X1 U2534 (.ZN(n1076), 
	.C2(n5527), 
	.C1(n5710), 
	.B(n1199), 
	.A(n1198));
   AOI222_X1 U2535 (.ZN(n1199), 
	.C2(n686), 
	.C1(n6000), 
	.B2(n1148), 
	.B1(n685), 
	.A2(n684), 
	.A1(n5747));
   AND2_X1 U2536 (.ZN(n686), 
	.A2(\UUT/Mpath/the_memhandle/N37 ), 
	.A1(n687));
   INV_X1 U2537 (.ZN(n1148), 
	.A(n5999));
   AND2_X1 U2538 (.ZN(n685), 
	.A2(n688), 
	.A1(n5757));
   AND2_X1 U2539 (.ZN(n684), 
	.A2(n1200), 
	.A1(n5710));
   OAI22_X1 U2540 (.ZN(n1200), 
	.B2(n1202), 
	.B1(\UUT/Mpath/the_memhandle/N34 ), 
	.A2(n1201), 
	.A1(n5985));
   INV_X1 U2541 (.ZN(n1202), 
	.A(n5755));
   AOI22_X1 U2542 (.ZN(n1198), 
	.B2(n688), 
	.B1(n5994), 
	.A2(n687), 
	.A1(n6001));
   INV_X1 U2543 (.ZN(n688), 
	.A(n660));
   NAND2_X1 U2544 (.ZN(n660), 
	.A2(n1201), 
	.A1(n5710));
   NOR2_X1 U2545 (.ZN(n687), 
	.A2(n489), 
	.A1(n1201));
   INV_X1 U2546 (.ZN(n489), 
	.A(n5710));
   INV_X1 U2547 (.ZN(n1201), 
	.A(\UUT/Mpath/the_memhandle/N34 ));
   NAND2_X1 U2549 (.ZN(n6197), 
	.A2(n1204), 
	.A1(n1203));
   AOI222_X1 U2550 (.ZN(n1204), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [31]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [31]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [31]));
   AOI22_X1 U2551 (.ZN(n1203), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [31]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [31]));
   INV_X1 U2554 (.ZN(n1209), 
	.A(\UUT/Mpath/the_alu/N21 ));
   AOI22_X1 U2555 (.ZN(n1206), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N94 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N126 ));
   AOI22_X1 U2556 (.ZN(n1205), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N190 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N158 ));
   INV_X1 U2557 (.ZN(n6116), 
	.A(n1216));
   NOR4_X1 U2558 (.ZN(n6076), 
	.A4(n6079), 
	.A3(n6067), 
	.A2(n1008), 
	.A1(n1217));
   INV_X1 U2559 (.ZN(n1008), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1945 ));
   INV_X1 U2560 (.ZN(n1217), 
	.A(n6285));
   NAND3_X1 U2561 (.ZN(n6074), 
	.A3(n857), 
	.A2(n445), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1975 ));
   INV_X1 U2562 (.ZN(n6073), 
	.A(n937));
   NOR2_X1 U2563 (.ZN(n937), 
	.A2(n1219), 
	.A1(n1218));
   INV_X1 U2564 (.ZN(n1218), 
	.A(n932));
   INV_X1 U2566 (.ZN(n6070), 
	.A(\UUT/Mcontrol/d_sampled_finstr [30]));
   INV_X1 U2567 (.ZN(n6069), 
	.A(\UUT/Mcontrol/d_sampled_finstr [31]));
   INV_X1 U2568 (.ZN(n6051), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2019 ));
   INV_X1 U2570 (.ZN(n6048), 
	.A(n6078));
   INV_X1 U2571 (.ZN(n6037), 
	.A(\UUT/Mcontrol/d_sampled_finstr [21]));
   INV_X1 U2572 (.ZN(n6034), 
	.A(\UUT/Mcontrol/d_sampled_finstr [17]));
   INV_X1 U2573 (.ZN(n6031), 
	.A(\UUT/Mcontrol/d_sampled_finstr [19]));
   INV_X1 U2574 (.ZN(n6029), 
	.A(\UUT/Mcontrol/d_sampled_finstr [20]));
   INV_X1 U2575 (.ZN(n6028), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2043 ));
   INV_X1 U2576 (.ZN(n6027), 
	.A(\UUT/Mcontrol/d_sampled_finstr [16]));
   INV_X1 U2577 (.ZN(n6026), 
	.A(\UUT/Mcontrol/d_sampled_finstr [18]));
   AOI22_X1 U2578 (.ZN(n5944), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[16]), 
	.A2(n5779), 
	.A1(dram_data_inbus[16]));
   AOI22_X1 U2579 (.ZN(n5919), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[17]), 
	.A2(n5779), 
	.A1(dram_data_inbus[17]));
   INV_X1 U2580 (.ZN(n5896), 
	.A(\UUT/Mcontrol/d_sampled_finstr [22]));
   AOI22_X1 U2581 (.ZN(n5890), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[24]), 
	.A2(n5779), 
	.A1(dram_data_inbus[24]));
   INV_X1 U2582 (.ZN(n5888), 
	.A(\UUT/Mcontrol/d_sampled_finstr [23]));
   AOI22_X1 U2583 (.ZN(n5882), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[25]), 
	.A2(n5779), 
	.A1(dram_data_inbus[25]));
   INV_X1 U2584 (.ZN(n5880), 
	.A(n5870));
   INV_X1 U2585 (.ZN(n5879), 
	.A(\UUT/Mcontrol/d_sampled_finstr [24]));
   AOI22_X1 U2586 (.ZN(n5873), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[26]), 
	.A2(n5779), 
	.A1(dram_data_inbus[26]));
   NAND2_X1 U2587 (.ZN(n5872), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A1(n1220));
   INV_X1 U2588 (.ZN(n1220), 
	.A(n6118));
   INV_X1 U2589 (.ZN(n5871), 
	.A(\UUT/Mcontrol/d_sampled_finstr [25]));
   AOI22_X1 U2590 (.ZN(n5863), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[27]), 
	.A2(n5779), 
	.A1(dram_data_inbus[27]));
   AOI22_X1 U2591 (.ZN(n5857), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[28]), 
	.A2(n5779), 
	.A1(dram_data_inbus[28]));
   AOI22_X1 U2592 (.ZN(n5851), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[29]), 
	.A2(n5779), 
	.A1(dram_data_inbus[29]));
   AOI22_X1 U2593 (.ZN(n5841), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[18]), 
	.A2(n5779), 
	.A1(dram_data_inbus[18]));
   AOI22_X1 U2594 (.ZN(n5832), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[30]), 
	.A2(n5779), 
	.A1(dram_data_inbus[30]));
   AOI22_X1 U2595 (.ZN(n5825), 
	.B2(BUS_DATA_INBUS[31]), 
	.B1(FE_OFN92_n5780), 
	.A2(dram_data_inbus[31]), 
	.A1(n5779));
   AOI22_X1 U2596 (.ZN(n5815), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[19]), 
	.A2(n5779), 
	.A1(dram_data_inbus[19]));
   AOI22_X1 U2597 (.ZN(n5802), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[20]), 
	.A2(n5779), 
	.A1(dram_data_inbus[20]));
   AOI22_X1 U2598 (.ZN(n5789), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[21]), 
	.A2(n5779), 
	.A1(dram_data_inbus[21]));
   AOI22_X1 U2599 (.ZN(n5772), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[22]), 
	.A2(n5779), 
	.A1(dram_data_inbus[22]));
   AOI22_X1 U2600 (.ZN(n5760), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[23]), 
	.A2(n5779), 
	.A1(dram_data_inbus[23]));
   OAI21_X1 U2601 (.ZN(n5754), 
	.B2(n5983), 
	.B1(n5984), 
	.A(\UUT/Mpath/the_memhandle/N34 ));
   NAND2_X1 U2602 (.ZN(n5613), 
	.A2(n1222), 
	.A1(n1221));
   AOI222_X1 U2603 (.ZN(n1222), 
	.C2(\UUT/Mpath/the_shift/sh_rol [0]), 
	.C1(n6199), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [0]), 
	.A2(\UUT/Mpath/the_shift/sh_ror [0]), 
	.A1(FE_OFN88_n6201));
   AOI22_X1 U2604 (.ZN(n1221), 
	.B2(\UUT/Mpath/the_shift/sh_sra [0]), 
	.B1(n6198), 
	.A2(\UUT/Mpath/the_shift/sh_sll [0]), 
	.A1(n6200));
   NAND3_X1 U2605 (.ZN(n5606), 
	.A3(n1225), 
	.A2(n1224), 
	.A1(n1223));
   AOI222_X1 U2606 (.ZN(n1225), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[24] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[24] ), 
	.A2(n1226), 
	.A1(n1208));
   INV_X1 U2607 (.ZN(n1226), 
	.A(\UUT/Mpath/the_alu/N35 ));
   AOI22_X1 U2608 (.ZN(n1224), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N101 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N133 ));
   AOI22_X1 U2609 (.ZN(n1223), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N197 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N165 ));
   NAND2_X1 U2610 (.ZN(n5605), 
	.A2(n1228), 
	.A1(n1227));
   AOI222_X1 U2611 (.ZN(n1228), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [24]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [24]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [24]));
   AOI22_X1 U2612 (.ZN(n1227), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [24]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [24]));
   NAND3_X1 U2613 (.ZN(n5599), 
	.A3(n1231), 
	.A2(n1230), 
	.A1(n1229));
   AOI222_X1 U2614 (.ZN(n1231), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[25] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[25] ), 
	.A2(n1232), 
	.A1(n1208));
   INV_X1 U2615 (.ZN(n1232), 
	.A(\UUT/Mpath/the_alu/N33 ));
   AOI22_X1 U2616 (.ZN(n1230), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N100 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N132 ));
   AOI22_X1 U2617 (.ZN(n1229), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N196 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N164 ));
   NAND2_X1 U2618 (.ZN(n5598), 
	.A2(n1234), 
	.A1(n1233));
   AOI222_X1 U2619 (.ZN(n1234), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [25]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [25]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [25]));
   AOI22_X1 U2620 (.ZN(n1233), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [25]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [25]));
   INV_X1 U2623 (.ZN(n1238), 
	.A(\UUT/Mpath/the_alu/N31 ));
   AOI22_X1 U2624 (.ZN(n1236), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N99 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N131 ));
   AOI22_X1 U2625 (.ZN(n1235), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N195 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N163 ));
   NAND2_X1 U2626 (.ZN(n5591), 
	.A2(n1240), 
	.A1(n1239));
   AOI222_X1 U2627 (.ZN(n1240), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [26]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [26]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [26]));
   AOI22_X1 U2628 (.ZN(n1239), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [26]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [26]));
   INV_X1 U2631 (.ZN(n1244), 
	.A(\UUT/Mpath/the_alu/N29 ));
   AOI22_X1 U2632 (.ZN(n1242), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N98 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N130 ));
   AOI22_X1 U2633 (.ZN(n1241), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N194 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N162 ));
   NAND2_X1 U2634 (.ZN(n5584), 
	.A2(n1246), 
	.A1(n1245));
   AOI222_X1 U2635 (.ZN(n1246), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [27]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [27]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [27]));
   AOI22_X1 U2636 (.ZN(n1245), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [27]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [27]));
   INV_X1 U2639 (.ZN(n1250), 
	.A(\UUT/Mpath/the_alu/N27 ));
   AOI22_X1 U2640 (.ZN(n1248), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N97 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N129 ));
   AOI22_X1 U2641 (.ZN(n1247), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N193 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N161 ));
   NAND2_X1 U2642 (.ZN(n5577), 
	.A2(n1252), 
	.A1(n1251));
   AOI222_X1 U2643 (.ZN(n1252), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [28]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [28]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [28]));
   AOI22_X1 U2644 (.ZN(n1251), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [28]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [28]));
   INV_X1 U2647 (.ZN(n1256), 
	.A(\UUT/Mpath/the_alu/N25 ));
   AOI22_X1 U2648 (.ZN(n1254), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N96 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N128 ));
   AOI22_X1 U2649 (.ZN(n1253), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N192 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N160 ));
   NAND2_X1 U2650 (.ZN(n5570), 
	.A2(n1258), 
	.A1(n1257));
   AOI222_X1 U2651 (.ZN(n1258), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [29]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [29]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [29]));
   AOI22_X1 U2652 (.ZN(n1257), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [29]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [29]));
   INV_X1 U2655 (.ZN(n1262), 
	.A(\UUT/Mpath/the_alu/N23 ));
   AOI22_X1 U2656 (.ZN(n1260), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N95 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N127 ));
   AOI22_X1 U2657 (.ZN(n1259), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N191 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N159 ));
   NAND2_X1 U2658 (.ZN(n5562), 
	.A2(n1264), 
	.A1(n1263));
   AOI222_X1 U2659 (.ZN(n1264), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [30]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [30]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [30]));
   AOI22_X1 U2660 (.ZN(n1263), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [30]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [30]));
   AND4_X1 U2661 (.ZN(n5526), 
	.A4(n1268), 
	.A3(n1267), 
	.A2(n1266), 
	.A1(n1265));
   NOR4_X1 U2662 (.ZN(n1268), 
	.A4(n1272), 
	.A3(n1271), 
	.A2(n1270), 
	.A1(n1269));
   NAND3_X1 U2663 (.ZN(n1272), 
	.A3(n6024), 
	.A2(n6015), 
	.A1(n6019));
   OAI211_X1 U2664 (.ZN(n1271), 
	.C2(n5412), 
	.C1(n5745), 
	.B(n6011), 
	.A(n6004));
   OAI222_X1 U2665 (.ZN(n1270), 
	.C2(n5380), 
	.C1(n5746), 
	.B2(n5252), 
	.B1(n5744), 
	.A2(n5284), 
	.A1(n5743));
   OAI221_X1 U2666 (.ZN(n1269), 
	.C2(n5220), 
	.C1(n5717), 
	.B2(n5188), 
	.B1(n5716), 
	.A(n1273));
   AOI22_X1 U2667 (.ZN(n1273), 
	.B2(n1277), 
	.B1(n1276), 
	.A2(n1275), 
	.A1(n1274));
   AOI211_X1 U2668 (.ZN(n1267), 
	.C2(n1279), 
	.C1(n1278), 
	.B(n1281), 
	.A(n1280));
   OAI22_X1 U2669 (.ZN(n1281), 
	.B2(n4740), 
	.B1(n5736), 
	.A2(n4836), 
	.A1(n5726));
   OAI222_X1 U2670 (.ZN(n1280), 
	.C2(n4708), 
	.C1(n5732), 
	.B2(n4644), 
	.B1(n5737), 
	.A2(n4676), 
	.A1(n5731));
   AOI221_X1 U2671 (.ZN(n1266), 
	.C2(n1285), 
	.C1(n1284), 
	.B2(n1283), 
	.B1(n1282), 
	.A(n1286));
   OAI22_X1 U2672 (.ZN(n1286), 
	.B2(n1288), 
	.B1(n5316), 
	.A2(n1287), 
	.A1(n4484));
   INV_X1 U2673 (.ZN(n1283), 
	.A(n5092));
   AOI222_X1 U2674 (.ZN(n1265), 
	.C2(n1294), 
	.C1(n1293), 
	.B2(n1292), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1289));
   AND4_X1 U2675 (.ZN(n5523), 
	.A4(n1298), 
	.A3(n1297), 
	.A2(n1296), 
	.A1(n1295));
   NOR4_X1 U2676 (.ZN(n1298), 
	.A4(n1302), 
	.A3(n1301), 
	.A2(n1300), 
	.A1(n1299));
   NAND3_X1 U2677 (.ZN(n1302), 
	.A3(n5993), 
	.A2(n5991), 
	.A1(n5992));
   OAI211_X1 U2678 (.ZN(n1301), 
	.C2(n5411), 
	.C1(n5745), 
	.B(n5990), 
	.A(n5989));
   OAI222_X1 U2679 (.ZN(n1300), 
	.C2(n5379), 
	.C1(n5746), 
	.B2(n5251), 
	.B1(n5744), 
	.A2(n5283), 
	.A1(n5743));
   OAI221_X1 U2680 (.ZN(n1299), 
	.C2(n5219), 
	.C1(n5717), 
	.B2(n5187), 
	.B1(n5716), 
	.A(n1303));
   AOI22_X1 U2681 (.ZN(n1303), 
	.B2(n1277), 
	.B1(n1305), 
	.A2(n1275), 
	.A1(n1304));
   AOI211_X1 U2682 (.ZN(n1297), 
	.C2(n1279), 
	.C1(n1306), 
	.B(n1308), 
	.A(n1307));
   OAI22_X1 U2683 (.ZN(n1308), 
	.B2(n4739), 
	.B1(n5736), 
	.A2(n4835), 
	.A1(n5726));
   OAI222_X1 U2684 (.ZN(n1307), 
	.C2(n4707), 
	.C1(n5732), 
	.B2(n4643), 
	.B1(n5737), 
	.A2(n4675), 
	.A1(n5731));
   AOI221_X1 U2685 (.ZN(n1296), 
	.C2(n1310), 
	.C1(n1284), 
	.B2(n1309), 
	.B1(n1282), 
	.A(n1311));
   OAI22_X1 U2686 (.ZN(n1311), 
	.B2(n1288), 
	.B1(n5315), 
	.A2(n1287), 
	.A1(n4483));
   INV_X1 U2687 (.ZN(n1309), 
	.A(n5091));
   AOI222_X1 U2688 (.ZN(n1295), 
	.C2(n1294), 
	.C1(n1314), 
	.B2(n1313), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1312));
   AND4_X1 U2689 (.ZN(n5520), 
	.A4(FE_OFN62_n1318), 
	.A3(n1317), 
	.A2(n1316), 
	.A1(n1315));
   NOR4_X1 U2690 (.ZN(n1318), 
	.A4(n1322), 
	.A3(n1321), 
	.A2(n1320), 
	.A1(n1319));
   NAND3_X1 U2691 (.ZN(n1322), 
	.A3(n5982), 
	.A2(n5980), 
	.A1(n5981));
   OAI211_X1 U2692 (.ZN(n1321), 
	.C2(n5410), 
	.C1(n5745), 
	.B(n5979), 
	.A(n5978));
   OAI222_X1 U2693 (.ZN(n1320), 
	.C2(n5378), 
	.C1(n5746), 
	.B2(n5250), 
	.B1(n5744), 
	.A2(n5282), 
	.A1(n5743));
   OAI221_X1 U2694 (.ZN(n1319), 
	.C2(n5218), 
	.C1(n5717), 
	.B2(n5186), 
	.B1(n5716), 
	.A(n1323));
   AOI22_X1 U2695 (.ZN(n1323), 
	.B2(n1277), 
	.B1(n1325), 
	.A2(n1275), 
	.A1(n1324));
   AOI211_X1 U2696 (.ZN(n1317), 
	.C2(n1279), 
	.C1(n1326), 
	.B(n1328), 
	.A(n1327));
   OAI22_X1 U2697 (.ZN(n1328), 
	.B2(n4738), 
	.B1(n5736), 
	.A2(n4834), 
	.A1(n5726));
   OAI222_X1 U2698 (.ZN(n1327), 
	.C2(n4706), 
	.C1(n5732), 
	.B2(n4642), 
	.B1(n5737), 
	.A2(n4674), 
	.A1(n5731));
   AOI221_X1 U2699 (.ZN(n1316), 
	.C2(n1330), 
	.C1(n1284), 
	.B2(n1329), 
	.B1(n1282), 
	.A(n1331));
   OAI22_X1 U2700 (.ZN(n1331), 
	.B2(n1288), 
	.B1(n5314), 
	.A2(n1287), 
	.A1(n4482));
   INV_X1 U2701 (.ZN(n1329), 
	.A(n5090));
   AOI222_X1 U2702 (.ZN(n1315), 
	.C2(n1294), 
	.C1(n1334), 
	.B2(n1333), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1332));
   AND4_X1 U2703 (.ZN(n5517), 
	.A4(FE_OFN59_n1338), 
	.A3(n1337), 
	.A2(n1336), 
	.A1(n1335));
   NOR4_X1 U2704 (.ZN(n1338), 
	.A4(n1342), 
	.A3(n1341), 
	.A2(n1340), 
	.A1(n1339));
   NAND3_X1 U2705 (.ZN(n1342), 
	.A3(n5977), 
	.A2(n5975), 
	.A1(n5976));
   OAI211_X1 U2706 (.ZN(n1341), 
	.C2(n5409), 
	.C1(n5745), 
	.B(n5974), 
	.A(n5973));
   OAI222_X1 U2707 (.ZN(n1340), 
	.C2(n5377), 
	.C1(n5746), 
	.B2(n5249), 
	.B1(n5744), 
	.A2(n5281), 
	.A1(n5743));
   OAI221_X1 U2708 (.ZN(n1339), 
	.C2(n5217), 
	.C1(n5717), 
	.B2(n5185), 
	.B1(n5716), 
	.A(n1343));
   AOI22_X1 U2709 (.ZN(n1343), 
	.B2(n1277), 
	.B1(n1345), 
	.A2(n1275), 
	.A1(n1344));
   AOI211_X1 U2710 (.ZN(n1337), 
	.C2(n1279), 
	.C1(n1346), 
	.B(n1348), 
	.A(n1347));
   OAI22_X1 U2711 (.ZN(n1348), 
	.B2(n4737), 
	.B1(n5736), 
	.A2(n4833), 
	.A1(n5726));
   OAI222_X1 U2712 (.ZN(n1347), 
	.C2(n4705), 
	.C1(n5732), 
	.B2(n4641), 
	.B1(n5737), 
	.A2(n4673), 
	.A1(n5731));
   AOI221_X1 U2713 (.ZN(n1336), 
	.C2(n1350), 
	.C1(n1284), 
	.B2(n1349), 
	.B1(n1282), 
	.A(n1351));
   OAI22_X1 U2714 (.ZN(n1351), 
	.B2(n1288), 
	.B1(n5313), 
	.A2(n1287), 
	.A1(n4481));
   INV_X1 U2715 (.ZN(n1349), 
	.A(n5089));
   AOI222_X1 U2716 (.ZN(n1335), 
	.C2(n1294), 
	.C1(n1354), 
	.B2(n1353), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1352));
   AND4_X1 U2717 (.ZN(n5514), 
	.A4(FE_OFN56_n1358), 
	.A3(n1357), 
	.A2(n1356), 
	.A1(n1355));
   NOR4_X1 U2718 (.ZN(n1358), 
	.A4(n1362), 
	.A3(n1361), 
	.A2(n1360), 
	.A1(n1359));
   NAND3_X1 U2719 (.ZN(n1362), 
	.A3(n5972), 
	.A2(n5970), 
	.A1(n5971));
   OAI211_X1 U2720 (.ZN(n1361), 
	.C2(n5408), 
	.C1(n5745), 
	.B(n5969), 
	.A(n5968));
   OAI222_X1 U2721 (.ZN(n1360), 
	.C2(n5376), 
	.C1(n5746), 
	.B2(n5248), 
	.B1(n5744), 
	.A2(n5280), 
	.A1(n5743));
   OAI221_X1 U2722 (.ZN(n1359), 
	.C2(n5216), 
	.C1(n5717), 
	.B2(n5184), 
	.B1(n5716), 
	.A(n1363));
   AOI22_X1 U2723 (.ZN(n1363), 
	.B2(n1277), 
	.B1(n1365), 
	.A2(n1275), 
	.A1(n1364));
   AOI211_X1 U2724 (.ZN(n1357), 
	.C2(n1279), 
	.C1(n1366), 
	.B(n1368), 
	.A(n1367));
   OAI22_X1 U2725 (.ZN(n1368), 
	.B2(n4736), 
	.B1(n5736), 
	.A2(n4832), 
	.A1(n5726));
   OAI222_X1 U2726 (.ZN(n1367), 
	.C2(n4704), 
	.C1(n5732), 
	.B2(n4640), 
	.B1(n5737), 
	.A2(n4672), 
	.A1(n5731));
   AOI221_X1 U2727 (.ZN(n1356), 
	.C2(n1370), 
	.C1(n1284), 
	.B2(n1369), 
	.B1(n1282), 
	.A(n1371));
   OAI22_X1 U2728 (.ZN(n1371), 
	.B2(n1288), 
	.B1(n5312), 
	.A2(n1287), 
	.A1(n4480));
   INV_X1 U2729 (.ZN(n1369), 
	.A(n5088));
   AOI222_X1 U2730 (.ZN(n1355), 
	.C2(n1294), 
	.C1(n1374), 
	.B2(n1373), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1372));
   AND4_X1 U2731 (.ZN(n5511), 
	.A4(FE_OFN53_n1378), 
	.A3(n1377), 
	.A2(n1376), 
	.A1(n1375));
   NOR4_X1 U2732 (.ZN(n1378), 
	.A4(n1382), 
	.A3(n1381), 
	.A2(n1380), 
	.A1(n1379));
   NAND3_X1 U2733 (.ZN(n1382), 
	.A3(n5967), 
	.A2(n5965), 
	.A1(n5966));
   OAI211_X1 U2734 (.ZN(n1381), 
	.C2(n5407), 
	.C1(n5745), 
	.B(n5964), 
	.A(n5963));
   OAI222_X1 U2735 (.ZN(n1380), 
	.C2(n5375), 
	.C1(n5746), 
	.B2(n5247), 
	.B1(n5744), 
	.A2(n5279), 
	.A1(n5743));
   OAI221_X1 U2736 (.ZN(n1379), 
	.C2(n5215), 
	.C1(n5717), 
	.B2(n5183), 
	.B1(n5716), 
	.A(n1383));
   AOI22_X1 U2737 (.ZN(n1383), 
	.B2(n1277), 
	.B1(n1385), 
	.A2(n1275), 
	.A1(n1384));
   AOI211_X1 U2738 (.ZN(n1377), 
	.C2(n1279), 
	.C1(n1386), 
	.B(n1388), 
	.A(n1387));
   OAI22_X1 U2739 (.ZN(n1388), 
	.B2(n4735), 
	.B1(n5736), 
	.A2(n4831), 
	.A1(n5726));
   OAI222_X1 U2740 (.ZN(n1387), 
	.C2(n4703), 
	.C1(n5732), 
	.B2(n4639), 
	.B1(n5737), 
	.A2(n4671), 
	.A1(n5731));
   AOI221_X1 U2741 (.ZN(n1376), 
	.C2(n1390), 
	.C1(n1284), 
	.B2(n1389), 
	.B1(n1282), 
	.A(n1391));
   OAI22_X1 U2742 (.ZN(n1391), 
	.B2(n1288), 
	.B1(n5311), 
	.A2(n1287), 
	.A1(n4479));
   INV_X1 U2743 (.ZN(n1389), 
	.A(n5087));
   AOI222_X1 U2744 (.ZN(n1375), 
	.C2(n1294), 
	.C1(n1394), 
	.B2(n1393), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1392));
   AND4_X1 U2745 (.ZN(n5508), 
	.A4(n1398), 
	.A3(n1397), 
	.A2(n1396), 
	.A1(n1395));
   NOR4_X1 U2746 (.ZN(n1398), 
	.A4(n1402), 
	.A3(n1401), 
	.A2(n1400), 
	.A1(n1399));
   NAND3_X1 U2747 (.ZN(n1402), 
	.A3(n5962), 
	.A2(n5960), 
	.A1(n5961));
   OAI211_X1 U2748 (.ZN(n1401), 
	.C2(n5406), 
	.C1(n5745), 
	.B(n5959), 
	.A(n5958));
   OAI222_X1 U2749 (.ZN(n1400), 
	.C2(n5374), 
	.C1(n5746), 
	.B2(n5246), 
	.B1(n5744), 
	.A2(n5278), 
	.A1(n5743));
   OAI221_X1 U2750 (.ZN(n1399), 
	.C2(n5214), 
	.C1(n5717), 
	.B2(n5182), 
	.B1(n5716), 
	.A(n1403));
   AOI22_X1 U2751 (.ZN(n1403), 
	.B2(n1277), 
	.B1(n1405), 
	.A2(n1275), 
	.A1(n1404));
   AOI211_X1 U2752 (.ZN(n1397), 
	.C2(n1279), 
	.C1(n1406), 
	.B(n1408), 
	.A(n1407));
   OAI22_X1 U2753 (.ZN(n1408), 
	.B2(n4734), 
	.B1(n5736), 
	.A2(n4830), 
	.A1(n5726));
   OAI222_X1 U2754 (.ZN(n1407), 
	.C2(n4702), 
	.C1(n5732), 
	.B2(n4638), 
	.B1(n5737), 
	.A2(n4670), 
	.A1(n5731));
   AOI221_X1 U2755 (.ZN(n1396), 
	.C2(n1410), 
	.C1(n1284), 
	.B2(n1409), 
	.B1(n1282), 
	.A(n1411));
   OAI22_X1 U2756 (.ZN(n1411), 
	.B2(n1288), 
	.B1(n5310), 
	.A2(n1287), 
	.A1(n4478));
   INV_X1 U2757 (.ZN(n1409), 
	.A(n5086));
   AOI222_X1 U2758 (.ZN(n1395), 
	.C2(n1294), 
	.C1(n1414), 
	.B2(n1413), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1412));
   AND4_X1 U2759 (.ZN(n5505), 
	.A4(FE_OFN49_n1418), 
	.A3(n1417), 
	.A2(n1416), 
	.A1(n1415));
   NOR4_X1 U2760 (.ZN(n1418), 
	.A4(n1422), 
	.A3(n1421), 
	.A2(n1420), 
	.A1(n1419));
   NAND3_X1 U2761 (.ZN(n1422), 
	.A3(n5956), 
	.A2(n5954), 
	.A1(n5955));
   OAI211_X1 U2762 (.ZN(n1421), 
	.C2(n5405), 
	.C1(n5745), 
	.B(n5953), 
	.A(n5952));
   OAI222_X1 U2763 (.ZN(n1420), 
	.C2(n5373), 
	.C1(n5746), 
	.B2(n5245), 
	.B1(n5744), 
	.A2(n5277), 
	.A1(n5743));
   OAI221_X1 U2764 (.ZN(n1419), 
	.C2(n5213), 
	.C1(n5717), 
	.B2(n5181), 
	.B1(n5716), 
	.A(n1423));
   AOI22_X1 U2765 (.ZN(n1423), 
	.B2(n1277), 
	.B1(n1425), 
	.A2(n1275), 
	.A1(n1424));
   AOI211_X1 U2766 (.ZN(n1417), 
	.C2(n1279), 
	.C1(n1426), 
	.B(n1428), 
	.A(n1427));
   OAI22_X1 U2767 (.ZN(n1428), 
	.B2(n4733), 
	.B1(n5736), 
	.A2(n4829), 
	.A1(n5726));
   OAI222_X1 U2768 (.ZN(n1427), 
	.C2(n4701), 
	.C1(n5732), 
	.B2(n4637), 
	.B1(n5737), 
	.A2(n4669), 
	.A1(n5731));
   AOI221_X1 U2769 (.ZN(n1416), 
	.C2(n1430), 
	.C1(n1284), 
	.B2(n1429), 
	.B1(n1282), 
	.A(n1431));
   OAI22_X1 U2770 (.ZN(n1431), 
	.B2(n1288), 
	.B1(n5309), 
	.A2(n1287), 
	.A1(n4477));
   INV_X1 U2771 (.ZN(n1429), 
	.A(n5085));
   AOI222_X1 U2772 (.ZN(n1415), 
	.C2(n1294), 
	.C1(n1434), 
	.B2(n1433), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1432));
   AND4_X1 U2773 (.ZN(n5502), 
	.A4(n1438), 
	.A3(n1437), 
	.A2(n1436), 
	.A1(n1435));
   NOR4_X1 U2774 (.ZN(n1438), 
	.A4(n1442), 
	.A3(n1441), 
	.A2(n1440), 
	.A1(n1439));
   NAND3_X1 U2775 (.ZN(n1442), 
	.A3(n5943), 
	.A2(n5941), 
	.A1(n5942));
   OAI211_X1 U2776 (.ZN(n1441), 
	.C2(n5404), 
	.C1(n5745), 
	.B(n5940), 
	.A(n5939));
   OAI222_X1 U2777 (.ZN(n1440), 
	.C2(n5372), 
	.C1(n5746), 
	.B2(n5244), 
	.B1(n5744), 
	.A2(n5276), 
	.A1(n5743));
   OAI221_X1 U2778 (.ZN(n1439), 
	.C2(n5212), 
	.C1(n5717), 
	.B2(n5180), 
	.B1(n5716), 
	.A(n1443));
   AOI22_X1 U2779 (.ZN(n1443), 
	.B2(n1277), 
	.B1(n1445), 
	.A2(n1275), 
	.A1(n1444));
   AOI211_X1 U2780 (.ZN(n1437), 
	.C2(n1279), 
	.C1(n1446), 
	.B(n1448), 
	.A(n1447));
   OAI22_X1 U2781 (.ZN(n1448), 
	.B2(n4732), 
	.B1(n5736), 
	.A2(n4828), 
	.A1(n5726));
   OAI222_X1 U2782 (.ZN(n1447), 
	.C2(n4700), 
	.C1(n5732), 
	.B2(n4636), 
	.B1(n5737), 
	.A2(n4668), 
	.A1(n5731));
   AOI221_X1 U2783 (.ZN(n1436), 
	.C2(n1450), 
	.C1(n1284), 
	.B2(n1449), 
	.B1(n1282), 
	.A(n1451));
   OAI22_X1 U2784 (.ZN(n1451), 
	.B2(n1288), 
	.B1(n5308), 
	.A2(n1287), 
	.A1(n4476));
   INV_X1 U2785 (.ZN(n1449), 
	.A(n5084));
   AOI222_X1 U2786 (.ZN(n1435), 
	.C2(n1294), 
	.C1(n1454), 
	.B2(n1453), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1452));
   AND4_X1 U2787 (.ZN(n5499), 
	.A4(n1458), 
	.A3(n1457), 
	.A2(n1456), 
	.A1(n1455));
   NOR4_X1 U2788 (.ZN(n1458), 
	.A4(n1462), 
	.A3(n1461), 
	.A2(n1460), 
	.A1(n1459));
   NAND3_X1 U2789 (.ZN(n1462), 
	.A3(n5938), 
	.A2(n5936), 
	.A1(n5937));
   OAI211_X1 U2790 (.ZN(n1461), 
	.C2(n5403), 
	.C1(n5745), 
	.B(n5935), 
	.A(n5934));
   OAI222_X1 U2791 (.ZN(n1460), 
	.C2(n5371), 
	.C1(n5746), 
	.B2(n5243), 
	.B1(n5744), 
	.A2(n5275), 
	.A1(n5743));
   OAI221_X1 U2792 (.ZN(n1459), 
	.C2(n5211), 
	.C1(n5717), 
	.B2(n5179), 
	.B1(n5716), 
	.A(n1463));
   AOI22_X1 U2793 (.ZN(n1463), 
	.B2(n1277), 
	.B1(n1465), 
	.A2(n1275), 
	.A1(n1464));
   AOI211_X1 U2794 (.ZN(n1457), 
	.C2(n1279), 
	.C1(n1466), 
	.B(n1468), 
	.A(n1467));
   OAI22_X1 U2795 (.ZN(n1468), 
	.B2(n4731), 
	.B1(n5736), 
	.A2(n4827), 
	.A1(n5726));
   OAI222_X1 U2796 (.ZN(n1467), 
	.C2(n4699), 
	.C1(n5732), 
	.B2(n4635), 
	.B1(n5737), 
	.A2(n4667), 
	.A1(n5731));
   AOI221_X1 U2797 (.ZN(n1456), 
	.C2(n1470), 
	.C1(n1284), 
	.B2(n1469), 
	.B1(n1282), 
	.A(n1471));
   OAI22_X1 U2798 (.ZN(n1471), 
	.B2(n1288), 
	.B1(n5307), 
	.A2(n1287), 
	.A1(n4475));
   INV_X1 U2799 (.ZN(n1469), 
	.A(n5083));
   AOI222_X1 U2800 (.ZN(n1455), 
	.C2(n1294), 
	.C1(n1474), 
	.B2(n1473), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1472));
   AND4_X1 U2801 (.ZN(n5496), 
	.A4(n1478), 
	.A3(n1477), 
	.A2(n1476), 
	.A1(n1475));
   NOR4_X1 U2802 (.ZN(n1478), 
	.A4(n1482), 
	.A3(n1481), 
	.A2(n1480), 
	.A1(n1479));
   NAND3_X1 U2803 (.ZN(n1482), 
	.A3(n5933), 
	.A2(n5931), 
	.A1(n5932));
   OAI211_X1 U2804 (.ZN(n1481), 
	.C2(n5402), 
	.C1(n5745), 
	.B(n5930), 
	.A(n5929));
   OAI222_X1 U2805 (.ZN(n1480), 
	.C2(n5370), 
	.C1(n5746), 
	.B2(n5242), 
	.B1(n5744), 
	.A2(n5274), 
	.A1(n5743));
   OAI221_X1 U2806 (.ZN(n1479), 
	.C2(n5210), 
	.C1(n5717), 
	.B2(n5178), 
	.B1(n5716), 
	.A(n1483));
   AOI22_X1 U2807 (.ZN(n1483), 
	.B2(n1277), 
	.B1(n1485), 
	.A2(n1275), 
	.A1(n1484));
   AOI211_X1 U2808 (.ZN(n1477), 
	.C2(n1279), 
	.C1(n1486), 
	.B(n1488), 
	.A(n1487));
   OAI22_X1 U2809 (.ZN(n1488), 
	.B2(n4730), 
	.B1(n5736), 
	.A2(n4826), 
	.A1(n5726));
   OAI222_X1 U2810 (.ZN(n1487), 
	.C2(n4698), 
	.C1(n5732), 
	.B2(n4634), 
	.B1(n5737), 
	.A2(n4666), 
	.A1(n5731));
   AOI221_X1 U2811 (.ZN(n1476), 
	.C2(n1490), 
	.C1(n1284), 
	.B2(n1489), 
	.B1(n1282), 
	.A(n1491));
   OAI22_X1 U2812 (.ZN(n1491), 
	.B2(n1288), 
	.B1(n5306), 
	.A2(n1287), 
	.A1(n4474));
   INV_X1 U2813 (.ZN(n1489), 
	.A(n5082));
   AOI222_X1 U2814 (.ZN(n1475), 
	.C2(n1294), 
	.C1(n1494), 
	.B2(n1493), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1492));
   AND4_X1 U2815 (.ZN(n5493), 
	.A4(FE_OFN84_n1498), 
	.A3(n1497), 
	.A2(n1496), 
	.A1(n1495));
   NOR4_X1 U2816 (.ZN(n1498), 
	.A4(n1502), 
	.A3(n1501), 
	.A2(n1500), 
	.A1(n1499));
   NAND3_X1 U2817 (.ZN(n1502), 
	.A3(n5928), 
	.A2(n5926), 
	.A1(n5927));
   OAI211_X1 U2818 (.ZN(n1501), 
	.C2(n5401), 
	.C1(n5745), 
	.B(n5925), 
	.A(n5924));
   OAI222_X1 U2819 (.ZN(n1500), 
	.C2(n5369), 
	.C1(n5746), 
	.B2(n5241), 
	.B1(n5744), 
	.A2(n5273), 
	.A1(n5743));
   OAI221_X1 U2820 (.ZN(n1499), 
	.C2(n5209), 
	.C1(n5717), 
	.B2(n5177), 
	.B1(n5716), 
	.A(n1503));
   AOI22_X1 U2821 (.ZN(n1503), 
	.B2(n1277), 
	.B1(n1505), 
	.A2(n1275), 
	.A1(n1504));
   AOI211_X1 U2822 (.ZN(n1497), 
	.C2(n1279), 
	.C1(n1506), 
	.B(n1508), 
	.A(n1507));
   OAI22_X1 U2823 (.ZN(n1508), 
	.B2(n4729), 
	.B1(n5736), 
	.A2(n4825), 
	.A1(n5726));
   OAI222_X1 U2824 (.ZN(n1507), 
	.C2(n4697), 
	.C1(n5732), 
	.B2(n4633), 
	.B1(n5737), 
	.A2(n4665), 
	.A1(n5731));
   AOI221_X1 U2825 (.ZN(n1496), 
	.C2(n1510), 
	.C1(n1284), 
	.B2(n1509), 
	.B1(n1282), 
	.A(n1511));
   OAI22_X1 U2826 (.ZN(n1511), 
	.B2(n1288), 
	.B1(n5305), 
	.A2(n1287), 
	.A1(n4473));
   INV_X1 U2827 (.ZN(n1509), 
	.A(n5081));
   AOI222_X1 U2828 (.ZN(n1495), 
	.C2(n1294), 
	.C1(n1514), 
	.B2(n1513), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1512));
   AND4_X1 U2829 (.ZN(n5490), 
	.A4(n1518), 
	.A3(n1517), 
	.A2(n1516), 
	.A1(n1515));
   NOR4_X1 U2830 (.ZN(n1518), 
	.A4(n1522), 
	.A3(n1521), 
	.A2(n1520), 
	.A1(n1519));
   NAND3_X1 U2831 (.ZN(n1522), 
	.A3(n5917), 
	.A2(n5915), 
	.A1(n5916));
   OAI211_X1 U2832 (.ZN(n1521), 
	.C2(n5400), 
	.C1(n5745), 
	.B(n5914), 
	.A(n5913));
   OAI222_X1 U2833 (.ZN(n1520), 
	.C2(n5368), 
	.C1(n5746), 
	.B2(n5240), 
	.B1(n5744), 
	.A2(n5272), 
	.A1(n5743));
   OAI221_X1 U2834 (.ZN(n1519), 
	.C2(n5208), 
	.C1(n5717), 
	.B2(n5176), 
	.B1(n5716), 
	.A(n1523));
   AOI22_X1 U2835 (.ZN(n1523), 
	.B2(n1277), 
	.B1(n1525), 
	.A2(n1275), 
	.A1(n1524));
   AOI211_X1 U2836 (.ZN(n1517), 
	.C2(n1279), 
	.C1(n1526), 
	.B(n1528), 
	.A(n1527));
   OAI22_X1 U2837 (.ZN(n1528), 
	.B2(n4728), 
	.B1(n5736), 
	.A2(n4824), 
	.A1(n5726));
   OAI222_X1 U2838 (.ZN(n1527), 
	.C2(n4696), 
	.C1(n5732), 
	.B2(n4632), 
	.B1(n5737), 
	.A2(n4664), 
	.A1(n5731));
   AOI221_X1 U2839 (.ZN(n1516), 
	.C2(n1530), 
	.C1(n1284), 
	.B2(n1529), 
	.B1(n1282), 
	.A(n1531));
   OAI22_X1 U2840 (.ZN(n1531), 
	.B2(n1288), 
	.B1(n5304), 
	.A2(n1287), 
	.A1(n4472));
   INV_X1 U2841 (.ZN(n1529), 
	.A(n5080));
   AOI222_X1 U2842 (.ZN(n1515), 
	.C2(n1294), 
	.C1(n1534), 
	.B2(n1533), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1532));
   AND4_X1 U2843 (.ZN(n5487), 
	.A4(n1538), 
	.A3(n1537), 
	.A2(n1536), 
	.A1(n1535));
   NOR4_X1 U2844 (.ZN(n1538), 
	.A4(n1542), 
	.A3(n1541), 
	.A2(n1540), 
	.A1(n1539));
   NAND3_X1 U2845 (.ZN(n1542), 
	.A3(n5912), 
	.A2(n5910), 
	.A1(n5911));
   OAI211_X1 U2846 (.ZN(n1541), 
	.C2(n5399), 
	.C1(n5745), 
	.B(n5909), 
	.A(n5908));
   OAI222_X1 U2847 (.ZN(n1540), 
	.C2(n5367), 
	.C1(n5746), 
	.B2(n5239), 
	.B1(n5744), 
	.A2(n5271), 
	.A1(n5743));
   OAI221_X1 U2848 (.ZN(n1539), 
	.C2(n5207), 
	.C1(n5717), 
	.B2(n5175), 
	.B1(n5716), 
	.A(n1543));
   AOI22_X1 U2849 (.ZN(n1543), 
	.B2(n1277), 
	.B1(n1545), 
	.A2(n1275), 
	.A1(n1544));
   AOI211_X1 U2850 (.ZN(n1537), 
	.C2(n1279), 
	.C1(n1546), 
	.B(n1548), 
	.A(n1547));
   OAI22_X1 U2851 (.ZN(n1548), 
	.B2(n4727), 
	.B1(n5736), 
	.A2(n4823), 
	.A1(n5726));
   OAI222_X1 U2852 (.ZN(n1547), 
	.C2(n4695), 
	.C1(n5732), 
	.B2(n4631), 
	.B1(n5737), 
	.A2(n4663), 
	.A1(n5731));
   AOI221_X1 U2853 (.ZN(n1536), 
	.C2(n1550), 
	.C1(n1284), 
	.B2(n1549), 
	.B1(n1282), 
	.A(n1551));
   OAI22_X1 U2854 (.ZN(n1551), 
	.B2(n1288), 
	.B1(n5303), 
	.A2(n1287), 
	.A1(n4471));
   INV_X1 U2855 (.ZN(n1549), 
	.A(n5079));
   AOI222_X1 U2856 (.ZN(n1535), 
	.C2(n1294), 
	.C1(n1554), 
	.B2(n1553), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1552));
   AND4_X1 U2857 (.ZN(n5484), 
	.A4(n1558), 
	.A3(n1557), 
	.A2(n1556), 
	.A1(n1555));
   NOR4_X1 U2858 (.ZN(n1558), 
	.A4(n1562), 
	.A3(n1561), 
	.A2(n1560), 
	.A1(n1559));
   NAND3_X1 U2859 (.ZN(n1562), 
	.A3(n5907), 
	.A2(n5905), 
	.A1(n5906));
   OAI211_X1 U2860 (.ZN(n1561), 
	.C2(n5398), 
	.C1(n5745), 
	.B(n5904), 
	.A(n5903));
   OAI222_X1 U2861 (.ZN(n1560), 
	.C2(n5366), 
	.C1(n5746), 
	.B2(n5238), 
	.B1(n5744), 
	.A2(n5270), 
	.A1(n5743));
   OAI221_X1 U2862 (.ZN(n1559), 
	.C2(n5206), 
	.C1(n5717), 
	.B2(n5174), 
	.B1(n5716), 
	.A(n1563));
   AOI22_X1 U2863 (.ZN(n1563), 
	.B2(n1277), 
	.B1(n1565), 
	.A2(n1275), 
	.A1(n1564));
   AOI211_X1 U2864 (.ZN(n1557), 
	.C2(n1279), 
	.C1(n1566), 
	.B(n1568), 
	.A(n1567));
   OAI22_X1 U2865 (.ZN(n1568), 
	.B2(n4726), 
	.B1(n5736), 
	.A2(n4822), 
	.A1(n5726));
   OAI222_X1 U2866 (.ZN(n1567), 
	.C2(n4694), 
	.C1(n5732), 
	.B2(n4630), 
	.B1(n5737), 
	.A2(n4662), 
	.A1(n5731));
   AOI221_X1 U2867 (.ZN(n1556), 
	.C2(n1570), 
	.C1(n1284), 
	.B2(n1569), 
	.B1(n1282), 
	.A(n1571));
   OAI22_X1 U2868 (.ZN(n1571), 
	.B2(n1288), 
	.B1(n5302), 
	.A2(n1287), 
	.A1(n4470));
   INV_X1 U2869 (.ZN(n1569), 
	.A(n5078));
   AOI222_X1 U2870 (.ZN(n1555), 
	.C2(n1294), 
	.C1(n1574), 
	.B2(n1573), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1572));
   AND4_X1 U2871 (.ZN(n5481), 
	.A4(n1578), 
	.A3(n1577), 
	.A2(n1576), 
	.A1(n1575));
   NOR4_X1 U2872 (.ZN(n1578), 
	.A4(n1582), 
	.A3(n1581), 
	.A2(n1580), 
	.A1(n1579));
   NAND3_X1 U2873 (.ZN(n1582), 
	.A3(n5902), 
	.A2(n5900), 
	.A1(n5901));
   OAI211_X1 U2874 (.ZN(n1581), 
	.C2(n5397), 
	.C1(n5745), 
	.B(n5899), 
	.A(n5898));
   OAI222_X1 U2875 (.ZN(n1580), 
	.C2(n5365), 
	.C1(n5746), 
	.B2(n5237), 
	.B1(n5744), 
	.A2(n5269), 
	.A1(n5743));
   OAI221_X1 U2876 (.ZN(n1579), 
	.C2(n5205), 
	.C1(n5717), 
	.B2(n5173), 
	.B1(n5716), 
	.A(n1583));
   AOI22_X1 U2877 (.ZN(n1583), 
	.B2(n1277), 
	.B1(n1585), 
	.A2(n1275), 
	.A1(n1584));
   AOI211_X1 U2878 (.ZN(n1577), 
	.C2(n1279), 
	.C1(n1586), 
	.B(n1588), 
	.A(n1587));
   OAI22_X1 U2879 (.ZN(n1588), 
	.B2(n4725), 
	.B1(n5736), 
	.A2(n4821), 
	.A1(n5726));
   OAI222_X1 U2880 (.ZN(n1587), 
	.C2(n4693), 
	.C1(n5732), 
	.B2(n4629), 
	.B1(n5737), 
	.A2(n4661), 
	.A1(n5731));
   AOI221_X1 U2881 (.ZN(n1576), 
	.C2(n1590), 
	.C1(n1284), 
	.B2(n1589), 
	.B1(n1282), 
	.A(n1591));
   OAI22_X1 U2882 (.ZN(n1591), 
	.B2(n1288), 
	.B1(n5301), 
	.A2(n1287), 
	.A1(n4469));
   INV_X1 U2883 (.ZN(n1589), 
	.A(n5077));
   AOI222_X1 U2884 (.ZN(n1575), 
	.C2(n1294), 
	.C1(n1594), 
	.B2(n1593), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1592));
   AND4_X1 U2885 (.ZN(n5478), 
	.A4(n1598), 
	.A3(n1597), 
	.A2(n1596), 
	.A1(n1595));
   NOR4_X1 U2886 (.ZN(n1598), 
	.A4(n1602), 
	.A3(n1601), 
	.A2(n1600), 
	.A1(n1599));
   NAND3_X1 U2887 (.ZN(n1602), 
	.A3(n5895), 
	.A2(n5893), 
	.A1(n5894));
   OAI211_X1 U2888 (.ZN(n1601), 
	.C2(n5396), 
	.C1(n5745), 
	.B(n5892), 
	.A(n5891));
   OAI222_X1 U2889 (.ZN(n1600), 
	.C2(n5364), 
	.C1(n5746), 
	.B2(n5236), 
	.B1(n5744), 
	.A2(n5268), 
	.A1(n5743));
   OAI221_X1 U2890 (.ZN(n1599), 
	.C2(n5204), 
	.C1(n5717), 
	.B2(n5172), 
	.B1(n5716), 
	.A(n1603));
   AOI22_X1 U2891 (.ZN(n1603), 
	.B2(n1277), 
	.B1(n1605), 
	.A2(n1275), 
	.A1(n1604));
   AOI211_X1 U2892 (.ZN(n1597), 
	.C2(n1279), 
	.C1(n1606), 
	.B(n1608), 
	.A(n1607));
   OAI22_X1 U2893 (.ZN(n1608), 
	.B2(n4724), 
	.B1(n5736), 
	.A2(n4820), 
	.A1(n5726));
   OAI222_X1 U2894 (.ZN(n1607), 
	.C2(n4692), 
	.C1(n5732), 
	.B2(n4628), 
	.B1(n5737), 
	.A2(n4660), 
	.A1(n5731));
   AOI221_X1 U2895 (.ZN(n1596), 
	.C2(n1610), 
	.C1(n1284), 
	.B2(n1609), 
	.B1(n1282), 
	.A(n1611));
   OAI22_X1 U2896 (.ZN(n1611), 
	.B2(n1288), 
	.B1(n5300), 
	.A2(n1287), 
	.A1(n4468));
   INV_X1 U2897 (.ZN(n1609), 
	.A(n5076));
   AOI222_X1 U2898 (.ZN(n1595), 
	.C2(n1294), 
	.C1(n1614), 
	.B2(n1613), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1612));
   AND4_X1 U2899 (.ZN(n5475), 
	.A4(n1618), 
	.A3(n1617), 
	.A2(n1616), 
	.A1(n1615));
   NOR4_X1 U2900 (.ZN(n1618), 
	.A4(n1622), 
	.A3(n1621), 
	.A2(n1620), 
	.A1(n1619));
   NAND3_X1 U2901 (.ZN(n1622), 
	.A3(n5887), 
	.A2(n5885), 
	.A1(n5886));
   OAI211_X1 U2902 (.ZN(n1621), 
	.C2(n5395), 
	.C1(n5745), 
	.B(n5884), 
	.A(n5883));
   OAI222_X1 U2903 (.ZN(n1620), 
	.C2(n5363), 
	.C1(n5746), 
	.B2(n5235), 
	.B1(n5744), 
	.A2(n5267), 
	.A1(n5743));
   OAI221_X1 U2904 (.ZN(n1619), 
	.C2(n5203), 
	.C1(n5717), 
	.B2(n5171), 
	.B1(n5716), 
	.A(n1623));
   AOI22_X1 U2905 (.ZN(n1623), 
	.B2(n1277), 
	.B1(n1625), 
	.A2(n1275), 
	.A1(n1624));
   AOI211_X1 U2906 (.ZN(n1617), 
	.C2(n1279), 
	.C1(n1626), 
	.B(n1628), 
	.A(n1627));
   OAI22_X1 U2907 (.ZN(n1628), 
	.B2(n4723), 
	.B1(n5736), 
	.A2(n4819), 
	.A1(n5726));
   OAI222_X1 U2908 (.ZN(n1627), 
	.C2(n4691), 
	.C1(n5732), 
	.B2(n4627), 
	.B1(n5737), 
	.A2(n4659), 
	.A1(n5731));
   AOI221_X1 U2909 (.ZN(n1616), 
	.C2(n1630), 
	.C1(n1284), 
	.B2(n1629), 
	.B1(n1282), 
	.A(n1631));
   OAI22_X1 U2910 (.ZN(n1631), 
	.B2(n1288), 
	.B1(n5299), 
	.A2(n1287), 
	.A1(n4467));
   INV_X1 U2911 (.ZN(n1629), 
	.A(n5075));
   AOI222_X1 U2912 (.ZN(n1615), 
	.C2(n1294), 
	.C1(n1634), 
	.B2(n1633), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1632));
   AND4_X1 U2913 (.ZN(n5472), 
	.A4(n1638), 
	.A3(n1637), 
	.A2(n1636), 
	.A1(n1635));
   NOR4_X1 U2914 (.ZN(n1638), 
	.A4(n1642), 
	.A3(n1641), 
	.A2(n1640), 
	.A1(n1639));
   NAND3_X1 U2915 (.ZN(n1642), 
	.A3(n5878), 
	.A2(n5876), 
	.A1(n5877));
   OAI211_X1 U2916 (.ZN(n1641), 
	.C2(n5394), 
	.C1(n5745), 
	.B(n5875), 
	.A(n5874));
   OAI222_X1 U2917 (.ZN(n1640), 
	.C2(n5362), 
	.C1(n5746), 
	.B2(n5234), 
	.B1(n5744), 
	.A2(n5266), 
	.A1(n5743));
   OAI221_X1 U2918 (.ZN(n1639), 
	.C2(n5202), 
	.C1(n5717), 
	.B2(n5170), 
	.B1(n5716), 
	.A(n1643));
   AOI22_X1 U2919 (.ZN(n1643), 
	.B2(n1277), 
	.B1(n1645), 
	.A2(n1275), 
	.A1(n1644));
   AOI211_X1 U2920 (.ZN(n1637), 
	.C2(n1279), 
	.C1(n1646), 
	.B(n1648), 
	.A(n1647));
   OAI22_X1 U2921 (.ZN(n1648), 
	.B2(n4722), 
	.B1(n5736), 
	.A2(n4818), 
	.A1(n5726));
   OAI222_X1 U2922 (.ZN(n1647), 
	.C2(n4690), 
	.C1(n5732), 
	.B2(n4626), 
	.B1(n5737), 
	.A2(n4658), 
	.A1(n5731));
   AOI221_X1 U2923 (.ZN(n1636), 
	.C2(n1650), 
	.C1(n1284), 
	.B2(n1649), 
	.B1(n1282), 
	.A(n1651));
   OAI22_X1 U2924 (.ZN(n1651), 
	.B2(n1288), 
	.B1(n5298), 
	.A2(n1287), 
	.A1(n4466));
   INV_X1 U2925 (.ZN(n1649), 
	.A(n5074));
   AOI222_X1 U2926 (.ZN(n1635), 
	.C2(n1294), 
	.C1(n1654), 
	.B2(n1653), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1652));
   AND4_X1 U2927 (.ZN(n5469), 
	.A4(n1658), 
	.A3(n1657), 
	.A2(n1656), 
	.A1(n1655));
   NOR4_X1 U2928 (.ZN(n1658), 
	.A4(n1662), 
	.A3(n1661), 
	.A2(n1660), 
	.A1(n1659));
   NAND3_X1 U2929 (.ZN(n1662), 
	.A3(n5868), 
	.A2(n5866), 
	.A1(n5867));
   OAI211_X1 U2930 (.ZN(n1661), 
	.C2(n5393), 
	.C1(n5745), 
	.B(n5865), 
	.A(n5864));
   OAI222_X1 U2931 (.ZN(n1660), 
	.C2(n5361), 
	.C1(n5746), 
	.B2(n5233), 
	.B1(n5744), 
	.A2(n5265), 
	.A1(n5743));
   OAI221_X1 U2932 (.ZN(n1659), 
	.C2(n5201), 
	.C1(n5717), 
	.B2(n5169), 
	.B1(n5716), 
	.A(n1663));
   AOI22_X1 U2933 (.ZN(n1663), 
	.B2(n1277), 
	.B1(n1665), 
	.A2(n1275), 
	.A1(n1664));
   AOI211_X1 U2934 (.ZN(n1657), 
	.C2(n1279), 
	.C1(n1666), 
	.B(n1668), 
	.A(n1667));
   OAI22_X1 U2935 (.ZN(n1668), 
	.B2(n4721), 
	.B1(n5736), 
	.A2(n4817), 
	.A1(n5726));
   OAI222_X1 U2936 (.ZN(n1667), 
	.C2(n4689), 
	.C1(n5732), 
	.B2(n4625), 
	.B1(n5737), 
	.A2(n4657), 
	.A1(n5731));
   AOI221_X1 U2937 (.ZN(n1656), 
	.C2(n1670), 
	.C1(n1284), 
	.B2(n1669), 
	.B1(n1282), 
	.A(n1671));
   OAI22_X1 U2938 (.ZN(n1671), 
	.B2(n1288), 
	.B1(n5297), 
	.A2(n1287), 
	.A1(n4465));
   INV_X1 U2939 (.ZN(n1669), 
	.A(n5073));
   AOI222_X1 U2940 (.ZN(n1655), 
	.C2(n1294), 
	.C1(n1674), 
	.B2(n1673), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1672));
   AND4_X1 U2941 (.ZN(n5466), 
	.A4(n1678), 
	.A3(n1677), 
	.A2(n1676), 
	.A1(n1675));
   NOR4_X1 U2942 (.ZN(n1678), 
	.A4(n1682), 
	.A3(n1681), 
	.A2(n1680), 
	.A1(n1679));
   NAND3_X1 U2943 (.ZN(n1682), 
	.A3(n5862), 
	.A2(n5860), 
	.A1(n5861));
   OAI211_X1 U2944 (.ZN(n1681), 
	.C2(n5392), 
	.C1(n5745), 
	.B(n5859), 
	.A(n5858));
   OAI222_X1 U2945 (.ZN(n1680), 
	.C2(n5360), 
	.C1(n5746), 
	.B2(n5232), 
	.B1(n5744), 
	.A2(n5264), 
	.A1(n5743));
   OAI221_X1 U2946 (.ZN(n1679), 
	.C2(n5200), 
	.C1(n5717), 
	.B2(n5168), 
	.B1(n5716), 
	.A(n1683));
   AOI22_X1 U2947 (.ZN(n1683), 
	.B2(n1277), 
	.B1(n1685), 
	.A2(n1275), 
	.A1(n1684));
   AOI211_X1 U2948 (.ZN(n1677), 
	.C2(n1279), 
	.C1(n1686), 
	.B(n1688), 
	.A(n1687));
   OAI22_X1 U2949 (.ZN(n1688), 
	.B2(n4720), 
	.B1(n5736), 
	.A2(n4816), 
	.A1(n5726));
   OAI222_X1 U2950 (.ZN(n1687), 
	.C2(n4688), 
	.C1(n5732), 
	.B2(n4624), 
	.B1(n5737), 
	.A2(n4656), 
	.A1(n5731));
   AOI221_X1 U2951 (.ZN(n1676), 
	.C2(n1690), 
	.C1(n1284), 
	.B2(n1689), 
	.B1(n1282), 
	.A(n1691));
   OAI22_X1 U2952 (.ZN(n1691), 
	.B2(n1288), 
	.B1(n5296), 
	.A2(n1287), 
	.A1(n4464));
   INV_X1 U2953 (.ZN(n1689), 
	.A(n5072));
   AOI222_X1 U2954 (.ZN(n1675), 
	.C2(n1294), 
	.C1(n1694), 
	.B2(n1693), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1692));
   AND4_X1 U2955 (.ZN(n5463), 
	.A4(n1698), 
	.A3(n1697), 
	.A2(n1696), 
	.A1(n1695));
   NOR4_X1 U2956 (.ZN(n1698), 
	.A4(n1702), 
	.A3(n1701), 
	.A2(n1700), 
	.A1(n1699));
   NAND3_X1 U2957 (.ZN(n1702), 
	.A3(n5856), 
	.A2(n5854), 
	.A1(n5855));
   OAI211_X1 U2958 (.ZN(n1701), 
	.C2(n5391), 
	.C1(n5745), 
	.B(n5853), 
	.A(n5852));
   OAI222_X1 U2959 (.ZN(n1700), 
	.C2(n5359), 
	.C1(n5746), 
	.B2(n5231), 
	.B1(n5744), 
	.A2(n5263), 
	.A1(n5743));
   OAI221_X1 U2960 (.ZN(n1699), 
	.C2(n5199), 
	.C1(n5717), 
	.B2(n5167), 
	.B1(n5716), 
	.A(n1703));
   AOI22_X1 U2961 (.ZN(n1703), 
	.B2(n1277), 
	.B1(n1705), 
	.A2(n1275), 
	.A1(n1704));
   AOI211_X1 U2962 (.ZN(n1697), 
	.C2(n1279), 
	.C1(n1706), 
	.B(n1708), 
	.A(n1707));
   OAI22_X1 U2963 (.ZN(n1708), 
	.B2(n4719), 
	.B1(n5736), 
	.A2(n4815), 
	.A1(n5726));
   OAI222_X1 U2964 (.ZN(n1707), 
	.C2(n4687), 
	.C1(n5732), 
	.B2(n4623), 
	.B1(n5737), 
	.A2(n4655), 
	.A1(n5731));
   AOI221_X1 U2965 (.ZN(n1696), 
	.C2(n1710), 
	.C1(n1284), 
	.B2(n1709), 
	.B1(n1282), 
	.A(n1711));
   OAI22_X1 U2966 (.ZN(n1711), 
	.B2(n1288), 
	.B1(n5295), 
	.A2(n1287), 
	.A1(n4463));
   INV_X1 U2967 (.ZN(n1709), 
	.A(n5071));
   AOI222_X1 U2968 (.ZN(n1695), 
	.C2(n1294), 
	.C1(n1714), 
	.B2(n1713), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1712));
   AND4_X1 U2969 (.ZN(n5460), 
	.A4(FE_OFN82_n1718), 
	.A3(n1717), 
	.A2(n1716), 
	.A1(n1715));
   NOR4_X1 U2970 (.ZN(n1718), 
	.A4(n1722), 
	.A3(n1721), 
	.A2(n1720), 
	.A1(n1719));
   NAND3_X1 U2971 (.ZN(n1722), 
	.A3(n5850), 
	.A2(n5848), 
	.A1(n5849));
   OAI211_X1 U2972 (.ZN(n1721), 
	.C2(n5390), 
	.C1(n5745), 
	.B(n5847), 
	.A(n5846));
   OAI222_X1 U2973 (.ZN(n1720), 
	.C2(n5358), 
	.C1(n5746), 
	.B2(n5230), 
	.B1(n5744), 
	.A2(n5262), 
	.A1(n5743));
   OAI221_X1 U2974 (.ZN(n1719), 
	.C2(n5198), 
	.C1(n5717), 
	.B2(n5166), 
	.B1(n5716), 
	.A(n1723));
   AOI22_X1 U2975 (.ZN(n1723), 
	.B2(n1277), 
	.B1(n1725), 
	.A2(n1275), 
	.A1(n1724));
   AOI211_X1 U2976 (.ZN(n1717), 
	.C2(n1279), 
	.C1(n1726), 
	.B(n1728), 
	.A(n1727));
   OAI22_X1 U2977 (.ZN(n1728), 
	.B2(n4718), 
	.B1(n5736), 
	.A2(n4814), 
	.A1(n5726));
   OAI222_X1 U2978 (.ZN(n1727), 
	.C2(n4686), 
	.C1(n5732), 
	.B2(n4622), 
	.B1(n5737), 
	.A2(n4654), 
	.A1(n5731));
   AOI221_X1 U2979 (.ZN(n1716), 
	.C2(n1730), 
	.C1(n1284), 
	.B2(n1729), 
	.B1(n1282), 
	.A(n1731));
   OAI22_X1 U2980 (.ZN(n1731), 
	.B2(n1288), 
	.B1(n5294), 
	.A2(n1287), 
	.A1(n4462));
   INV_X1 U2981 (.ZN(n1729), 
	.A(n5070));
   AOI222_X1 U2982 (.ZN(n1715), 
	.C2(n1294), 
	.C1(n1734), 
	.B2(n1733), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1732));
   AND4_X1 U2983 (.ZN(n5457), 
	.A4(n1738), 
	.A3(n1737), 
	.A2(n1736), 
	.A1(n1735));
   NOR4_X1 U2984 (.ZN(n1738), 
	.A4(n1742), 
	.A3(n1741), 
	.A2(n1740), 
	.A1(n1739));
   NAND3_X1 U2985 (.ZN(n1742), 
	.A3(n5837), 
	.A2(n5835), 
	.A1(n5836));
   OAI211_X1 U2986 (.ZN(n1741), 
	.C2(n5389), 
	.C1(n5745), 
	.B(n5834), 
	.A(n5833));
   OAI222_X1 U2987 (.ZN(n1740), 
	.C2(n5357), 
	.C1(n5746), 
	.B2(n5229), 
	.B1(n5744), 
	.A2(n5261), 
	.A1(n5743));
   OAI221_X1 U2988 (.ZN(n1739), 
	.C2(n5197), 
	.C1(n5717), 
	.B2(n5165), 
	.B1(n5716), 
	.A(n1743));
   AOI22_X1 U2989 (.ZN(n1743), 
	.B2(n1277), 
	.B1(n1745), 
	.A2(n1275), 
	.A1(n1744));
   AOI211_X1 U2990 (.ZN(n1737), 
	.C2(n1279), 
	.C1(n1746), 
	.B(n1748), 
	.A(n1747));
   OAI22_X1 U2991 (.ZN(n1748), 
	.B2(n4717), 
	.B1(n5736), 
	.A2(n4813), 
	.A1(n5726));
   OAI222_X1 U2992 (.ZN(n1747), 
	.C2(n4685), 
	.C1(n5732), 
	.B2(n4621), 
	.B1(n5737), 
	.A2(n4653), 
	.A1(n5731));
   AOI221_X1 U2993 (.ZN(n1736), 
	.C2(n1750), 
	.C1(n1284), 
	.B2(n1749), 
	.B1(n1282), 
	.A(n1751));
   OAI22_X1 U2994 (.ZN(n1751), 
	.B2(n1288), 
	.B1(n5293), 
	.A2(n1287), 
	.A1(n4461));
   INV_X1 U2995 (.ZN(n1749), 
	.A(n5069));
   AOI222_X1 U2996 (.ZN(n1735), 
	.C2(n1294), 
	.C1(n1754), 
	.B2(n1753), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1752));
   AND4_X1 U2997 (.ZN(n5454), 
	.A4(n1758), 
	.A3(n1757), 
	.A2(n1756), 
	.A1(n1755));
   NOR4_X1 U2998 (.ZN(n1758), 
	.A4(n1762), 
	.A3(n1761), 
	.A2(n1760), 
	.A1(n1759));
   NAND3_X1 U2999 (.ZN(n1762), 
	.A3(n5830), 
	.A2(n5828), 
	.A1(n5829));
   OAI211_X1 U3000 (.ZN(n1761), 
	.C2(n5388), 
	.C1(n5745), 
	.B(n5827), 
	.A(n5826));
   OAI222_X1 U3001 (.ZN(n1760), 
	.C2(n5356), 
	.C1(n5746), 
	.B2(n5228), 
	.B1(n5744), 
	.A2(n5260), 
	.A1(n5743));
   OAI221_X1 U3002 (.ZN(n1759), 
	.C2(n5196), 
	.C1(n5717), 
	.B2(n5164), 
	.B1(n5716), 
	.A(n1763));
   AOI22_X1 U3003 (.ZN(n1763), 
	.B2(n1277), 
	.B1(n1765), 
	.A2(n1275), 
	.A1(n1764));
   AOI211_X1 U3004 (.ZN(n1757), 
	.C2(n1279), 
	.C1(n1766), 
	.B(n1768), 
	.A(n1767));
   OAI22_X1 U3005 (.ZN(n1768), 
	.B2(n4716), 
	.B1(n5736), 
	.A2(n4812), 
	.A1(n5726));
   OAI222_X1 U3006 (.ZN(n1767), 
	.C2(n4684), 
	.C1(n5732), 
	.B2(n4620), 
	.B1(n5737), 
	.A2(n4652), 
	.A1(n5731));
   AOI221_X1 U3007 (.ZN(n1756), 
	.C2(n1770), 
	.C1(n1284), 
	.B2(n1769), 
	.B1(n1282), 
	.A(n1771));
   OAI22_X1 U3008 (.ZN(n1771), 
	.B2(n1288), 
	.B1(n5292), 
	.A2(n1287), 
	.A1(n4460));
   INV_X1 U3009 (.ZN(n1769), 
	.A(n5068));
   AOI222_X1 U3010 (.ZN(n1755), 
	.C2(n1294), 
	.C1(n1774), 
	.B2(n1773), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1772));
   AND4_X1 U3011 (.ZN(n5451), 
	.A4(FE_OFN79_n1778), 
	.A3(n1777), 
	.A2(n1776), 
	.A1(n1775));
   NOR4_X1 U3012 (.ZN(n1778), 
	.A4(n1782), 
	.A3(n1781), 
	.A2(n1780), 
	.A1(n1779));
   NAND3_X1 U3013 (.ZN(n1782), 
	.A3(n5824), 
	.A2(n5822), 
	.A1(n5823));
   OAI211_X1 U3014 (.ZN(n1781), 
	.C2(n5387), 
	.C1(n5745), 
	.B(n5821), 
	.A(n5820));
   OAI222_X1 U3015 (.ZN(n1780), 
	.C2(n5355), 
	.C1(n5746), 
	.B2(n5227), 
	.B1(n5744), 
	.A2(n5259), 
	.A1(n5743));
   OAI221_X1 U3016 (.ZN(n1779), 
	.C2(n5195), 
	.C1(n5717), 
	.B2(n5163), 
	.B1(n5716), 
	.A(n1783));
   AOI22_X1 U3017 (.ZN(n1783), 
	.B2(n1277), 
	.B1(n1785), 
	.A2(n1275), 
	.A1(n1784));
   AOI211_X1 U3018 (.ZN(n1777), 
	.C2(n1279), 
	.C1(n1786), 
	.B(n1788), 
	.A(n1787));
   OAI22_X1 U3019 (.ZN(n1788), 
	.B2(n4715), 
	.B1(n5736), 
	.A2(n4811), 
	.A1(n5726));
   OAI222_X1 U3020 (.ZN(n1787), 
	.C2(n4683), 
	.C1(n5732), 
	.B2(n4619), 
	.B1(n5737), 
	.A2(n4651), 
	.A1(n5731));
   AOI221_X1 U3021 (.ZN(n1776), 
	.C2(n1790), 
	.C1(n1284), 
	.B2(n1789), 
	.B1(n1282), 
	.A(n1791));
   OAI22_X1 U3022 (.ZN(n1791), 
	.B2(n1288), 
	.B1(n5291), 
	.A2(n1287), 
	.A1(n4459));
   INV_X1 U3023 (.ZN(n1789), 
	.A(n5067));
   AOI222_X1 U3024 (.ZN(n1775), 
	.C2(n1294), 
	.C1(n1794), 
	.B2(n1793), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1792));
   AND4_X1 U3025 (.ZN(n5448), 
	.A4(FE_OFN76_n1798), 
	.A3(n1797), 
	.A2(n1796), 
	.A1(n1795));
   NOR4_X1 U3026 (.ZN(n1798), 
	.A4(n1802), 
	.A3(n1801), 
	.A2(n1800), 
	.A1(n1799));
   NAND3_X1 U3027 (.ZN(n1802), 
	.A3(n5811), 
	.A2(n5809), 
	.A1(n5810));
   OAI211_X1 U3028 (.ZN(n1801), 
	.C2(n5386), 
	.C1(n5745), 
	.B(n5808), 
	.A(n5807));
   OAI222_X1 U3029 (.ZN(n1800), 
	.C2(n5354), 
	.C1(n5746), 
	.B2(n5226), 
	.B1(n5744), 
	.A2(n5258), 
	.A1(n5743));
   OAI221_X1 U3030 (.ZN(n1799), 
	.C2(n5194), 
	.C1(n5717), 
	.B2(n5162), 
	.B1(n5716), 
	.A(n1803));
   AOI22_X1 U3031 (.ZN(n1803), 
	.B2(n1277), 
	.B1(n1805), 
	.A2(n1275), 
	.A1(n1804));
   AOI211_X1 U3032 (.ZN(n1797), 
	.C2(n1279), 
	.C1(n1806), 
	.B(n1808), 
	.A(n1807));
   OAI22_X1 U3033 (.ZN(n1808), 
	.B2(n4714), 
	.B1(n5736), 
	.A2(n4810), 
	.A1(n5726));
   OAI222_X1 U3034 (.ZN(n1807), 
	.C2(n4682), 
	.C1(n5732), 
	.B2(n4618), 
	.B1(n5737), 
	.A2(n4650), 
	.A1(n5731));
   AOI221_X1 U3035 (.ZN(n1796), 
	.C2(n1810), 
	.C1(n1284), 
	.B2(n1809), 
	.B1(n1282), 
	.A(n1811));
   OAI22_X1 U3036 (.ZN(n1811), 
	.B2(n1288), 
	.B1(n5290), 
	.A2(n1287), 
	.A1(n4458));
   INV_X1 U3037 (.ZN(n1809), 
	.A(n5066));
   AOI222_X1 U3038 (.ZN(n1795), 
	.C2(n1294), 
	.C1(n1814), 
	.B2(n1813), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1812));
   AND4_X1 U3039 (.ZN(n5445), 
	.A4(FE_OFN73_n1818), 
	.A3(n1817), 
	.A2(n1816), 
	.A1(n1815));
   NOR4_X1 U3040 (.ZN(n1818), 
	.A4(n1822), 
	.A3(n1821), 
	.A2(n1820), 
	.A1(n1819));
   NAND3_X1 U3041 (.ZN(n1822), 
	.A3(n5798), 
	.A2(n5796), 
	.A1(n5797));
   OAI211_X1 U3042 (.ZN(n1821), 
	.C2(n5385), 
	.C1(n5745), 
	.B(n5795), 
	.A(n5794));
   OAI222_X1 U3043 (.ZN(n1820), 
	.C2(n5353), 
	.C1(n5746), 
	.B2(n5225), 
	.B1(n5744), 
	.A2(n5257), 
	.A1(n5743));
   OAI221_X1 U3044 (.ZN(n1819), 
	.C2(n5193), 
	.C1(n5717), 
	.B2(n5161), 
	.B1(n5716), 
	.A(n1823));
   AOI22_X1 U3045 (.ZN(n1823), 
	.B2(n1277), 
	.B1(n1825), 
	.A2(n1275), 
	.A1(n1824));
   AOI211_X1 U3046 (.ZN(n1817), 
	.C2(n1279), 
	.C1(n1826), 
	.B(n1828), 
	.A(n1827));
   OAI22_X1 U3047 (.ZN(n1828), 
	.B2(n4713), 
	.B1(n5736), 
	.A2(n4809), 
	.A1(n5726));
   OAI222_X1 U3048 (.ZN(n1827), 
	.C2(n4681), 
	.C1(n5732), 
	.B2(n4617), 
	.B1(n5737), 
	.A2(n4649), 
	.A1(n5731));
   AOI221_X1 U3049 (.ZN(n1816), 
	.C2(n1830), 
	.C1(n1284), 
	.B2(n1829), 
	.B1(n1282), 
	.A(n1831));
   OAI22_X1 U3050 (.ZN(n1831), 
	.B2(n1288), 
	.B1(n5289), 
	.A2(n1287), 
	.A1(n4457));
   INV_X1 U3051 (.ZN(n1829), 
	.A(n5065));
   AOI222_X1 U3052 (.ZN(n1815), 
	.C2(n1294), 
	.C1(n1834), 
	.B2(n1833), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1832));
   AND4_X1 U3053 (.ZN(n5442), 
	.A4(n1838), 
	.A3(n1837), 
	.A2(n1836), 
	.A1(n1835));
   NOR4_X1 U3054 (.ZN(n1838), 
	.A4(n1842), 
	.A3(n1841), 
	.A2(n1840), 
	.A1(n1839));
   NAND3_X1 U3055 (.ZN(n1842), 
	.A3(n5785), 
	.A2(n5783), 
	.A1(n5784));
   OAI211_X1 U3056 (.ZN(n1841), 
	.C2(n5384), 
	.C1(n5745), 
	.B(n5782), 
	.A(n5781));
   OAI222_X1 U3057 (.ZN(n1840), 
	.C2(n5352), 
	.C1(n5746), 
	.B2(n5224), 
	.B1(n5744), 
	.A2(n5256), 
	.A1(n5743));
   OAI221_X1 U3058 (.ZN(n1839), 
	.C2(n5192), 
	.C1(n5717), 
	.B2(n5160), 
	.B1(n5716), 
	.A(n1843));
   AOI22_X1 U3059 (.ZN(n1843), 
	.B2(n1277), 
	.B1(n1845), 
	.A2(n1275), 
	.A1(n1844));
   AOI211_X1 U3060 (.ZN(n1837), 
	.C2(n1279), 
	.C1(n1846), 
	.B(n1848), 
	.A(n1847));
   OAI22_X1 U3061 (.ZN(n1848), 
	.B2(n4712), 
	.B1(n5736), 
	.A2(n4808), 
	.A1(n5726));
   OAI222_X1 U3062 (.ZN(n1847), 
	.C2(n4680), 
	.C1(n5732), 
	.B2(n4616), 
	.B1(n5737), 
	.A2(n4648), 
	.A1(n5731));
   AOI221_X1 U3063 (.ZN(n1836), 
	.C2(n1850), 
	.C1(n1284), 
	.B2(n1849), 
	.B1(n1282), 
	.A(n1851));
   OAI22_X1 U3064 (.ZN(n1851), 
	.B2(n1288), 
	.B1(n5288), 
	.A2(n1287), 
	.A1(n4456));
   INV_X1 U3065 (.ZN(n1849), 
	.A(n5064));
   AOI222_X1 U3066 (.ZN(n1835), 
	.C2(n1294), 
	.C1(n1854), 
	.B2(n1853), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1852));
   AND4_X1 U3067 (.ZN(n5439), 
	.A4(FE_OFN68_n1858), 
	.A3(n1857), 
	.A2(n1856), 
	.A1(n1855));
   NOR4_X1 U3068 (.ZN(n1858), 
	.A4(n1862), 
	.A3(n1861), 
	.A2(n1860), 
	.A1(n1859));
   NAND3_X1 U3069 (.ZN(n1862), 
	.A3(n5768), 
	.A2(n5766), 
	.A1(n5767));
   OAI211_X1 U3070 (.ZN(n1861), 
	.C2(n5383), 
	.C1(n5745), 
	.B(n5765), 
	.A(n5764));
   OAI222_X1 U3071 (.ZN(n1860), 
	.C2(n5351), 
	.C1(n5746), 
	.B2(n5223), 
	.B1(n5744), 
	.A2(n5255), 
	.A1(n5743));
   OAI221_X1 U3072 (.ZN(n1859), 
	.C2(n5191), 
	.C1(n5717), 
	.B2(n5159), 
	.B1(n5716), 
	.A(n1863));
   AOI22_X1 U3073 (.ZN(n1863), 
	.B2(n1277), 
	.B1(n1865), 
	.A2(n1275), 
	.A1(n1864));
   AOI211_X1 U3074 (.ZN(n1857), 
	.C2(n1279), 
	.C1(n1866), 
	.B(n1868), 
	.A(n1867));
   OAI22_X1 U3075 (.ZN(n1868), 
	.B2(n4711), 
	.B1(n5736), 
	.A2(n4807), 
	.A1(n5726));
   OAI222_X1 U3076 (.ZN(n1867), 
	.C2(n4679), 
	.C1(n5732), 
	.B2(n4615), 
	.B1(n5737), 
	.A2(n4647), 
	.A1(n5731));
   AOI221_X1 U3077 (.ZN(n1856), 
	.C2(n1870), 
	.C1(n1284), 
	.B2(n1869), 
	.B1(n1282), 
	.A(n1871));
   OAI22_X1 U3078 (.ZN(n1871), 
	.B2(n1288), 
	.B1(n5287), 
	.A2(n1287), 
	.A1(n4455));
   INV_X1 U3079 (.ZN(n1869), 
	.A(n5063));
   AOI222_X1 U3080 (.ZN(n1855), 
	.C2(n1294), 
	.C1(n1874), 
	.B2(n1873), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1872));
   AND4_X1 U3081 (.ZN(n5436), 
	.A4(FE_OFN93_n1878), 
	.A3(n1877), 
	.A2(n1876), 
	.A1(n1875));
   NOR4_X1 U3082 (.ZN(n1878), 
	.A4(n1882), 
	.A3(n1881), 
	.A2(n1880), 
	.A1(n1879));
   NAND3_X1 U3083 (.ZN(n1882), 
	.A3(n5753), 
	.A2(n5751), 
	.A1(n5752));
   OAI211_X1 U3084 (.ZN(n1881), 
	.C2(n5382), 
	.C1(n5745), 
	.B(n5750), 
	.A(n5749));
   OAI222_X1 U3085 (.ZN(n1880), 
	.C2(n5350), 
	.C1(n5746), 
	.B2(n5222), 
	.B1(n5744), 
	.A2(n5254), 
	.A1(n5743));
   OAI221_X1 U3086 (.ZN(n1879), 
	.C2(n5190), 
	.C1(n5717), 
	.B2(n5158), 
	.B1(n5716), 
	.A(n1883));
   AOI22_X1 U3087 (.ZN(n1883), 
	.B2(n1277), 
	.B1(n1885), 
	.A2(n1275), 
	.A1(n1884));
   AOI211_X1 U3088 (.ZN(n1877), 
	.C2(n1279), 
	.C1(n1886), 
	.B(n1888), 
	.A(n1887));
   OAI22_X1 U3089 (.ZN(n1888), 
	.B2(n4710), 
	.B1(n5736), 
	.A2(n4806), 
	.A1(n5726));
   OAI222_X1 U3090 (.ZN(n1887), 
	.C2(n4678), 
	.C1(n5732), 
	.B2(n4614), 
	.B1(n5737), 
	.A2(n4646), 
	.A1(n5731));
   AOI221_X1 U3091 (.ZN(n1876), 
	.C2(n1890), 
	.C1(n1284), 
	.B2(n1889), 
	.B1(n1282), 
	.A(n1891));
   OAI22_X1 U3092 (.ZN(n1891), 
	.B2(n1288), 
	.B1(n5286), 
	.A2(n1287), 
	.A1(n4454));
   INV_X1 U3093 (.ZN(n1889), 
	.A(n5062));
   AOI222_X1 U3094 (.ZN(n1875), 
	.C2(n1294), 
	.C1(n1894), 
	.B2(n1893), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1892));
   AND4_X1 U3095 (.ZN(n5431), 
	.A4(n1898), 
	.A3(n1897), 
	.A2(n1896), 
	.A1(n1895));
   NOR4_X1 U3096 (.ZN(n1898), 
	.A4(n1902), 
	.A3(n1901), 
	.A2(n1900), 
	.A1(n1899));
   NAND3_X1 U3097 (.ZN(n1902), 
	.A3(n5740), 
	.A2(n5728), 
	.A1(n5733));
   OAI211_X1 U3098 (.ZN(n1901), 
	.C2(n5381), 
	.C1(n5745), 
	.B(n5723), 
	.A(n5718));
   OAI222_X1 U3099 (.ZN(n1900), 
	.C2(n5349), 
	.C1(n5746), 
	.B2(n5221), 
	.B1(n5744), 
	.A2(n5253), 
	.A1(n5743));
   OAI221_X1 U3100 (.ZN(n1899), 
	.C2(n5189), 
	.C1(n5717), 
	.B2(n5157), 
	.B1(n5716), 
	.A(n1903));
   AOI22_X1 U3101 (.ZN(n1903), 
	.B2(n1277), 
	.B1(n1905), 
	.A2(n1275), 
	.A1(n1904));
   AOI211_X1 U3104 (.ZN(n1897), 
	.C2(n1279), 
	.C1(n1906), 
	.B(n1908), 
	.A(n1907));
   OAI22_X1 U3105 (.ZN(n1908), 
	.B2(n4709), 
	.B1(n5736), 
	.A2(n4805), 
	.A1(n5726));
   OAI222_X1 U3106 (.ZN(n1907), 
	.C2(n4677), 
	.C1(n5732), 
	.B2(n4613), 
	.B1(n5737), 
	.A2(n4645), 
	.A1(n5731));
   AOI221_X1 U3108 (.ZN(n1896), 
	.C2(n1910), 
	.C1(n1284), 
	.B2(n1909), 
	.B1(n1282), 
	.A(n1911));
   OAI22_X1 U3109 (.ZN(n1911), 
	.B2(n1288), 
	.B1(n5285), 
	.A2(n1287), 
	.A1(n4453));
   INV_X1 U3114 (.ZN(n1909), 
	.A(n5061));
   AOI222_X1 U3116 (.ZN(n1895), 
	.C2(n1294), 
	.C1(n1915), 
	.B2(n1914), 
	.B1(n1291), 
	.A2(n1290), 
	.A1(n1913));
   INV_X1 U3120 (.ZN(n5424), 
	.A(\UUT/Mcontrol/d_sampled_finstr [4]));
   INV_X1 U3121 (.ZN(n5422), 
	.A(n1075));
   NAND4_X1 U3122 (.ZN(n1075), 
	.A4(n1919), 
	.A3(n1918), 
	.A2(n1917), 
	.A1(n1916));
   NOR4_X1 U3123 (.ZN(n1919), 
	.A4(n1923), 
	.A3(n1922), 
	.A2(n1921), 
	.A1(n1920));
   NAND3_X1 U3124 (.ZN(n1923), 
	.A3(n5611), 
	.A2(n5609), 
	.A1(n5610));
   OAI211_X1 U3125 (.ZN(n1922), 
	.C2(n5412), 
	.C1(n5560), 
	.B(n5608), 
	.A(n5607));
   OAI222_X1 U3126 (.ZN(n1921), 
	.C2(n5380), 
	.C1(n5561), 
	.B2(n5252), 
	.B1(n5559), 
	.A2(n5284), 
	.A1(n5558));
   OAI221_X1 U3127 (.ZN(n1920), 
	.C2(n5220), 
	.C1(n5532), 
	.B2(n5188), 
	.B1(n5531), 
	.A(n1924));
   AOI22_X1 U3128 (.ZN(n1924), 
	.B2(n1926), 
	.B1(n1276), 
	.A2(n1925), 
	.A1(n1274));
   INV_X1 U3129 (.ZN(n1276), 
	.A(n4996));
   INV_X1 U3130 (.ZN(n1274), 
	.A(n4964));
   AOI211_X1 U3131 (.ZN(n1918), 
	.C2(n1927), 
	.C1(n1278), 
	.B(n1929), 
	.A(n1928));
   OAI22_X1 U3132 (.ZN(n1929), 
	.B2(n4740), 
	.B1(n5551), 
	.A2(n4836), 
	.A1(n5541));
   OAI222_X1 U3133 (.ZN(n1928), 
	.C2(n4708), 
	.C1(n5547), 
	.B2(n4644), 
	.B1(n5552), 
	.A2(n4676), 
	.A1(n5546));
   INV_X1 U3134 (.ZN(n1278), 
	.A(n4868));
   AOI221_X1 U3135 (.ZN(n1917), 
	.C2(n1932), 
	.C1(n1931), 
	.B2(n1285), 
	.B1(n1930), 
	.A(n1933));
   OAI22_X1 U3136 (.ZN(n1933), 
	.B2(n6373), 
	.B1(n5092), 
	.A2(n1934), 
	.A1(n4484));
   INV_X1 U3137 (.ZN(n1932), 
	.A(n5316));
   INV_X1 U3138 (.ZN(n1285), 
	.A(n5348));
   AOI222_X1 U3139 (.ZN(n1916), 
	.C2(n1938), 
	.C1(n1293), 
	.B2(n1292), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1289));
   INV_X1 U3140 (.ZN(n1293), 
	.A(n4516));
   INV_X1 U3141 (.ZN(n1292), 
	.A(n4452));
   INV_X1 U3142 (.ZN(n1289), 
	.A(n4548));
   AND4_X1 U3143 (.ZN(n5421), 
	.A4(n1942), 
	.A3(n1941), 
	.A2(n1940), 
	.A1(n1939));
   NOR4_X1 U3144 (.ZN(n1942), 
	.A4(n1946), 
	.A3(n1945), 
	.A2(n1944), 
	.A1(n1943));
   NAND3_X1 U3145 (.ZN(n1946), 
	.A3(n5604), 
	.A2(n5602), 
	.A1(n5603));
   OAI211_X1 U3146 (.ZN(n1945), 
	.C2(n5396), 
	.C1(n5560), 
	.B(n5601), 
	.A(n5600));
   OAI222_X1 U3147 (.ZN(n1944), 
	.C2(n5364), 
	.C1(n5561), 
	.B2(n5236), 
	.B1(n5559), 
	.A2(n5268), 
	.A1(n5558));
   OAI221_X1 U3148 (.ZN(n1943), 
	.C2(n5204), 
	.C1(n5532), 
	.B2(n5172), 
	.B1(n5531), 
	.A(n1947));
   AOI22_X1 U3149 (.ZN(n1947), 
	.B2(n1926), 
	.B1(n1605), 
	.A2(n1925), 
	.A1(n1604));
   INV_X1 U3150 (.ZN(n1605), 
	.A(n4980));
   INV_X1 U3151 (.ZN(n1604), 
	.A(n4948));
   AOI211_X1 U3152 (.ZN(n1941), 
	.C2(n1927), 
	.C1(n1606), 
	.B(n1949), 
	.A(n1948));
   OAI22_X1 U3153 (.ZN(n1949), 
	.B2(n4724), 
	.B1(n5551), 
	.A2(n4820), 
	.A1(n5541));
   OAI222_X1 U3154 (.ZN(n1948), 
	.C2(n4692), 
	.C1(n5547), 
	.B2(n4628), 
	.B1(n5552), 
	.A2(n4660), 
	.A1(n5546));
   INV_X1 U3155 (.ZN(n1606), 
	.A(n4852));
   AOI221_X1 U3156 (.ZN(n1940), 
	.C2(n1950), 
	.C1(n1931), 
	.B2(n1610), 
	.B1(n1930), 
	.A(n1951));
   OAI22_X1 U3157 (.ZN(n1951), 
	.B2(n6373), 
	.B1(n5076), 
	.A2(n1934), 
	.A1(n4468));
   INV_X1 U3158 (.ZN(n1950), 
	.A(n5300));
   INV_X1 U3159 (.ZN(n1610), 
	.A(n5332));
   AOI222_X1 U3160 (.ZN(n1939), 
	.C2(n1938), 
	.C1(n1614), 
	.B2(n1613), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1612));
   INV_X1 U3161 (.ZN(n1614), 
	.A(n4500));
   INV_X1 U3162 (.ZN(n1613), 
	.A(n4436));
   INV_X1 U3163 (.ZN(n1612), 
	.A(n4532));
   AND4_X1 U3164 (.ZN(n5420), 
	.A4(n1955), 
	.A3(n1954), 
	.A2(n1953), 
	.A1(n1952));
   NOR4_X1 U3165 (.ZN(n1955), 
	.A4(n1959), 
	.A3(n1958), 
	.A2(n1957), 
	.A1(n1956));
   NAND3_X1 U3166 (.ZN(n1959), 
	.A3(n5597), 
	.A2(n5595), 
	.A1(n5596));
   OAI211_X1 U3167 (.ZN(n1958), 
	.C2(n5395), 
	.C1(n5560), 
	.B(n5594), 
	.A(n5593));
   OAI222_X1 U3168 (.ZN(n1957), 
	.C2(n5363), 
	.C1(n5561), 
	.B2(n5235), 
	.B1(n5559), 
	.A2(n5267), 
	.A1(n5558));
   OAI221_X1 U3169 (.ZN(n1956), 
	.C2(n5203), 
	.C1(n5532), 
	.B2(n5171), 
	.B1(n5531), 
	.A(n1960));
   AOI22_X1 U3170 (.ZN(n1960), 
	.B2(n1926), 
	.B1(n1625), 
	.A2(n1925), 
	.A1(n1624));
   INV_X1 U3171 (.ZN(n1625), 
	.A(n4979));
   INV_X1 U3172 (.ZN(n1624), 
	.A(n4947));
   AOI211_X1 U3173 (.ZN(n1954), 
	.C2(n1927), 
	.C1(n1626), 
	.B(n1962), 
	.A(n1961));
   OAI22_X1 U3174 (.ZN(n1962), 
	.B2(n4723), 
	.B1(n5551), 
	.A2(n4819), 
	.A1(n5541));
   OAI222_X1 U3175 (.ZN(n1961), 
	.C2(n4691), 
	.C1(n5547), 
	.B2(n4627), 
	.B1(n5552), 
	.A2(n4659), 
	.A1(n5546));
   INV_X1 U3176 (.ZN(n1626), 
	.A(n4851));
   AOI221_X1 U3177 (.ZN(n1953), 
	.C2(n1963), 
	.C1(n1931), 
	.B2(n1630), 
	.B1(n1930), 
	.A(n1964));
   OAI22_X1 U3178 (.ZN(n1964), 
	.B2(n6373), 
	.B1(n5075), 
	.A2(n1934), 
	.A1(n4467));
   INV_X1 U3179 (.ZN(n1963), 
	.A(n5299));
   INV_X1 U3180 (.ZN(n1630), 
	.A(n5331));
   AOI222_X1 U3181 (.ZN(n1952), 
	.C2(n1938), 
	.C1(n1634), 
	.B2(n1633), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1632));
   INV_X1 U3182 (.ZN(n1634), 
	.A(n4499));
   INV_X1 U3183 (.ZN(n1633), 
	.A(n4435));
   INV_X1 U3184 (.ZN(n1632), 
	.A(n4531));
   AND4_X1 U3185 (.ZN(n5419), 
	.A4(n1968), 
	.A3(n1967), 
	.A2(n1966), 
	.A1(n1965));
   NOR4_X1 U3186 (.ZN(n1968), 
	.A4(n1972), 
	.A3(n1971), 
	.A2(n1970), 
	.A1(n1969));
   NAND3_X1 U3187 (.ZN(n1972), 
	.A3(n5590), 
	.A2(n5588), 
	.A1(n5589));
   OAI211_X1 U3188 (.ZN(n1971), 
	.C2(n5394), 
	.C1(n5560), 
	.B(n5587), 
	.A(n5586));
   OAI222_X1 U3189 (.ZN(n1970), 
	.C2(n5362), 
	.C1(n5561), 
	.B2(n5234), 
	.B1(n5559), 
	.A2(n5266), 
	.A1(n5558));
   OAI221_X1 U3190 (.ZN(n1969), 
	.C2(n5202), 
	.C1(n5532), 
	.B2(n5170), 
	.B1(n5531), 
	.A(n1973));
   AOI22_X1 U3191 (.ZN(n1973), 
	.B2(n1926), 
	.B1(n1645), 
	.A2(n1925), 
	.A1(n1644));
   INV_X1 U3192 (.ZN(n1645), 
	.A(n4978));
   INV_X1 U3193 (.ZN(n1644), 
	.A(n4946));
   AOI211_X1 U3194 (.ZN(n1967), 
	.C2(n1927), 
	.C1(n1646), 
	.B(n1975), 
	.A(n1974));
   OAI22_X1 U3195 (.ZN(n1975), 
	.B2(n4722), 
	.B1(n5551), 
	.A2(n4818), 
	.A1(n5541));
   OAI222_X1 U3196 (.ZN(n1974), 
	.C2(n4690), 
	.C1(n5547), 
	.B2(n4626), 
	.B1(n5552), 
	.A2(n4658), 
	.A1(n5546));
   INV_X1 U3197 (.ZN(n1646), 
	.A(n4850));
   AOI221_X1 U3198 (.ZN(n1966), 
	.C2(n1976), 
	.C1(n1931), 
	.B2(n1650), 
	.B1(n1930), 
	.A(n1977));
   OAI22_X1 U3199 (.ZN(n1977), 
	.B2(n6373), 
	.B1(n5074), 
	.A2(n1934), 
	.A1(n4466));
   INV_X1 U3200 (.ZN(n1976), 
	.A(n5298));
   INV_X1 U3201 (.ZN(n1650), 
	.A(n5330));
   AOI222_X1 U3202 (.ZN(n1965), 
	.C2(n1938), 
	.C1(n1654), 
	.B2(n1653), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1652));
   INV_X1 U3203 (.ZN(n1654), 
	.A(n4498));
   INV_X1 U3204 (.ZN(n1653), 
	.A(n4434));
   INV_X1 U3205 (.ZN(n1652), 
	.A(n4530));
   AND4_X1 U3206 (.ZN(n5418), 
	.A4(n1981), 
	.A3(n1980), 
	.A2(n1979), 
	.A1(n1978));
   NOR4_X1 U3207 (.ZN(n1981), 
	.A4(n1985), 
	.A3(n1984), 
	.A2(n1983), 
	.A1(n1982));
   NAND3_X1 U3208 (.ZN(n1985), 
	.A3(n5583), 
	.A2(n5581), 
	.A1(n5582));
   OAI211_X1 U3209 (.ZN(n1984), 
	.C2(n5393), 
	.C1(n5560), 
	.B(n5580), 
	.A(n5579));
   OAI222_X1 U3210 (.ZN(n1983), 
	.C2(n5361), 
	.C1(n5561), 
	.B2(n5233), 
	.B1(n5559), 
	.A2(n5265), 
	.A1(n5558));
   OAI221_X1 U3211 (.ZN(n1982), 
	.C2(n5201), 
	.C1(n5532), 
	.B2(n5169), 
	.B1(n5531), 
	.A(n1986));
   AOI22_X1 U3212 (.ZN(n1986), 
	.B2(n1926), 
	.B1(n1665), 
	.A2(n1925), 
	.A1(n1664));
   INV_X1 U3213 (.ZN(n1665), 
	.A(n4977));
   INV_X1 U3214 (.ZN(n1664), 
	.A(n4945));
   AOI211_X1 U3215 (.ZN(n1980), 
	.C2(n1927), 
	.C1(n1666), 
	.B(n1988), 
	.A(n1987));
   OAI22_X1 U3216 (.ZN(n1988), 
	.B2(n4721), 
	.B1(n5551), 
	.A2(n4817), 
	.A1(n5541));
   OAI222_X1 U3217 (.ZN(n1987), 
	.C2(n4689), 
	.C1(n5547), 
	.B2(n4625), 
	.B1(n5552), 
	.A2(n4657), 
	.A1(n5546));
   INV_X1 U3218 (.ZN(n1666), 
	.A(n4849));
   AOI221_X1 U3219 (.ZN(n1979), 
	.C2(n1989), 
	.C1(n1931), 
	.B2(n1670), 
	.B1(n1930), 
	.A(n1990));
   OAI22_X1 U3220 (.ZN(n1990), 
	.B2(n6373), 
	.B1(n5073), 
	.A2(n1934), 
	.A1(n4465));
   INV_X1 U3221 (.ZN(n1989), 
	.A(n5297));
   INV_X1 U3222 (.ZN(n1670), 
	.A(n5329));
   AOI222_X1 U3223 (.ZN(n1978), 
	.C2(n1938), 
	.C1(n1674), 
	.B2(n1673), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1672));
   INV_X1 U3224 (.ZN(n1674), 
	.A(n4497));
   INV_X1 U3225 (.ZN(n1673), 
	.A(n4433));
   INV_X1 U3226 (.ZN(n1672), 
	.A(n4529));
   AND4_X1 U3227 (.ZN(n5417), 
	.A4(n1994), 
	.A3(n1993), 
	.A2(n1992), 
	.A1(n1991));
   NOR4_X1 U3228 (.ZN(n1994), 
	.A4(n1998), 
	.A3(n1997), 
	.A2(n1996), 
	.A1(n1995));
   NAND3_X1 U3229 (.ZN(n1998), 
	.A3(n5576), 
	.A2(n5574), 
	.A1(n5575));
   OAI211_X1 U3230 (.ZN(n1997), 
	.C2(n5392), 
	.C1(n5560), 
	.B(n5573), 
	.A(n5572));
   OAI222_X1 U3231 (.ZN(n1996), 
	.C2(n5360), 
	.C1(n5561), 
	.B2(n5232), 
	.B1(n5559), 
	.A2(n5264), 
	.A1(n5558));
   OAI221_X1 U3232 (.ZN(n1995), 
	.C2(n5200), 
	.C1(n5532), 
	.B2(n5168), 
	.B1(n5531), 
	.A(n1999));
   AOI22_X1 U3233 (.ZN(n1999), 
	.B2(n1926), 
	.B1(n1685), 
	.A2(n1925), 
	.A1(n1684));
   INV_X1 U3234 (.ZN(n1685), 
	.A(n4976));
   INV_X1 U3235 (.ZN(n1684), 
	.A(n4944));
   AOI211_X1 U3236 (.ZN(n1993), 
	.C2(n1927), 
	.C1(n1686), 
	.B(n2001), 
	.A(n2000));
   OAI22_X1 U3237 (.ZN(n2001), 
	.B2(n4720), 
	.B1(n5551), 
	.A2(n4816), 
	.A1(n5541));
   OAI222_X1 U3238 (.ZN(n2000), 
	.C2(n4688), 
	.C1(n5547), 
	.B2(n4624), 
	.B1(n5552), 
	.A2(n4656), 
	.A1(n5546));
   INV_X1 U3239 (.ZN(n1686), 
	.A(n4848));
   AOI221_X1 U3240 (.ZN(n1992), 
	.C2(n2002), 
	.C1(n1931), 
	.B2(n1690), 
	.B1(n1930), 
	.A(n2003));
   OAI22_X1 U3241 (.ZN(n2003), 
	.B2(n6373), 
	.B1(n5072), 
	.A2(n1934), 
	.A1(n4464));
   INV_X1 U3242 (.ZN(n2002), 
	.A(n5296));
   INV_X1 U3243 (.ZN(n1690), 
	.A(n5328));
   AOI222_X1 U3244 (.ZN(n1991), 
	.C2(n1938), 
	.C1(n1694), 
	.B2(n1693), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1692));
   INV_X1 U3245 (.ZN(n1694), 
	.A(n4496));
   INV_X1 U3246 (.ZN(n1693), 
	.A(n4432));
   INV_X1 U3247 (.ZN(n1692), 
	.A(n4528));
   AND4_X1 U3248 (.ZN(n5416), 
	.A4(n2007), 
	.A3(n2006), 
	.A2(n2005), 
	.A1(n2004));
   NOR4_X1 U3249 (.ZN(n2007), 
	.A4(n2011), 
	.A3(n2010), 
	.A2(n2009), 
	.A1(n2008));
   NAND3_X1 U3250 (.ZN(n2011), 
	.A3(n5569), 
	.A2(n5567), 
	.A1(n5568));
   OAI211_X1 U3251 (.ZN(n2010), 
	.C2(n5391), 
	.C1(n5560), 
	.B(n5566), 
	.A(n5565));
   OAI222_X1 U3252 (.ZN(n2009), 
	.C2(n5359), 
	.C1(n5561), 
	.B2(n5231), 
	.B1(n5559), 
	.A2(n5263), 
	.A1(n5558));
   OAI221_X1 U3253 (.ZN(n2008), 
	.C2(n5199), 
	.C1(n5532), 
	.B2(n5167), 
	.B1(n5531), 
	.A(n2012));
   AOI22_X1 U3254 (.ZN(n2012), 
	.B2(n1926), 
	.B1(n1705), 
	.A2(n1925), 
	.A1(n1704));
   INV_X1 U3255 (.ZN(n1705), 
	.A(n4975));
   INV_X1 U3256 (.ZN(n1704), 
	.A(n4943));
   AOI211_X1 U3257 (.ZN(n2006), 
	.C2(n1927), 
	.C1(n1706), 
	.B(n2014), 
	.A(n2013));
   OAI22_X1 U3258 (.ZN(n2014), 
	.B2(n4719), 
	.B1(n5551), 
	.A2(n4815), 
	.A1(n5541));
   OAI222_X1 U3259 (.ZN(n2013), 
	.C2(n4687), 
	.C1(n5547), 
	.B2(n4623), 
	.B1(n5552), 
	.A2(n4655), 
	.A1(n5546));
   INV_X1 U3260 (.ZN(n1706), 
	.A(n4847));
   AOI221_X1 U3261 (.ZN(n2005), 
	.C2(n2015), 
	.C1(n1931), 
	.B2(n1710), 
	.B1(n1930), 
	.A(n2016));
   OAI22_X1 U3262 (.ZN(n2016), 
	.B2(n6373), 
	.B1(n5071), 
	.A2(n1934), 
	.A1(n4463));
   INV_X1 U3263 (.ZN(n2015), 
	.A(n5295));
   INV_X1 U3264 (.ZN(n1710), 
	.A(n5327));
   AOI222_X1 U3265 (.ZN(n2004), 
	.C2(n1938), 
	.C1(n1714), 
	.B2(n1713), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1712));
   INV_X1 U3266 (.ZN(n1714), 
	.A(n4495));
   INV_X1 U3267 (.ZN(n1713), 
	.A(n4431));
   INV_X1 U3268 (.ZN(n1712), 
	.A(n4527));
   AND4_X1 U3269 (.ZN(n5415), 
	.A4(n2020), 
	.A3(n2019), 
	.A2(n2018), 
	.A1(n2017));
   NOR4_X1 U3270 (.ZN(n2020), 
	.A4(n2024), 
	.A3(n2023), 
	.A2(n2022), 
	.A1(n2021));
   NAND3_X1 U3271 (.ZN(n2024), 
	.A3(n5555), 
	.A2(n5543), 
	.A1(n5548));
   OAI211_X1 U3272 (.ZN(n2023), 
	.C2(n5389), 
	.C1(n5560), 
	.B(n5538), 
	.A(n5533));
   OAI222_X1 U3273 (.ZN(n2022), 
	.C2(n5357), 
	.C1(n5561), 
	.B2(n5229), 
	.B1(n5559), 
	.A2(n5261), 
	.A1(n5558));
   OAI221_X1 U3274 (.ZN(n2021), 
	.C2(n5197), 
	.C1(n5532), 
	.B2(n5165), 
	.B1(n5531), 
	.A(n2025));
   AOI22_X1 U3275 (.ZN(n2025), 
	.B2(n1926), 
	.B1(n1745), 
	.A2(n1925), 
	.A1(n1744));
   INV_X1 U3276 (.ZN(n1745), 
	.A(n4973));
   INV_X1 U3277 (.ZN(n1744), 
	.A(n4941));
   AOI211_X1 U3278 (.ZN(n2019), 
	.C2(n1927), 
	.C1(n1746), 
	.B(n2027), 
	.A(n2026));
   OAI22_X1 U3279 (.ZN(n2027), 
	.B2(n4717), 
	.B1(n5551), 
	.A2(n4813), 
	.A1(n5541));
   OAI222_X1 U3280 (.ZN(n2026), 
	.C2(n4685), 
	.C1(n5547), 
	.B2(n4621), 
	.B1(n5552), 
	.A2(n4653), 
	.A1(n5546));
   INV_X1 U3281 (.ZN(n1746), 
	.A(n4845));
   AOI221_X1 U3282 (.ZN(n2018), 
	.C2(n2028), 
	.C1(n1931), 
	.B2(n1750), 
	.B1(n1930), 
	.A(n2029));
   OAI22_X1 U3283 (.ZN(n2029), 
	.B2(n6373), 
	.B1(n5069), 
	.A2(n1934), 
	.A1(n4461));
   INV_X1 U3284 (.ZN(n2028), 
	.A(n5293));
   INV_X1 U3285 (.ZN(n1750), 
	.A(n5325));
   AOI222_X1 U3286 (.ZN(n2017), 
	.C2(n1938), 
	.C1(n1754), 
	.B2(n1753), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1752));
   INV_X1 U3287 (.ZN(n1754), 
	.A(n4493));
   INV_X1 U3288 (.ZN(n1753), 
	.A(n4429));
   INV_X1 U3289 (.ZN(n1752), 
	.A(n4525));
   AND4_X1 U3290 (.ZN(n5414), 
	.A4(n2033), 
	.A3(n2032), 
	.A2(n2031), 
	.A1(n2030));
   NOR4_X1 U3291 (.ZN(n2033), 
	.A4(n2037), 
	.A3(n2036), 
	.A2(n2035), 
	.A1(n2034));
   NAND3_X1 U3292 (.ZN(n2037), 
	.A3(n6320), 
	.A2(n6311), 
	.A1(n6315));
   OAI211_X1 U3293 (.ZN(n2036), 
	.C2(n5388), 
	.C1(n5560), 
	.B(n6307), 
	.A(n6300));
   OAI222_X1 U3294 (.ZN(n2035), 
	.C2(n5356), 
	.C1(n5561), 
	.B2(n5228), 
	.B1(n5559), 
	.A2(n5260), 
	.A1(n5558));
   OAI221_X1 U3295 (.ZN(n2034), 
	.C2(n5196), 
	.C1(n5532), 
	.B2(n5164), 
	.B1(n5531), 
	.A(n2038));
   AOI22_X1 U3296 (.ZN(n2038), 
	.B2(n1926), 
	.B1(n1765), 
	.A2(n1925), 
	.A1(n1764));
   INV_X1 U3297 (.ZN(n1765), 
	.A(n4972));
   INV_X1 U3298 (.ZN(n1764), 
	.A(n4940));
   AOI211_X1 U3299 (.ZN(n2032), 
	.C2(n1927), 
	.C1(n1766), 
	.B(n2040), 
	.A(n2039));
   OAI22_X1 U3300 (.ZN(n2040), 
	.B2(n4716), 
	.B1(n5551), 
	.A2(n4812), 
	.A1(n5541));
   OAI222_X1 U3301 (.ZN(n2039), 
	.C2(n4684), 
	.C1(n5547), 
	.B2(n4620), 
	.B1(n5552), 
	.A2(n4652), 
	.A1(n5546));
   INV_X1 U3302 (.ZN(n1766), 
	.A(n4844));
   AOI221_X1 U3303 (.ZN(n2031), 
	.C2(n2041), 
	.C1(n1931), 
	.B2(n1770), 
	.B1(n1930), 
	.A(n2042));
   OAI22_X1 U3304 (.ZN(n2042), 
	.B2(n6373), 
	.B1(n5068), 
	.A2(n1934), 
	.A1(n4460));
   INV_X1 U3305 (.ZN(n2041), 
	.A(n5292));
   INV_X1 U3306 (.ZN(n1770), 
	.A(n5324));
   AOI222_X1 U3307 (.ZN(n2030), 
	.C2(n1938), 
	.C1(n1774), 
	.B2(n1773), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1772));
   INV_X1 U3308 (.ZN(n1774), 
	.A(n4492));
   INV_X1 U3309 (.ZN(n1773), 
	.A(n4428));
   INV_X1 U3310 (.ZN(n1772), 
	.A(n4524));
   NAND2_X1 U3311 (.ZN(dmem_read), 
	.A2(n1059), 
	.A1(\UUT/Mcontrol/bp_logicA/N9 ));
   INV_X1 U3312 (.ZN(n1059), 
	.A(\UUT/Mcontrol/x_sampled_dmem_command[MR] ));
   NAND2_X1 U3313 (.ZN(dmem_ishalf), 
	.A2(n1054), 
	.A1(\UUT/Mcontrol/bp_logicA/N9 ));
   INV_X1 U3314 (.ZN(n1054), 
	.A(\UUT/Mcontrol/x_sampled_dmem_command[MH] ));
   NAND2_X1 U3315 (.ZN(dmem_isbyte), 
	.A2(n1047), 
	.A1(\UUT/Mcontrol/bp_logicA/N9 ));
   INV_X1 U3316 (.ZN(n1047), 
	.A(\UUT/Mcontrol/x_sampled_dmem_command[MB] ));
   NOR2_X1 U3318 (.ZN(\UUT/regfile/N269 ), 
	.A2(n2043), 
	.A1(\UUT/regfile/N267 ));
   INV_X1 U3319 (.ZN(n2043), 
	.A(n6007));
   NAND2_X1 U3320 (.ZN(\UUT/daddr_out [0]), 
	.A2(n2045), 
	.A1(n2044));
   AOI21_X1 U3321 (.ZN(n2045), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[0] ), 
	.A(n2046));
   NOR3_X1 U3322 (.ZN(n2046), 
	.A3(FE_OFN87_n1211), 
	.A2(n2048), 
	.A1(n2047));
   AOI22_X1 U3323 (.ZN(n2048), 
	.B2(n2050), 
	.B1(\UUT/Mpath/the_alu/N91 ), 
	.A2(\UUT/Mpath/the_alu/N93 ), 
	.A1(n2049));
   AND2_X1 U3324 (.ZN(n2049), 
	.A2(\UUT/Mpath/the_alu/N503 ), 
	.A1(\UUT/Mpath/the_alu/N498 ));
   AOI22_X1 U3325 (.ZN(n2044), 
	.B2(n6348), 
	.B1(n6351), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[0] ));
   INV_X1 U3326 (.ZN(\UUT/d_mul_command [5]), 
	.A(n1025));
   NAND2_X1 U3327 (.ZN(n1025), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [5]), 
	.A1(n2051));
   INV_X1 U3328 (.ZN(\UUT/d_mul_command [4]), 
	.A(n1022));
   NAND2_X1 U3329 (.ZN(n1022), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [4]), 
	.A1(n2051));
   NAND2_X1 U3330 (.ZN(\UUT/d_mul_command [3]), 
	.A2(n5425), 
	.A1(n2051));
   NAND2_X1 U3331 (.ZN(\UUT/d_mul_command [2]), 
	.A2(n5426), 
	.A1(n2051));
   NAND2_X1 U3332 (.ZN(\UUT/d_mul_command [1]), 
	.A2(n5427), 
	.A1(n2051));
   NAND2_X1 U3333 (.ZN(\UUT/d_mul_command [0]), 
	.A2(n5428), 
	.A1(n2051));
   AND2_X1 U3334 (.ZN(n2051), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2043 ), 
	.A1(n927));
   INV_X1 U3335 (.ZN(\UUT/byp_controlB[0] ), 
	.A(\UUT/Mcontrol/st_logic/N42 ));
   INV_X1 U3336 (.ZN(\UUT/break_code[23] ), 
	.A(FE_OFN102_n117));
   AOI221_X1 U3337 (.ZN(n117), 
	.C2(n2053), 
	.C1(\UUT/Mcontrol/d_instr [7]), 
	.B2(n2052), 
	.B1(n6093), 
	.A(n2054));
   INV_X1 U3338 (.ZN(\UUT/break_code[22] ), 
	.A(FE_OFN101_n292));
   AOI221_X1 U3339 (.ZN(n292), 
	.C2(\UUT/Mcontrol/d_instr [6]), 
	.C1(n2053), 
	.B2(n2052), 
	.B1(n6101), 
	.A(n2054));
   INV_X1 U3340 (.ZN(\UUT/break_code[21] ), 
	.A(FE_OFN100_n327));
   AOI221_X1 U3341 (.ZN(n327), 
	.C2(n2053), 
	.C1(\UUT/Mcontrol/d_instr [5]), 
	.B2(n2052), 
	.B1(n6108), 
	.A(n2054));
   INV_X1 U3342 (.ZN(\UUT/break_code[20] ), 
	.A(FE_OFN99_n348));
   AOI221_X1 U3343 (.ZN(n348), 
	.C2(n2053), 
	.C1(\UUT/Mcontrol/d_instr [4]), 
	.B2(n2052), 
	.B1(n6115), 
	.A(n2054));
   OAI21_X1 U3344 (.ZN(n2054), 
	.B2(n855), 
	.B1(n1169), 
	.A(n2055));
   INV_X1 U3345 (.ZN(n2055), 
	.A(n448));
   NAND3_X1 U3346 (.ZN(n855), 
	.A3(n857), 
	.A2(n1216), 
	.A1(\UUT/Mcontrol/d_sampled_finstr [15]));
   NOR2_X1 U3347 (.ZN(n2052), 
	.A2(n1169), 
	.A1(n1168));
   INV_X1 U3348 (.ZN(n1168), 
	.A(n1167));
   NOR2_X1 U3349 (.ZN(n1167), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
	.A1(n1216));
   NAND4_X1 U3350 (.ZN(n1216), 
	.A4(\UUT/Mcontrol/Operation_decoding32/N1994 ), 
	.A3(n6042), 
	.A2(n1061), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1987 ));
   INV_X1 U3351 (.ZN(n6042), 
	.A(n1064));
   NOR3_X1 U3352 (.ZN(n1064), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1992 ), 
	.A1(\UUT/Mcontrol/d_instr [27]));
   OAI21_X1 U3353 (.ZN(n1061), 
	.B2(n2056), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.A(n2057));
   NAND3_X1 U3354 (.ZN(n2057), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1993 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2005 ));
   INV_X1 U3355 (.ZN(n2056), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1974 ));
   NAND2_X1 U3356 (.ZN(\UUT/break_code[1] ), 
	.A2(n2059), 
	.A1(n2058));
   NAND3_X1 U3357 (.ZN(n2059), 
	.A3(\UUT/Mcontrol/d_instr [7]), 
	.A2(n935), 
	.A1(n6086));
   NAND2_X1 U3358 (.ZN(n2058), 
	.A2(n2060), 
	.A1(\UUT/Mcontrol/d_instr [1]));
   INV_X1 U3359 (.ZN(n2060), 
	.A(n2061));
   OAI221_X1 U3360 (.ZN(\UUT/break_code[19] ), 
	.C2(n2064), 
	.C1(n5425), 
	.B2(n2063), 
	.B1(n2062), 
	.A(n2065));
   INV_X1 U3361 (.ZN(n5425), 
	.A(\UUT/Mcontrol/d_sampled_finstr [3]));
   INV_X1 U3362 (.ZN(n2063), 
	.A(n6126));
   OAI221_X1 U3363 (.ZN(\UUT/break_code[18] ), 
	.C2(n2064), 
	.C1(n5426), 
	.B2(n2066), 
	.B1(n2062), 
	.A(n2065));
   INV_X1 U3364 (.ZN(n5426), 
	.A(\UUT/Mcontrol/d_sampled_finstr [2]));
   INV_X1 U3365 (.ZN(n2066), 
	.A(n6135));
   OAI221_X1 U3366 (.ZN(\UUT/break_code[17] ), 
	.C2(n2064), 
	.C1(n5427), 
	.B2(n2067), 
	.B1(n2062), 
	.A(n2065));
   INV_X1 U3367 (.ZN(n5427), 
	.A(\UUT/Mcontrol/d_sampled_finstr [1]));
   INV_X1 U3368 (.ZN(n2067), 
	.A(n6153));
   OAI221_X1 U3369 (.ZN(\UUT/break_code[16] ), 
	.C2(n2064), 
	.C1(n5428), 
	.B2(n2068), 
	.B1(n2062), 
	.A(n2065));
   AOI21_X1 U3370 (.ZN(n2065), 
	.B2(n6127), 
	.B1(n6050), 
	.A(n448));
   NOR3_X1 U3371 (.ZN(n448), 
	.A3(n929), 
	.A2(n5831), 
	.A1(n933));
   INV_X1 U3372 (.ZN(n2064), 
	.A(n2053));
   NOR2_X1 U3373 (.ZN(n2053), 
	.A2(n1169), 
	.A1(n857));
   INV_X1 U3374 (.ZN(n857), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2025 ));
   INV_X1 U3375 (.ZN(n5428), 
	.A(\UUT/Mcontrol/d_sampled_finstr [0]));
   INV_X1 U3376 (.ZN(n2068), 
	.A(n6162));
   NAND2_X1 U3377 (.ZN(n2062), 
	.A2(n445), 
	.A1(n6050));
   NOR2_X1 U3378 (.ZN(n6050), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
	.A1(n1169));
   NAND2_X1 U3379 (.ZN(n1169), 
	.A2(n931), 
	.A1(n927));
   INV_X1 U3381 (.ZN(n943), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2030 ));
   NOR2_X1 U3382 (.ZN(n927), 
	.A2(n6170), 
	.A1(n933));
   INV_X1 U3383 (.ZN(\UUT/break_code[15] ), 
	.A(n466));
   NAND2_X1 U3384 (.ZN(n466), 
	.A2(n6030), 
	.A1(n2069));
   OAI22_X1 U3385 (.ZN(n2069), 
	.B2(n2071), 
	.B1(n5831), 
	.A2(n2070), 
	.A1(n6173));
   INV_X1 U3386 (.ZN(n2071), 
	.A(n6170));
   INV_X1 U3387 (.ZN(n5831), 
	.A(\UUT/Mcontrol/d_sampled_finstr [15]));
   OAI21_X1 U3388 (.ZN(\UUT/break_code[14] ), 
	.B2(n2072), 
	.B1(n6032), 
	.A(n2073));
   NAND2_X1 U3389 (.ZN(n2073), 
	.A2(n2074), 
	.A1(n6181));
   INV_X1 U3390 (.ZN(n6032), 
	.A(\UUT/Mcontrol/d_sampled_finstr [14]));
   OAI21_X1 U3391 (.ZN(\UUT/break_code[13] ), 
	.B2(n2072), 
	.B1(n6033), 
	.A(n2075));
   NAND2_X1 U3392 (.ZN(n2075), 
	.A2(n2074), 
	.A1(n6188));
   INV_X1 U3393 (.ZN(n6033), 
	.A(\UUT/Mcontrol/d_sampled_finstr [13]));
   OAI21_X1 U3394 (.ZN(\UUT/break_code[0] ), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N1901 ), 
	.B1(n2061), 
	.A(n2076));
   NOR2_X1 U3397 (.ZN(n935), 
	.A2(n933), 
	.A1(n2077));
   AOI222_X1 U3399 (.ZN(n5480), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[23] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n878), 
	.A2(n5564), 
	.A1(n6092));
   NAND2_X1 U3400 (.ZN(n878), 
	.A2(n2080), 
	.A1(n2079));
   AOI222_X1 U3401 (.ZN(n2080), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [23]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [23]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [23]));
   AOI22_X1 U3402 (.ZN(n2079), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [23]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [23]));
   NAND3_X1 U3403 (.ZN(n6092), 
	.A3(n2083), 
	.A2(n2082), 
	.A1(n2081));
   AOI222_X1 U3404 (.ZN(n2083), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[23] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[23] ), 
	.A2(n2084), 
	.A1(n1208));
   INV_X1 U3405 (.ZN(n2084), 
	.A(\UUT/Mpath/the_alu/N37 ));
   AOI22_X1 U3406 (.ZN(n2082), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N102 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N134 ));
   AOI22_X1 U3407 (.ZN(n2081), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N198 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N166 ));
   INV_X1 U3408 (.ZN(n2078), 
	.A(n811));
   NAND4_X1 U3409 (.ZN(n811), 
	.A4(n2088), 
	.A3(n2087), 
	.A2(n2086), 
	.A1(n2085));
   NOR4_X1 U3410 (.ZN(n2088), 
	.A4(n2092), 
	.A3(n2091), 
	.A2(n2090), 
	.A1(n2089));
   NAND3_X1 U3411 (.ZN(n2092), 
	.A3(n6091), 
	.A2(n6089), 
	.A1(n6090));
   OAI211_X1 U3412 (.ZN(n2091), 
	.C2(n5397), 
	.C1(n5560), 
	.B(n6088), 
	.A(n6087));
   OAI222_X1 U3413 (.ZN(n2090), 
	.C2(n5365), 
	.C1(n5561), 
	.B2(n5237), 
	.B1(n5559), 
	.A2(n5269), 
	.A1(n5558));
   OAI221_X1 U3414 (.ZN(n2089), 
	.C2(n5205), 
	.C1(n5532), 
	.B2(n5173), 
	.B1(n5531), 
	.A(n2093));
   AOI22_X1 U3415 (.ZN(n2093), 
	.B2(n1926), 
	.B1(n1585), 
	.A2(n1925), 
	.A1(n1584));
   INV_X1 U3416 (.ZN(n1585), 
	.A(n4981));
   INV_X1 U3417 (.ZN(n1584), 
	.A(n4949));
   AOI211_X1 U3418 (.ZN(n2087), 
	.C2(n1927), 
	.C1(n1586), 
	.B(n2095), 
	.A(n2094));
   OAI22_X1 U3419 (.ZN(n2095), 
	.B2(n4725), 
	.B1(n5551), 
	.A2(n4821), 
	.A1(n5541));
   OAI222_X1 U3420 (.ZN(n2094), 
	.C2(n4693), 
	.C1(n5547), 
	.B2(n4629), 
	.B1(n5552), 
	.A2(n4661), 
	.A1(n5546));
   INV_X1 U3421 (.ZN(n1586), 
	.A(n4853));
   AOI221_X1 U3422 (.ZN(n2086), 
	.C2(n2096), 
	.C1(n1931), 
	.B2(n1590), 
	.B1(n1930), 
	.A(n2097));
   OAI22_X1 U3423 (.ZN(n2097), 
	.B2(n6373), 
	.B1(n5077), 
	.A2(n1934), 
	.A1(n4469));
   INV_X1 U3424 (.ZN(n2096), 
	.A(n5301));
   INV_X1 U3425 (.ZN(n1590), 
	.A(n5333));
   AOI222_X1 U3426 (.ZN(n2085), 
	.C2(n1938), 
	.C1(n1594), 
	.B2(n1593), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1592));
   INV_X1 U3427 (.ZN(n1594), 
	.A(n4501));
   INV_X1 U3428 (.ZN(n1593), 
	.A(n4437));
   INV_X1 U3429 (.ZN(n1592), 
	.A(n4533));
   AOI222_X1 U3431 (.ZN(n5483), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[22] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n324), 
	.A2(n5564), 
	.A1(n6100));
   NAND2_X1 U3432 (.ZN(n324), 
	.A2(n2100), 
	.A1(n2099));
   AOI222_X1 U3433 (.ZN(n2100), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [22]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [22]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [22]));
   AOI22_X1 U3434 (.ZN(n2099), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [22]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [22]));
   NAND3_X1 U3435 (.ZN(n6100), 
	.A3(n2103), 
	.A2(n2102), 
	.A1(n2101));
   AOI222_X1 U3436 (.ZN(n2103), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[22] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[22] ), 
	.A2(n2104), 
	.A1(n1208));
   INV_X1 U3437 (.ZN(n2104), 
	.A(\UUT/Mpath/the_alu/N39 ));
   AOI22_X1 U3438 (.ZN(n2102), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N103 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N135 ));
   AOI22_X1 U3439 (.ZN(n2101), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N199 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N167 ));
   INV_X1 U3440 (.ZN(n2098), 
	.A(n313));
   NAND4_X1 U3441 (.ZN(n313), 
	.A4(n2108), 
	.A3(n2107), 
	.A2(n2106), 
	.A1(n2105));
   NOR4_X1 U3442 (.ZN(n2108), 
	.A4(n2112), 
	.A3(n2111), 
	.A2(n2110), 
	.A1(n2109));
   NAND3_X1 U3443 (.ZN(n2112), 
	.A3(n6099), 
	.A2(n6097), 
	.A1(n6098));
   OAI211_X1 U3444 (.ZN(n2111), 
	.C2(n5398), 
	.C1(n5560), 
	.B(n6096), 
	.A(n6095));
   OAI222_X1 U3445 (.ZN(n2110), 
	.C2(n5366), 
	.C1(n5561), 
	.B2(n5238), 
	.B1(n5559), 
	.A2(n5270), 
	.A1(n5558));
   OAI221_X1 U3446 (.ZN(n2109), 
	.C2(n5206), 
	.C1(n5532), 
	.B2(n5174), 
	.B1(n5531), 
	.A(n2113));
   AOI22_X1 U3447 (.ZN(n2113), 
	.B2(n1926), 
	.B1(n1565), 
	.A2(n1925), 
	.A1(n1564));
   INV_X1 U3448 (.ZN(n1565), 
	.A(n4982));
   INV_X1 U3449 (.ZN(n1564), 
	.A(n4950));
   AOI211_X1 U3450 (.ZN(n2107), 
	.C2(n1927), 
	.C1(n1566), 
	.B(n2115), 
	.A(n2114));
   OAI22_X1 U3451 (.ZN(n2115), 
	.B2(n4726), 
	.B1(n5551), 
	.A2(n4822), 
	.A1(n5541));
   OAI222_X1 U3452 (.ZN(n2114), 
	.C2(n4694), 
	.C1(n5547), 
	.B2(n4630), 
	.B1(n5552), 
	.A2(n4662), 
	.A1(n5546));
   INV_X1 U3453 (.ZN(n1566), 
	.A(n4854));
   AOI221_X1 U3454 (.ZN(n2106), 
	.C2(n2116), 
	.C1(n1931), 
	.B2(n1570), 
	.B1(n1930), 
	.A(n2117));
   OAI22_X1 U3455 (.ZN(n2117), 
	.B2(n6373), 
	.B1(n5078), 
	.A2(n1934), 
	.A1(n4470));
   INV_X1 U3456 (.ZN(n2116), 
	.A(n5302));
   INV_X1 U3457 (.ZN(n1570), 
	.A(n5334));
   AOI222_X1 U3458 (.ZN(n2105), 
	.C2(n1938), 
	.C1(n1574), 
	.B2(n1573), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1572));
   INV_X1 U3459 (.ZN(n1574), 
	.A(n4502));
   INV_X1 U3460 (.ZN(n1573), 
	.A(n4438));
   INV_X1 U3461 (.ZN(n1572), 
	.A(n4534));
   OAI222_X1 U3462 (.ZN(\UUT/branch_rega [21]), 
	.C2(n5486), 
	.C1(n5528), 
	.B2(n2118), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5488));
   NAND2_X1 U3464 (.ZN(n346), 
	.A2(n2120), 
	.A1(n2119));
   AOI222_X1 U3465 (.ZN(n2120), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [21]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [21]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [21]));
   AOI22_X1 U3466 (.ZN(n2119), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [21]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [21]));
   NAND3_X1 U3467 (.ZN(n6107), 
	.A3(n2123), 
	.A2(n2122), 
	.A1(n2121));
   AOI222_X1 U3468 (.ZN(n2123), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[21] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[21] ), 
	.A2(n2124), 
	.A1(n1208));
   INV_X1 U3469 (.ZN(n2124), 
	.A(\UUT/Mpath/the_alu/N41 ));
   AOI22_X1 U3470 (.ZN(n2122), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N104 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N136 ));
   AOI22_X1 U3471 (.ZN(n2121), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N200 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N168 ));
   INV_X1 U3472 (.ZN(n2118), 
	.A(n340));
   NAND4_X1 U3473 (.ZN(n340), 
	.A4(n2128), 
	.A3(n2127), 
	.A2(n2126), 
	.A1(n2125));
   NOR4_X1 U3474 (.ZN(n2128), 
	.A4(n2132), 
	.A3(n2131), 
	.A2(n2130), 
	.A1(n2129));
   NAND3_X1 U3475 (.ZN(n2132), 
	.A3(n6106), 
	.A2(n6104), 
	.A1(n6105));
   OAI211_X1 U3476 (.ZN(n2131), 
	.C2(n5399), 
	.C1(n5560), 
	.B(n6103), 
	.A(n6102));
   OAI222_X1 U3477 (.ZN(n2130), 
	.C2(n5367), 
	.C1(n5561), 
	.B2(n5239), 
	.B1(n5559), 
	.A2(n5271), 
	.A1(n5558));
   OAI221_X1 U3478 (.ZN(n2129), 
	.C2(n5207), 
	.C1(n5532), 
	.B2(n5175), 
	.B1(n5531), 
	.A(n2133));
   AOI22_X1 U3479 (.ZN(n2133), 
	.B2(n1926), 
	.B1(n1545), 
	.A2(n1925), 
	.A1(n1544));
   INV_X1 U3480 (.ZN(n1545), 
	.A(n4983));
   INV_X1 U3481 (.ZN(n1544), 
	.A(n4951));
   AOI211_X1 U3482 (.ZN(n2127), 
	.C2(n1927), 
	.C1(n1546), 
	.B(n2135), 
	.A(n2134));
   OAI22_X1 U3483 (.ZN(n2135), 
	.B2(n4727), 
	.B1(n5551), 
	.A2(n4823), 
	.A1(n5541));
   OAI222_X1 U3484 (.ZN(n2134), 
	.C2(n4695), 
	.C1(n5547), 
	.B2(n4631), 
	.B1(n5552), 
	.A2(n4663), 
	.A1(n5546));
   INV_X1 U3485 (.ZN(n1546), 
	.A(n4855));
   AOI221_X1 U3486 (.ZN(n2126), 
	.C2(n2136), 
	.C1(n1931), 
	.B2(n1550), 
	.B1(n1930), 
	.A(n2137));
   OAI22_X1 U3487 (.ZN(n2137), 
	.B2(n6373), 
	.B1(n5079), 
	.A2(n1934), 
	.A1(n4471));
   INV_X1 U3488 (.ZN(n2136), 
	.A(n5303));
   INV_X1 U3489 (.ZN(n1550), 
	.A(n5335));
   AOI222_X1 U3490 (.ZN(n2125), 
	.C2(n1938), 
	.C1(n1554), 
	.B2(n1553), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1552));
   INV_X1 U3491 (.ZN(n1554), 
	.A(n4503));
   INV_X1 U3492 (.ZN(n1553), 
	.A(n4439));
   INV_X1 U3493 (.ZN(n1552), 
	.A(n4535));
   OAI222_X1 U3494 (.ZN(\UUT/branch_rega [20]), 
	.C2(n5489), 
	.C1(n5528), 
	.B2(n2138), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5491));
   AOI222_X1 U3495 (.ZN(n5489), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[20] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n367), 
	.A2(n5564), 
	.A1(n6114));
   NAND2_X1 U3496 (.ZN(n367), 
	.A2(n2140), 
	.A1(n2139));
   AOI222_X1 U3497 (.ZN(n2140), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [20]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [20]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [20]));
   AOI22_X1 U3498 (.ZN(n2139), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [20]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [20]));
   NAND3_X1 U3499 (.ZN(n6114), 
	.A3(n2143), 
	.A2(n2142), 
	.A1(n2141));
   AOI222_X1 U3500 (.ZN(n2143), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[20] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[20] ), 
	.A2(n2144), 
	.A1(n1208));
   INV_X1 U3501 (.ZN(n2144), 
	.A(\UUT/Mpath/the_alu/N43 ));
   AOI22_X1 U3502 (.ZN(n2142), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N105 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N137 ));
   AOI22_X1 U3503 (.ZN(n2141), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N201 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N169 ));
   INV_X1 U3504 (.ZN(n2138), 
	.A(n361));
   NAND4_X1 U3505 (.ZN(n361), 
	.A4(n2148), 
	.A3(n2147), 
	.A2(n2146), 
	.A1(n2145));
   NOR4_X1 U3506 (.ZN(n2148), 
	.A4(n2152), 
	.A3(n2151), 
	.A2(n2150), 
	.A1(n2149));
   NAND3_X1 U3507 (.ZN(n2152), 
	.A3(n6113), 
	.A2(n6111), 
	.A1(n6112));
   OAI211_X1 U3508 (.ZN(n2151), 
	.C2(n5400), 
	.C1(n5560), 
	.B(n6110), 
	.A(n6109));
   OAI222_X1 U3509 (.ZN(n2150), 
	.C2(n5368), 
	.C1(n5561), 
	.B2(n5240), 
	.B1(n5559), 
	.A2(n5272), 
	.A1(n5558));
   OAI221_X1 U3510 (.ZN(n2149), 
	.C2(n5208), 
	.C1(n5532), 
	.B2(n5176), 
	.B1(n5531), 
	.A(n2153));
   AOI22_X1 U3511 (.ZN(n2153), 
	.B2(n1926), 
	.B1(n1525), 
	.A2(n1925), 
	.A1(n1524));
   INV_X1 U3512 (.ZN(n1525), 
	.A(n4984));
   INV_X1 U3513 (.ZN(n1524), 
	.A(n4952));
   AOI211_X1 U3514 (.ZN(n2147), 
	.C2(n1927), 
	.C1(n1526), 
	.B(n2155), 
	.A(n2154));
   OAI22_X1 U3515 (.ZN(n2155), 
	.B2(n4728), 
	.B1(n5551), 
	.A2(n4824), 
	.A1(n5541));
   OAI222_X1 U3516 (.ZN(n2154), 
	.C2(n4696), 
	.C1(n5547), 
	.B2(n4632), 
	.B1(n5552), 
	.A2(n4664), 
	.A1(n5546));
   INV_X1 U3517 (.ZN(n1526), 
	.A(n4856));
   AOI221_X1 U3518 (.ZN(n2146), 
	.C2(n2156), 
	.C1(n1931), 
	.B2(n1530), 
	.B1(n1930), 
	.A(n2157));
   OAI22_X1 U3519 (.ZN(n2157), 
	.B2(n6373), 
	.B1(n5080), 
	.A2(n1934), 
	.A1(n4472));
   INV_X1 U3520 (.ZN(n2156), 
	.A(n5304));
   INV_X1 U3521 (.ZN(n1530), 
	.A(n5336));
   AOI222_X1 U3522 (.ZN(n2145), 
	.C2(n1938), 
	.C1(n1534), 
	.B2(n1533), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1532));
   INV_X1 U3523 (.ZN(n1534), 
	.A(n4504));
   INV_X1 U3524 (.ZN(n1533), 
	.A(n4440));
   INV_X1 U3525 (.ZN(n1532), 
	.A(n4536));
   OAI222_X1 U3526 (.ZN(\UUT/branch_rega [1]), 
	.C2(FE_OFN188_n5492), 
	.C1(n5528), 
	.B2(n2158), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5494));
   AOI222_X1 U3527 (.ZN(n5492), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[1] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n822), 
	.A2(n5564), 
	.A1(\UUT/daddr_out [1]));
   NAND2_X1 U3528 (.ZN(n822), 
	.A2(n2160), 
	.A1(n2159));
   AOI222_X1 U3529 (.ZN(n2160), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [1]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [1]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [1]));
   AOI22_X1 U3530 (.ZN(n2159), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [1]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [1]));
   OAI211_X1 U3531 (.ZN(\UUT/daddr_out [1]), 
	.C2(n2161), 
	.C1(\UUT/Mpath/the_alu/N81 ), 
	.B(n2163), 
	.A(n2162));
   AOI22_X1 U3532 (.ZN(n2163), 
	.B2(FE_OFN87_n1211), 
	.B1(\UUT/Mpath/the_alu/sum[1] ), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[1] ));
   AOI22_X1 U3533 (.ZN(n2162), 
	.B2(n2166), 
	.B1(n2165), 
	.A2(\UUT/Mpath/the_alu/N82 ), 
	.A1(n2164));
   INV_X1 U3534 (.ZN(n2165), 
	.A(n2167));
   AOI21_X1 U3535 (.ZN(n2167), 
	.B2(\UUT/Mpath/the_alu/N81 ), 
	.B1(FE_OFN86_n1214), 
	.A(n1212));
   AND2_X1 U3536 (.ZN(n2164), 
	.A2(\UUT/Mpath/the_alu/N81 ), 
	.A1(n1215));
   NOR3_X1 U3537 (.ZN(n2161), 
	.A3(n1212), 
	.A2(n1208), 
	.A1(n2168));
   INV_X1 U3538 (.ZN(n2168), 
	.A(n2169));
   AOI22_X1 U3539 (.ZN(n2169), 
	.B2(n1213), 
	.B1(n2166), 
	.A2(\UUT/Mpath/the_alu/N82 ), 
	.A1(FE_OFN86_n1214));
   INV_X1 U3540 (.ZN(n2166), 
	.A(\UUT/Mpath/the_alu/N82 ));
   INV_X1 U3541 (.ZN(n2158), 
	.A(n799));
   NAND4_X1 U3542 (.ZN(n799), 
	.A4(FE_OFN85_n2173), 
	.A3(n2172), 
	.A2(n2171), 
	.A1(n2170));
   NOR4_X1 U3543 (.ZN(n2173), 
	.A4(n2177), 
	.A3(n2176), 
	.A2(n2175), 
	.A1(n2174));
   NAND3_X1 U3544 (.ZN(n2177), 
	.A3(n6084), 
	.A2(n6082), 
	.A1(n6083));
   OAI211_X1 U3545 (.ZN(n2176), 
	.C2(n5401), 
	.C1(n5560), 
	.B(n6081), 
	.A(n6080));
   OAI222_X1 U3546 (.ZN(n2175), 
	.C2(n5369), 
	.C1(n5561), 
	.B2(n5241), 
	.B1(n5559), 
	.A2(n5273), 
	.A1(n5558));
   OAI221_X1 U3547 (.ZN(n2174), 
	.C2(n5209), 
	.C1(n5532), 
	.B2(n5177), 
	.B1(n5531), 
	.A(n2178));
   AOI22_X1 U3548 (.ZN(n2178), 
	.B2(n1926), 
	.B1(n1505), 
	.A2(n1925), 
	.A1(n1504));
   INV_X1 U3549 (.ZN(n1505), 
	.A(n4985));
   INV_X1 U3550 (.ZN(n1504), 
	.A(n4953));
   AOI211_X1 U3551 (.ZN(n2172), 
	.C2(n1927), 
	.C1(n1506), 
	.B(n2180), 
	.A(n2179));
   OAI22_X1 U3552 (.ZN(n2180), 
	.B2(n4729), 
	.B1(n5551), 
	.A2(n4825), 
	.A1(n5541));
   OAI222_X1 U3553 (.ZN(n2179), 
	.C2(n4697), 
	.C1(n5547), 
	.B2(n4633), 
	.B1(n5552), 
	.A2(n4665), 
	.A1(n5546));
   INV_X1 U3554 (.ZN(n1506), 
	.A(n4857));
   AOI221_X1 U3555 (.ZN(n2171), 
	.C2(n2181), 
	.C1(n1931), 
	.B2(n1510), 
	.B1(n1930), 
	.A(n2182));
   OAI22_X1 U3556 (.ZN(n2182), 
	.B2(n6373), 
	.B1(n5081), 
	.A2(n1934), 
	.A1(n4473));
   INV_X1 U3557 (.ZN(n2181), 
	.A(n5305));
   INV_X1 U3558 (.ZN(n1510), 
	.A(n5337));
   AOI222_X1 U3559 (.ZN(n2170), 
	.C2(n1938), 
	.C1(n1514), 
	.B2(n1513), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1512));
   INV_X1 U3560 (.ZN(n1514), 
	.A(n4505));
   INV_X1 U3561 (.ZN(n1513), 
	.A(n4441));
   INV_X1 U3562 (.ZN(n1512), 
	.A(n4537));
   OAI222_X1 U3563 (.ZN(\UUT/branch_rega [19]), 
	.C2(n5495), 
	.C1(n5528), 
	.B2(n2183), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5497));
   AOI222_X1 U3564 (.ZN(n5495), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[19] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n393), 
	.A2(n5564), 
	.A1(n6124));
   NAND2_X1 U3565 (.ZN(n393), 
	.A2(n2185), 
	.A1(n2184));
   AOI222_X1 U3566 (.ZN(n2185), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [19]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [19]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [19]));
   AOI22_X1 U3567 (.ZN(n2184), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [19]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [19]));
   NAND3_X1 U3568 (.ZN(n6124), 
	.A3(n2188), 
	.A2(n2187), 
	.A1(n2186));
   AOI222_X1 U3569 (.ZN(n2188), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[19] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[19] ), 
	.A2(n2189), 
	.A1(n1208));
   INV_X1 U3570 (.ZN(n2189), 
	.A(\UUT/Mpath/the_alu/N45 ));
   AOI22_X1 U3571 (.ZN(n2187), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N106 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N138 ));
   AOI22_X1 U3572 (.ZN(n2186), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N202 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N170 ));
   INV_X1 U3573 (.ZN(n2183), 
	.A(n387));
   NAND4_X1 U3574 (.ZN(n387), 
	.A4(n2193), 
	.A3(n2192), 
	.A2(n2191), 
	.A1(n2190));
   NOR4_X1 U3575 (.ZN(n2193), 
	.A4(n2197), 
	.A3(n2196), 
	.A2(n2195), 
	.A1(n2194));
   NAND3_X1 U3576 (.ZN(n2197), 
	.A3(n6123), 
	.A2(n6121), 
	.A1(n6122));
   OAI211_X1 U3577 (.ZN(n2196), 
	.C2(n5402), 
	.C1(n5560), 
	.B(n6120), 
	.A(n6119));
   OAI222_X1 U3578 (.ZN(n2195), 
	.C2(n5370), 
	.C1(n5561), 
	.B2(n5242), 
	.B1(n5559), 
	.A2(n5274), 
	.A1(n5558));
   OAI221_X1 U3579 (.ZN(n2194), 
	.C2(n5210), 
	.C1(n5532), 
	.B2(n5178), 
	.B1(n5531), 
	.A(n2198));
   AOI22_X1 U3580 (.ZN(n2198), 
	.B2(n1926), 
	.B1(n1485), 
	.A2(n1925), 
	.A1(n1484));
   INV_X1 U3581 (.ZN(n1485), 
	.A(n4986));
   INV_X1 U3582 (.ZN(n1484), 
	.A(n4954));
   AOI211_X1 U3583 (.ZN(n2192), 
	.C2(n1927), 
	.C1(n1486), 
	.B(n2200), 
	.A(n2199));
   OAI22_X1 U3584 (.ZN(n2200), 
	.B2(n4730), 
	.B1(n5551), 
	.A2(n4826), 
	.A1(n5541));
   OAI222_X1 U3585 (.ZN(n2199), 
	.C2(n4698), 
	.C1(n5547), 
	.B2(n4634), 
	.B1(n5552), 
	.A2(n4666), 
	.A1(n5546));
   INV_X1 U3586 (.ZN(n1486), 
	.A(n4858));
   AOI221_X1 U3587 (.ZN(n2191), 
	.C2(n2201), 
	.C1(n1931), 
	.B2(n1490), 
	.B1(n1930), 
	.A(n2202));
   OAI22_X1 U3588 (.ZN(n2202), 
	.B2(n6373), 
	.B1(n5082), 
	.A2(n1934), 
	.A1(n4474));
   INV_X1 U3589 (.ZN(n2201), 
	.A(n5306));
   INV_X1 U3590 (.ZN(n1490), 
	.A(n5338));
   AOI222_X1 U3591 (.ZN(n2190), 
	.C2(n1938), 
	.C1(n1494), 
	.B2(n1493), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1492));
   INV_X1 U3592 (.ZN(n1494), 
	.A(n4506));
   INV_X1 U3593 (.ZN(n1493), 
	.A(n4442));
   INV_X1 U3594 (.ZN(n1492), 
	.A(n4538));
   NAND2_X1 U3597 (.ZN(n415), 
	.A2(n2205), 
	.A1(n2204));
   AOI222_X1 U3598 (.ZN(n2205), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [18]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [18]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [18]));
   AOI22_X1 U3599 (.ZN(n2204), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [18]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [18]));
   NAND3_X1 U3600 (.ZN(n6134), 
	.A3(n2208), 
	.A2(n2207), 
	.A1(n2206));
   AOI222_X1 U3601 (.ZN(n2208), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[18] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[18] ), 
	.A2(n2209), 
	.A1(n1208));
   INV_X1 U3602 (.ZN(n2209), 
	.A(\UUT/Mpath/the_alu/N47 ));
   AOI22_X1 U3603 (.ZN(n2207), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N107 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N139 ));
   AOI22_X1 U3604 (.ZN(n2206), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N203 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N171 ));
   INV_X1 U3605 (.ZN(n2203), 
	.A(n409));
   NAND4_X1 U3606 (.ZN(n409), 
	.A4(n2213), 
	.A3(n2212), 
	.A2(n2211), 
	.A1(n2210));
   NOR4_X1 U3607 (.ZN(n2213), 
	.A4(n2217), 
	.A3(n2216), 
	.A2(n2215), 
	.A1(n2214));
   NAND3_X1 U3608 (.ZN(n2217), 
	.A3(n6133), 
	.A2(n6131), 
	.A1(n6132));
   OAI211_X1 U3609 (.ZN(n2216), 
	.C2(n5403), 
	.C1(n5560), 
	.B(n6130), 
	.A(n6129));
   OAI222_X1 U3610 (.ZN(n2215), 
	.C2(n5371), 
	.C1(n5561), 
	.B2(n5243), 
	.B1(n5559), 
	.A2(n5275), 
	.A1(n5558));
   OAI221_X1 U3611 (.ZN(n2214), 
	.C2(n5211), 
	.C1(n5532), 
	.B2(n5179), 
	.B1(n5531), 
	.A(n2218));
   AOI22_X1 U3612 (.ZN(n2218), 
	.B2(n1926), 
	.B1(n1465), 
	.A2(n1925), 
	.A1(n1464));
   INV_X1 U3613 (.ZN(n1465), 
	.A(n4987));
   INV_X1 U3614 (.ZN(n1464), 
	.A(n4955));
   AOI211_X1 U3615 (.ZN(n2212), 
	.C2(n1927), 
	.C1(n1466), 
	.B(n2220), 
	.A(n2219));
   OAI22_X1 U3616 (.ZN(n2220), 
	.B2(n4731), 
	.B1(n5551), 
	.A2(n4827), 
	.A1(n5541));
   OAI222_X1 U3617 (.ZN(n2219), 
	.C2(n4699), 
	.C1(n5547), 
	.B2(n4635), 
	.B1(n5552), 
	.A2(n4667), 
	.A1(n5546));
   INV_X1 U3618 (.ZN(n1466), 
	.A(n4859));
   AOI221_X1 U3619 (.ZN(n2211), 
	.C2(n2221), 
	.C1(n1931), 
	.B2(n1470), 
	.B1(n1930), 
	.A(n2222));
   OAI22_X1 U3620 (.ZN(n2222), 
	.B2(n6373), 
	.B1(n5083), 
	.A2(n1934), 
	.A1(n4475));
   INV_X1 U3621 (.ZN(n2221), 
	.A(n5307));
   INV_X1 U3622 (.ZN(n1470), 
	.A(n5339));
   AOI222_X1 U3623 (.ZN(n2210), 
	.C2(n1938), 
	.C1(n1474), 
	.B2(n1473), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1472));
   INV_X1 U3624 (.ZN(n1474), 
	.A(n4507));
   INV_X1 U3625 (.ZN(n1473), 
	.A(n4443));
   INV_X1 U3626 (.ZN(n1472), 
	.A(n4539));
   AOI222_X1 U3628 (.ZN(n5501), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[17] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n437), 
	.A2(n5564), 
	.A1(n6152));
   NAND2_X1 U3629 (.ZN(n437), 
	.A2(n2225), 
	.A1(n2224));
   AOI222_X1 U3630 (.ZN(n2225), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [17]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [17]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [17]));
   AOI22_X1 U3631 (.ZN(n2224), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [17]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [17]));
   NAND3_X1 U3632 (.ZN(n6152), 
	.A3(n2228), 
	.A2(n2227), 
	.A1(n2226));
   AOI222_X1 U3633 (.ZN(n2228), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[17] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[17] ), 
	.A2(n2229), 
	.A1(n1208));
   INV_X1 U3634 (.ZN(n2229), 
	.A(\UUT/Mpath/the_alu/N49 ));
   AOI22_X1 U3635 (.ZN(n2227), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N108 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N140 ));
   AOI22_X1 U3636 (.ZN(n2226), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N204 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N172 ));
   INV_X1 U3637 (.ZN(n2223), 
	.A(n431));
   NAND4_X1 U3638 (.ZN(n431), 
	.A4(n2233), 
	.A3(n2232), 
	.A2(n2231), 
	.A1(n2230));
   NOR4_X1 U3639 (.ZN(n2233), 
	.A4(n2237), 
	.A3(n2236), 
	.A2(n2235), 
	.A1(n2234));
   NAND3_X1 U3640 (.ZN(n2237), 
	.A3(n6151), 
	.A2(n6149), 
	.A1(n6150));
   OAI211_X1 U3641 (.ZN(n2236), 
	.C2(n5404), 
	.C1(n5560), 
	.B(n6148), 
	.A(n6147));
   OAI222_X1 U3642 (.ZN(n2235), 
	.C2(n5372), 
	.C1(n5561), 
	.B2(n5244), 
	.B1(n5559), 
	.A2(n5276), 
	.A1(n5558));
   OAI221_X1 U3643 (.ZN(n2234), 
	.C2(n5212), 
	.C1(n5532), 
	.B2(n5180), 
	.B1(n5531), 
	.A(n2238));
   AOI22_X1 U3644 (.ZN(n2238), 
	.B2(n1926), 
	.B1(n1445), 
	.A2(n1925), 
	.A1(n1444));
   INV_X1 U3645 (.ZN(n1445), 
	.A(n4988));
   INV_X1 U3646 (.ZN(n1444), 
	.A(n4956));
   AOI211_X1 U3647 (.ZN(n2232), 
	.C2(n1927), 
	.C1(n1446), 
	.B(n2240), 
	.A(n2239));
   OAI22_X1 U3648 (.ZN(n2240), 
	.B2(n4732), 
	.B1(n5551), 
	.A2(n4828), 
	.A1(n5541));
   OAI222_X1 U3649 (.ZN(n2239), 
	.C2(n4700), 
	.C1(n5547), 
	.B2(n4636), 
	.B1(n5552), 
	.A2(n4668), 
	.A1(n5546));
   INV_X1 U3650 (.ZN(n1446), 
	.A(n4860));
   AOI221_X1 U3651 (.ZN(n2231), 
	.C2(n2241), 
	.C1(n1931), 
	.B2(n1450), 
	.B1(n1930), 
	.A(n2242));
   OAI22_X1 U3652 (.ZN(n2242), 
	.B2(n6373), 
	.B1(n5084), 
	.A2(n1934), 
	.A1(n4476));
   INV_X1 U3653 (.ZN(n2241), 
	.A(n5308));
   INV_X1 U3654 (.ZN(n1450), 
	.A(n5340));
   AOI222_X1 U3655 (.ZN(n2230), 
	.C2(n1938), 
	.C1(n1454), 
	.B2(n1453), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1452));
   INV_X1 U3656 (.ZN(n1454), 
	.A(n4508));
   INV_X1 U3657 (.ZN(n1453), 
	.A(n4444));
   INV_X1 U3658 (.ZN(n1452), 
	.A(n4540));
   AOI222_X1 U3660 (.ZN(n5504), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[16] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n464), 
	.A2(n5564), 
	.A1(n6161));
   NAND2_X1 U3661 (.ZN(n464), 
	.A2(n2245), 
	.A1(n2244));
   AOI222_X1 U3662 (.ZN(n2245), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [16]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [16]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [16]));
   AOI22_X1 U3663 (.ZN(n2244), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [16]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [16]));
   NAND3_X1 U3664 (.ZN(n6161), 
	.A3(n2248), 
	.A2(n2247), 
	.A1(n2246));
   AOI222_X1 U3665 (.ZN(n2248), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[16] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[16] ), 
	.A2(n2249), 
	.A1(n1208));
   INV_X1 U3666 (.ZN(n2249), 
	.A(\UUT/Mpath/the_alu/N51 ));
   AOI22_X1 U3667 (.ZN(n2247), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N109 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N141 ));
   AOI22_X1 U3668 (.ZN(n2246), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N205 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N173 ));
   INV_X1 U3669 (.ZN(n2243), 
	.A(n458));
   NAND4_X1 U3670 (.ZN(n458), 
	.A4(FE_OFN50_n2253), 
	.A3(n2252), 
	.A2(n2251), 
	.A1(n2250));
   NOR4_X1 U3671 (.ZN(n2253), 
	.A4(n2257), 
	.A3(n2256), 
	.A2(n2255), 
	.A1(n2254));
   NAND3_X1 U3672 (.ZN(n2257), 
	.A3(n6160), 
	.A2(n6158), 
	.A1(n6159));
   OAI211_X1 U3673 (.ZN(n2256), 
	.C2(n5405), 
	.C1(n5560), 
	.B(n6157), 
	.A(n6156));
   OAI222_X1 U3674 (.ZN(n2255), 
	.C2(n5373), 
	.C1(n5561), 
	.B2(n5245), 
	.B1(n5559), 
	.A2(n5277), 
	.A1(n5558));
   OAI221_X1 U3675 (.ZN(n2254), 
	.C2(n5213), 
	.C1(n5532), 
	.B2(n5181), 
	.B1(n5531), 
	.A(n2258));
   AOI22_X1 U3676 (.ZN(n2258), 
	.B2(n1926), 
	.B1(n1425), 
	.A2(n1925), 
	.A1(n1424));
   INV_X1 U3677 (.ZN(n1425), 
	.A(n4989));
   INV_X1 U3678 (.ZN(n1424), 
	.A(n4957));
   AOI211_X1 U3679 (.ZN(n2252), 
	.C2(n1927), 
	.C1(n1426), 
	.B(n2260), 
	.A(n2259));
   OAI22_X1 U3680 (.ZN(n2260), 
	.B2(n4733), 
	.B1(n5551), 
	.A2(n4829), 
	.A1(n5541));
   OAI222_X1 U3681 (.ZN(n2259), 
	.C2(n4701), 
	.C1(n5547), 
	.B2(n4637), 
	.B1(n5552), 
	.A2(n4669), 
	.A1(n5546));
   INV_X1 U3682 (.ZN(n1426), 
	.A(n4861));
   AOI221_X1 U3683 (.ZN(n2251), 
	.C2(n2261), 
	.C1(n1931), 
	.B2(n1430), 
	.B1(n1930), 
	.A(n2262));
   OAI22_X1 U3684 (.ZN(n2262), 
	.B2(n6373), 
	.B1(n5085), 
	.A2(n1934), 
	.A1(n4477));
   INV_X1 U3685 (.ZN(n2261), 
	.A(n5309));
   INV_X1 U3686 (.ZN(n1430), 
	.A(n5341));
   AOI222_X1 U3687 (.ZN(n2250), 
	.C2(n1938), 
	.C1(n1434), 
	.B2(n1433), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1432));
   INV_X1 U3688 (.ZN(n1434), 
	.A(n4509));
   INV_X1 U3689 (.ZN(n1433), 
	.A(n4445));
   INV_X1 U3690 (.ZN(n1432), 
	.A(n4541));
   AOI222_X1 U3692 (.ZN(n5507), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[15] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n493), 
	.A2(n5564), 
	.A1(n6169));
   NAND2_X1 U3693 (.ZN(n493), 
	.A2(n2265), 
	.A1(n2264));
   AOI222_X1 U3694 (.ZN(n2265), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [15]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [15]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [15]));
   AOI22_X1 U3695 (.ZN(n2264), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [15]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [15]));
   NAND3_X1 U3696 (.ZN(n6169), 
	.A3(n2268), 
	.A2(n2267), 
	.A1(n2266));
   AOI222_X1 U3697 (.ZN(n2268), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[15] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[15] ), 
	.A2(n2269), 
	.A1(n1208));
   INV_X1 U3698 (.ZN(n2269), 
	.A(\UUT/Mpath/the_alu/N53 ));
   AOI22_X1 U3699 (.ZN(n2267), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N110 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N142 ));
   AOI22_X1 U3700 (.ZN(n2266), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N206 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N174 ));
   INV_X1 U3701 (.ZN(n2263), 
	.A(n479));
   NAND4_X1 U3702 (.ZN(n479), 
	.A4(n2273), 
	.A3(n2272), 
	.A2(n2271), 
	.A1(n2270));
   NOR4_X1 U3703 (.ZN(n2273), 
	.A4(n2277), 
	.A3(n2276), 
	.A2(n2275), 
	.A1(n2274));
   NAND3_X1 U3704 (.ZN(n2277), 
	.A3(n6168), 
	.A2(n6166), 
	.A1(n6167));
   OAI211_X1 U3705 (.ZN(n2276), 
	.C2(n5406), 
	.C1(n5560), 
	.B(n6165), 
	.A(n6164));
   OAI222_X1 U3706 (.ZN(n2275), 
	.C2(n5374), 
	.C1(n5561), 
	.B2(n5246), 
	.B1(n5559), 
	.A2(n5278), 
	.A1(n5558));
   OAI221_X1 U3707 (.ZN(n2274), 
	.C2(n5214), 
	.C1(n5532), 
	.B2(n5182), 
	.B1(n5531), 
	.A(n2278));
   AOI22_X1 U3708 (.ZN(n2278), 
	.B2(n1926), 
	.B1(n1405), 
	.A2(n1925), 
	.A1(n1404));
   INV_X1 U3709 (.ZN(n1405), 
	.A(n4990));
   INV_X1 U3710 (.ZN(n1404), 
	.A(n4958));
   AOI211_X1 U3711 (.ZN(n2272), 
	.C2(n1927), 
	.C1(n1406), 
	.B(n2280), 
	.A(n2279));
   OAI22_X1 U3712 (.ZN(n2280), 
	.B2(n4734), 
	.B1(n5551), 
	.A2(n4830), 
	.A1(n5541));
   OAI222_X1 U3713 (.ZN(n2279), 
	.C2(n4702), 
	.C1(n5547), 
	.B2(n4638), 
	.B1(n5552), 
	.A2(n4670), 
	.A1(n5546));
   INV_X1 U3714 (.ZN(n1406), 
	.A(n4862));
   AOI221_X1 U3715 (.ZN(n2271), 
	.C2(n2281), 
	.C1(n1931), 
	.B2(n1410), 
	.B1(n1930), 
	.A(n2282));
   OAI22_X1 U3716 (.ZN(n2282), 
	.B2(n6373), 
	.B1(n5086), 
	.A2(n1934), 
	.A1(n4478));
   INV_X1 U3717 (.ZN(n2281), 
	.A(n5310));
   INV_X1 U3718 (.ZN(n1410), 
	.A(n5342));
   AOI222_X1 U3719 (.ZN(n2270), 
	.C2(n1938), 
	.C1(n1414), 
	.B2(n1413), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1412));
   INV_X1 U3720 (.ZN(n1414), 
	.A(n4510));
   INV_X1 U3721 (.ZN(n1413), 
	.A(n4446));
   INV_X1 U3722 (.ZN(n1412), 
	.A(n4542));
   AOI222_X1 U3724 (.ZN(n5510), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[14] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n518), 
	.A2(n5564), 
	.A1(n6180));
   NAND2_X1 U3725 (.ZN(n518), 
	.A2(n2285), 
	.A1(n2284));
   AOI222_X1 U3726 (.ZN(n2285), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [14]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [14]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [14]));
   AOI22_X1 U3727 (.ZN(n2284), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [14]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [14]));
   NAND3_X1 U3728 (.ZN(n6180), 
	.A3(n2288), 
	.A2(n2287), 
	.A1(n2286));
   AOI222_X1 U3729 (.ZN(n2288), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[14] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[14] ), 
	.A2(n2289), 
	.A1(n1208));
   INV_X1 U3730 (.ZN(n2289), 
	.A(\UUT/Mpath/the_alu/N55 ));
   AOI22_X1 U3731 (.ZN(n2287), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N111 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N143 ));
   AOI22_X1 U3732 (.ZN(n2286), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N207 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N175 ));
   INV_X1 U3733 (.ZN(n2283), 
	.A(n508));
   NAND4_X1 U3734 (.ZN(n508), 
	.A4(FE_OFN54_n2293), 
	.A3(n2292), 
	.A2(n2291), 
	.A1(n2290));
   NOR4_X1 U3735 (.ZN(n2293), 
	.A4(n2297), 
	.A3(n2296), 
	.A2(n2295), 
	.A1(n2294));
   NAND3_X1 U3736 (.ZN(n2297), 
	.A3(n6179), 
	.A2(n6177), 
	.A1(n6178));
   OAI211_X1 U3737 (.ZN(n2296), 
	.C2(n5407), 
	.C1(n5560), 
	.B(n6176), 
	.A(n6175));
   OAI222_X1 U3738 (.ZN(n2295), 
	.C2(n5375), 
	.C1(n5561), 
	.B2(n5247), 
	.B1(n5559), 
	.A2(n5279), 
	.A1(n5558));
   OAI221_X1 U3739 (.ZN(n2294), 
	.C2(n5215), 
	.C1(n5532), 
	.B2(n5183), 
	.B1(n5531), 
	.A(n2298));
   AOI22_X1 U3740 (.ZN(n2298), 
	.B2(n1926), 
	.B1(n1385), 
	.A2(n1925), 
	.A1(n1384));
   INV_X1 U3741 (.ZN(n1385), 
	.A(n4991));
   INV_X1 U3742 (.ZN(n1384), 
	.A(n4959));
   AOI211_X1 U3743 (.ZN(n2292), 
	.C2(n1927), 
	.C1(n1386), 
	.B(n2300), 
	.A(n2299));
   OAI22_X1 U3744 (.ZN(n2300), 
	.B2(n4735), 
	.B1(n5551), 
	.A2(n4831), 
	.A1(n5541));
   OAI222_X1 U3745 (.ZN(n2299), 
	.C2(n4703), 
	.C1(n5547), 
	.B2(n4639), 
	.B1(n5552), 
	.A2(n4671), 
	.A1(n5546));
   INV_X1 U3746 (.ZN(n1386), 
	.A(n4863));
   AOI221_X1 U3747 (.ZN(n2291), 
	.C2(n2301), 
	.C1(n1931), 
	.B2(n1390), 
	.B1(n1930), 
	.A(n2302));
   OAI22_X1 U3748 (.ZN(n2302), 
	.B2(n6373), 
	.B1(n5087), 
	.A2(n1934), 
	.A1(n4479));
   INV_X1 U3749 (.ZN(n2301), 
	.A(n5311));
   INV_X1 U3750 (.ZN(n1390), 
	.A(n5343));
   AOI222_X1 U3751 (.ZN(n2290), 
	.C2(n1938), 
	.C1(n1394), 
	.B2(n1393), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1392));
   INV_X1 U3752 (.ZN(n1394), 
	.A(n4511));
   INV_X1 U3753 (.ZN(n1393), 
	.A(n4447));
   INV_X1 U3754 (.ZN(n1392), 
	.A(n4543));
   AOI222_X1 U3756 (.ZN(n5513), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[13] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n543), 
	.A2(n5564), 
	.A1(n6187));
   NAND2_X1 U3757 (.ZN(n543), 
	.A2(n2305), 
	.A1(n2304));
   AOI222_X1 U3758 (.ZN(n2305), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [13]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [13]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [13]));
   AOI22_X1 U3759 (.ZN(n2304), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [13]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [13]));
   NAND3_X1 U3760 (.ZN(n6187), 
	.A3(n2308), 
	.A2(n2307), 
	.A1(n2306));
   AOI222_X1 U3761 (.ZN(n2308), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[13] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[13] ), 
	.A2(n2309), 
	.A1(n1208));
   INV_X1 U3762 (.ZN(n2309), 
	.A(\UUT/Mpath/the_alu/N57 ));
   AOI22_X1 U3763 (.ZN(n2307), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N112 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N144 ));
   AOI22_X1 U3764 (.ZN(n2306), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N208 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N176 ));
   INV_X1 U3765 (.ZN(n2303), 
	.A(n533));
   NAND4_X1 U3766 (.ZN(n533), 
	.A4(FE_OFN57_n2313), 
	.A3(n2312), 
	.A2(n2311), 
	.A1(n2310));
   NOR4_X1 U3767 (.ZN(n2313), 
	.A4(n2317), 
	.A3(n2316), 
	.A2(n2315), 
	.A1(n2314));
   NAND3_X1 U3768 (.ZN(n2317), 
	.A3(n6186), 
	.A2(n6184), 
	.A1(n6185));
   OAI211_X1 U3769 (.ZN(n2316), 
	.C2(n5408), 
	.C1(n5560), 
	.B(n6183), 
	.A(n6182));
   OAI222_X1 U3770 (.ZN(n2315), 
	.C2(n5376), 
	.C1(n5561), 
	.B2(n5248), 
	.B1(n5559), 
	.A2(n5280), 
	.A1(n5558));
   OAI221_X1 U3771 (.ZN(n2314), 
	.C2(n5216), 
	.C1(n5532), 
	.B2(n5184), 
	.B1(n5531), 
	.A(n2318));
   AOI22_X1 U3772 (.ZN(n2318), 
	.B2(n1926), 
	.B1(n1365), 
	.A2(n1925), 
	.A1(n1364));
   INV_X1 U3773 (.ZN(n1365), 
	.A(n4992));
   INV_X1 U3774 (.ZN(n1364), 
	.A(n4960));
   AOI211_X1 U3775 (.ZN(n2312), 
	.C2(n1927), 
	.C1(n1366), 
	.B(n2320), 
	.A(n2319));
   OAI22_X1 U3776 (.ZN(n2320), 
	.B2(n4736), 
	.B1(n5551), 
	.A2(n4832), 
	.A1(n5541));
   OAI222_X1 U3777 (.ZN(n2319), 
	.C2(n4704), 
	.C1(n5547), 
	.B2(n4640), 
	.B1(n5552), 
	.A2(n4672), 
	.A1(n5546));
   INV_X1 U3778 (.ZN(n1366), 
	.A(n4864));
   AOI221_X1 U3779 (.ZN(n2311), 
	.C2(n2321), 
	.C1(n1931), 
	.B2(n1370), 
	.B1(n1930), 
	.A(n2322));
   OAI22_X1 U3780 (.ZN(n2322), 
	.B2(n6373), 
	.B1(n5088), 
	.A2(n1934), 
	.A1(n4480));
   INV_X1 U3781 (.ZN(n2321), 
	.A(n5312));
   INV_X1 U3782 (.ZN(n1370), 
	.A(n5344));
   AOI222_X1 U3783 (.ZN(n2310), 
	.C2(n1938), 
	.C1(n1374), 
	.B2(n1373), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1372));
   INV_X1 U3784 (.ZN(n1374), 
	.A(n4512));
   INV_X1 U3785 (.ZN(n1373), 
	.A(n4448));
   INV_X1 U3786 (.ZN(n1372), 
	.A(n4544));
   NAND2_X1 U3787 (.ZN(\UUT/Mcontrol/st_logic/N42 ), 
	.A2(n2323), 
	.A1(\UUT/Mcontrol/bp_logicB/memory_main ));
   INV_X1 U3788 (.ZN(n2323), 
	.A(\UUT/Mcontrol/bp_logicB/exec_main ));
   INV_X1 U3793 (.ZN(\UUT/break_code[2] ), 
	.A(FE_OFN196_n764));
   AOI222_X1 U3796 (.ZN(n5459), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[2] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n785), 
	.A2(n5564), 
	.A1(n6202));
   NAND2_X1 U3797 (.ZN(n785), 
	.A2(n2332), 
	.A1(n2331));
   AOI222_X1 U3798 (.ZN(n2332), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [2]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [2]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [2]));
   AOI22_X1 U3799 (.ZN(n2331), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [2]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [2]));
   NAND3_X1 U3800 (.ZN(n6202), 
	.A3(n2335), 
	.A2(n2334), 
	.A1(n2333));
   AOI222_X1 U3801 (.ZN(n2335), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[2] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[2] ), 
	.A2(n2336), 
	.A1(n1208));
   INV_X1 U3802 (.ZN(n2336), 
	.A(\UUT/Mpath/the_alu/N79 ));
   AOI22_X1 U3803 (.ZN(n2334), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N123 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N155 ));
   AOI22_X1 U3804 (.ZN(n2333), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N219 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N187 ));
   INV_X1 U3805 (.ZN(n2330), 
	.A(n776));
   NAND4_X1 U3806 (.ZN(n776), 
	.A4(FE_OFN83_n2340), 
	.A3(n2339), 
	.A2(n2338), 
	.A1(n2337));
   NOR4_X1 U3807 (.ZN(n2340), 
	.A4(n2344), 
	.A3(n2343), 
	.A2(n2342), 
	.A1(n2341));
   NAND3_X1 U3808 (.ZN(n2344), 
	.A3(n6262), 
	.A2(n6260), 
	.A1(n6261));
   OAI211_X1 U3809 (.ZN(n2343), 
	.C2(n5390), 
	.C1(n5560), 
	.B(n6259), 
	.A(n6258));
   OAI222_X1 U3810 (.ZN(n2342), 
	.C2(n5358), 
	.C1(n5561), 
	.B2(n5230), 
	.B1(n5559), 
	.A2(n5262), 
	.A1(n5558));
   OAI221_X1 U3811 (.ZN(n2341), 
	.C2(n5198), 
	.C1(n5532), 
	.B2(n5166), 
	.B1(n5531), 
	.A(n2345));
   AOI22_X1 U3812 (.ZN(n2345), 
	.B2(n1926), 
	.B1(n1725), 
	.A2(n1925), 
	.A1(n1724));
   INV_X1 U3813 (.ZN(n1725), 
	.A(n4974));
   INV_X1 U3814 (.ZN(n1724), 
	.A(n4942));
   AOI211_X1 U3815 (.ZN(n2339), 
	.C2(n1927), 
	.C1(n1726), 
	.B(n2347), 
	.A(n2346));
   OAI22_X1 U3816 (.ZN(n2347), 
	.B2(n4718), 
	.B1(n5551), 
	.A2(n4814), 
	.A1(n5541));
   OAI222_X1 U3817 (.ZN(n2346), 
	.C2(n4686), 
	.C1(n5547), 
	.B2(n4622), 
	.B1(n5552), 
	.A2(n4654), 
	.A1(n5546));
   INV_X1 U3818 (.ZN(n1726), 
	.A(n4846));
   AOI221_X1 U3819 (.ZN(n2338), 
	.C2(n2348), 
	.C1(n1931), 
	.B2(n1730), 
	.B1(n1930), 
	.A(n2349));
   OAI22_X1 U3820 (.ZN(n2349), 
	.B2(n6373), 
	.B1(n5070), 
	.A2(n1934), 
	.A1(n4462));
   INV_X1 U3821 (.ZN(n2348), 
	.A(n5294));
   INV_X1 U3822 (.ZN(n1730), 
	.A(n5326));
   AOI222_X1 U3823 (.ZN(n2337), 
	.C2(n1938), 
	.C1(n1734), 
	.B2(n1733), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1732));
   INV_X1 U3824 (.ZN(n1734), 
	.A(n4494));
   INV_X1 U3825 (.ZN(n1733), 
	.A(n4430));
   INV_X1 U3826 (.ZN(n1732), 
	.A(n4526));
   AOI22_X1 U3830 (.ZN(n2351), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [12]), 
	.B1(n6449), 
	.A2(\UUT/break_code[12] ), 
	.A1(n908));
   OAI21_X1 U3831 (.ZN(\UUT/break_code[12] ), 
	.B2(n2072), 
	.B1(n6035), 
	.A(n2352));
   NAND2_X1 U3832 (.ZN(n2352), 
	.A2(n2074), 
	.A1(n6272));
   INV_X1 U3833 (.ZN(n6035), 
	.A(\UUT/Mcontrol/d_sampled_finstr [12]));
   AOI222_X1 U3835 (.ZN(n5516), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[12] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n569), 
	.A2(n5564), 
	.A1(n6203));
   NAND2_X1 U3836 (.ZN(n569), 
	.A2(n2355), 
	.A1(n2354));
   AOI222_X1 U3837 (.ZN(n2355), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [12]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [12]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [12]));
   AOI22_X1 U3838 (.ZN(n2354), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [12]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [12]));
   NAND3_X1 U3839 (.ZN(n6203), 
	.A3(n2358), 
	.A2(n2357), 
	.A1(n2356));
   AOI222_X1 U3840 (.ZN(n2358), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[12] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[12] ), 
	.A2(n2359), 
	.A1(n1208));
   INV_X1 U3841 (.ZN(n2359), 
	.A(\UUT/Mpath/the_alu/N59 ));
   AOI22_X1 U3842 (.ZN(n2357), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N113 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N145 ));
   AOI22_X1 U3843 (.ZN(n2356), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N209 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N177 ));
   INV_X1 U3844 (.ZN(n2353), 
	.A(n559));
   NAND4_X1 U3845 (.ZN(n559), 
	.A4(FE_OFN60_n2363), 
	.A3(n2362), 
	.A2(n2361), 
	.A1(n2360));
   NOR4_X1 U3846 (.ZN(n2363), 
	.A4(n2367), 
	.A3(n2366), 
	.A2(n2365), 
	.A1(n2364));
   NAND3_X1 U3847 (.ZN(n2367), 
	.A3(n6271), 
	.A2(n6269), 
	.A1(n6270));
   OAI211_X1 U3848 (.ZN(n2366), 
	.C2(n5409), 
	.C1(n5560), 
	.B(n6268), 
	.A(n6267));
   OAI222_X1 U3849 (.ZN(n2365), 
	.C2(n5377), 
	.C1(n5561), 
	.B2(n5249), 
	.B1(n5559), 
	.A2(n5281), 
	.A1(n5558));
   OAI221_X1 U3850 (.ZN(n2364), 
	.C2(n5217), 
	.C1(n5532), 
	.B2(n5185), 
	.B1(n5531), 
	.A(n2368));
   AOI22_X1 U3851 (.ZN(n2368), 
	.B2(n1926), 
	.B1(n1345), 
	.A2(n1925), 
	.A1(n1344));
   INV_X1 U3852 (.ZN(n1345), 
	.A(n4993));
   INV_X1 U3853 (.ZN(n1344), 
	.A(n4961));
   AOI211_X1 U3854 (.ZN(n2362), 
	.C2(n1927), 
	.C1(n1346), 
	.B(n2370), 
	.A(n2369));
   OAI22_X1 U3855 (.ZN(n2370), 
	.B2(n4737), 
	.B1(n5551), 
	.A2(n4833), 
	.A1(n5541));
   OAI222_X1 U3856 (.ZN(n2369), 
	.C2(n4705), 
	.C1(n5547), 
	.B2(n4641), 
	.B1(n5552), 
	.A2(n4673), 
	.A1(n5546));
   INV_X1 U3857 (.ZN(n1346), 
	.A(n4865));
   AOI221_X1 U3858 (.ZN(n2361), 
	.C2(n2371), 
	.C1(n1931), 
	.B2(n1350), 
	.B1(n1930), 
	.A(n2372));
   OAI22_X1 U3859 (.ZN(n2372), 
	.B2(n6373), 
	.B1(n5089), 
	.A2(n1934), 
	.A1(n4481));
   INV_X1 U3860 (.ZN(n2371), 
	.A(n5313));
   INV_X1 U3861 (.ZN(n1350), 
	.A(n5345));
   AOI222_X1 U3862 (.ZN(n2360), 
	.C2(n1938), 
	.C1(n1354), 
	.B2(n1353), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1352));
   INV_X1 U3863 (.ZN(n1354), 
	.A(n4513));
   INV_X1 U3864 (.ZN(n1353), 
	.A(n4449));
   INV_X1 U3865 (.ZN(n1352), 
	.A(n4545));
   AOI22_X1 U3869 (.ZN(n2374), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [11]), 
	.B1(n6449), 
	.A2(\UUT/break_code[11] ), 
	.A1(n908));
   OAI21_X1 U3870 (.ZN(\UUT/break_code[11] ), 
	.B2(n2072), 
	.B1(n6036), 
	.A(n2375));
   NAND2_X1 U3871 (.ZN(n2375), 
	.A2(n2074), 
	.A1(n6278));
   INV_X1 U3872 (.ZN(n6036), 
	.A(\UUT/Mcontrol/d_sampled_finstr [11]));
   AOI222_X1 U3874 (.ZN(n5519), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[11] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n594), 
	.A2(n5564), 
	.A1(n6204));
   NAND2_X1 U3875 (.ZN(n594), 
	.A2(n2378), 
	.A1(n2377));
   AOI222_X1 U3876 (.ZN(n2378), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [11]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [11]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [11]));
   AOI22_X1 U3877 (.ZN(n2377), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [11]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [11]));
   NAND3_X1 U3878 (.ZN(n6204), 
	.A3(n2381), 
	.A2(n2380), 
	.A1(n2379));
   AOI222_X1 U3879 (.ZN(n2381), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[11] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[11] ), 
	.A2(n2382), 
	.A1(n1208));
   INV_X1 U3880 (.ZN(n2382), 
	.A(\UUT/Mpath/the_alu/N61 ));
   AOI22_X1 U3881 (.ZN(n2380), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N114 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N146 ));
   AOI22_X1 U3882 (.ZN(n2379), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N210 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N178 ));
   INV_X1 U3883 (.ZN(n2376), 
	.A(n584));
   NAND4_X1 U3884 (.ZN(n584), 
	.A4(FE_OFN63_n2386), 
	.A3(n2385), 
	.A2(n2384), 
	.A1(n2383));
   NOR4_X1 U3885 (.ZN(n2386), 
	.A4(n2390), 
	.A3(n2389), 
	.A2(n2388), 
	.A1(n2387));
   NAND3_X1 U3886 (.ZN(n2390), 
	.A3(n6277), 
	.A2(n6275), 
	.A1(n6276));
   OAI211_X1 U3887 (.ZN(n2389), 
	.C2(n5410), 
	.C1(n5560), 
	.B(n6274), 
	.A(n6273));
   OAI222_X1 U3888 (.ZN(n2388), 
	.C2(n5378), 
	.C1(n5561), 
	.B2(n5250), 
	.B1(n5559), 
	.A2(n5282), 
	.A1(n5558));
   OAI221_X1 U3889 (.ZN(n2387), 
	.C2(n5218), 
	.C1(n5532), 
	.B2(n5186), 
	.B1(n5531), 
	.A(n2391));
   AOI22_X1 U3890 (.ZN(n2391), 
	.B2(n1926), 
	.B1(n1325), 
	.A2(n1925), 
	.A1(n1324));
   INV_X1 U3891 (.ZN(n1325), 
	.A(n4994));
   INV_X1 U3892 (.ZN(n1324), 
	.A(n4962));
   AOI211_X1 U3893 (.ZN(n2385), 
	.C2(n1927), 
	.C1(n1326), 
	.B(n2393), 
	.A(n2392));
   OAI22_X1 U3894 (.ZN(n2393), 
	.B2(n4738), 
	.B1(n5551), 
	.A2(n4834), 
	.A1(n5541));
   OAI222_X1 U3895 (.ZN(n2392), 
	.C2(n4706), 
	.C1(n5547), 
	.B2(n4642), 
	.B1(n5552), 
	.A2(n4674), 
	.A1(n5546));
   INV_X1 U3896 (.ZN(n1326), 
	.A(n4866));
   AOI221_X1 U3897 (.ZN(n2384), 
	.C2(n2394), 
	.C1(n1931), 
	.B2(n1330), 
	.B1(n1930), 
	.A(n2395));
   OAI22_X1 U3898 (.ZN(n2395), 
	.B2(n6373), 
	.B1(n5090), 
	.A2(n1934), 
	.A1(n4482));
   INV_X1 U3899 (.ZN(n2394), 
	.A(n5314));
   INV_X1 U3900 (.ZN(n1330), 
	.A(n5346));
   AOI222_X1 U3901 (.ZN(n2383), 
	.C2(n1938), 
	.C1(n1334), 
	.B2(n1333), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1332));
   INV_X1 U3902 (.ZN(n1334), 
	.A(n4514));
   INV_X1 U3903 (.ZN(n1333), 
	.A(n4450));
   INV_X1 U3904 (.ZN(n1332), 
	.A(n4546));
   INV_X1 U3905 (.ZN(\UUT/Mcontrol/Program_counter/N24 ), 
	.A(n979));
   OAI21_X1 U3909 (.ZN(\UUT/break_code[10] ), 
	.B2(n2072), 
	.B1(n5881), 
	.A(n2398));
   NAND2_X1 U3910 (.ZN(n2398), 
	.A2(n2074), 
	.A1(n6327));
   INV_X1 U3911 (.ZN(n5881), 
	.A(\UUT/Mcontrol/d_sampled_finstr [10]));
   AOI222_X1 U3913 (.ZN(n5522), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[10] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n1162), 
	.A2(n5564), 
	.A1(n6205));
   NAND2_X1 U3914 (.ZN(n1162), 
	.A2(n2401), 
	.A1(n2400));
   AOI222_X1 U3915 (.ZN(n2401), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [10]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [10]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [10]));
   AOI22_X1 U3916 (.ZN(n2400), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [10]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [10]));
   NAND3_X1 U3917 (.ZN(n6205), 
	.A3(n2404), 
	.A2(n2403), 
	.A1(n2402));
   AOI222_X1 U3918 (.ZN(n2404), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[10] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[10] ), 
	.A2(n2405), 
	.A1(n1208));
   INV_X1 U3919 (.ZN(n2405), 
	.A(\UUT/Mpath/the_alu/N63 ));
   AOI22_X1 U3920 (.ZN(n2403), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N115 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N147 ));
   AOI22_X1 U3921 (.ZN(n2402), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N211 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N179 ));
   INV_X1 U3922 (.ZN(n2399), 
	.A(n604));
   NAND4_X1 U3923 (.ZN(n604), 
	.A4(FE_OFN95_n2409), 
	.A3(n2408), 
	.A2(n2407), 
	.A1(n2406));
   NOR4_X1 U3924 (.ZN(n2409), 
	.A4(n2413), 
	.A3(n2412), 
	.A2(n2411), 
	.A1(n2410));
   NAND3_X1 U3925 (.ZN(n2413), 
	.A3(n6283), 
	.A2(n6281), 
	.A1(n6282));
   OAI211_X1 U3926 (.ZN(n2412), 
	.C2(n5411), 
	.C1(n5560), 
	.B(n6280), 
	.A(n6279));
   OAI222_X1 U3927 (.ZN(n2411), 
	.C2(n5379), 
	.C1(n5561), 
	.B2(n5251), 
	.B1(n5559), 
	.A2(n5283), 
	.A1(n5558));
   OAI221_X1 U3928 (.ZN(n2410), 
	.C2(n5219), 
	.C1(n5532), 
	.B2(n5187), 
	.B1(n5531), 
	.A(n2414));
   AOI22_X1 U3929 (.ZN(n2414), 
	.B2(n1926), 
	.B1(n1305), 
	.A2(n1925), 
	.A1(n1304));
   INV_X1 U3930 (.ZN(n1305), 
	.A(n4995));
   INV_X1 U3931 (.ZN(n1304), 
	.A(n4963));
   AOI211_X1 U3932 (.ZN(n2408), 
	.C2(n1927), 
	.C1(n1306), 
	.B(n2416), 
	.A(n2415));
   OAI22_X1 U3933 (.ZN(n2416), 
	.B2(n4739), 
	.B1(n5551), 
	.A2(n4835), 
	.A1(n5541));
   OAI222_X1 U3934 (.ZN(n2415), 
	.C2(n4707), 
	.C1(n5547), 
	.B2(n4643), 
	.B1(n5552), 
	.A2(n4675), 
	.A1(n5546));
   INV_X1 U3935 (.ZN(n1306), 
	.A(n4867));
   AOI221_X1 U3936 (.ZN(n2407), 
	.C2(n2417), 
	.C1(n1931), 
	.B2(n1310), 
	.B1(n1930), 
	.A(n2418));
   OAI22_X1 U3937 (.ZN(n2418), 
	.B2(n6373), 
	.B1(n5091), 
	.A2(n1934), 
	.A1(n4483));
   INV_X1 U3938 (.ZN(n2417), 
	.A(n5315));
   INV_X1 U3939 (.ZN(n1310), 
	.A(n5347));
   AOI222_X1 U3940 (.ZN(n2406), 
	.C2(n1938), 
	.C1(n1314), 
	.B2(n1313), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1312));
   INV_X1 U3941 (.ZN(n1314), 
	.A(n4515));
   INV_X1 U3942 (.ZN(n1313), 
	.A(n4451));
   INV_X1 U3943 (.ZN(n1312), 
	.A(n4547));
   INV_X1 U3944 (.ZN(\UUT/Mcontrol/Program_counter/N22 ), 
	.A(n909));
   OAI21_X1 U3948 (.ZN(\UUT/break_code[9] ), 
	.B2(n2072), 
	.B1(n5889), 
	.A(n2421));
   NAND2_X1 U3949 (.ZN(n2421), 
	.A2(n2074), 
	.A1(n6216));
   INV_X1 U3950 (.ZN(n5889), 
	.A(\UUT/Mcontrol/d_sampled_finstr [9]));
   OAI222_X1 U3951 (.ZN(\UUT/branch_rega [9]), 
	.C2(FE_OFN194_n5429), 
	.C1(n5528), 
	.B2(n2422), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5433));
   AOI222_X1 U3952 (.ZN(n5429), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[9] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n629), 
	.A2(n5564), 
	.A1(n6189));
   NAND2_X1 U3953 (.ZN(n629), 
	.A2(n2424), 
	.A1(n2423));
   AOI222_X1 U3954 (.ZN(n2424), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [9]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [9]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [9]));
   AOI22_X1 U3955 (.ZN(n2423), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [9]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [9]));
   NAND3_X1 U3956 (.ZN(n6189), 
	.A3(n2427), 
	.A2(n2426), 
	.A1(n2425));
   AOI222_X1 U3957 (.ZN(n2427), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[9] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[9] ), 
	.A2(n2428), 
	.A1(n1208));
   INV_X1 U3958 (.ZN(n2428), 
	.A(\UUT/Mpath/the_alu/N65 ));
   AOI22_X1 U3959 (.ZN(n2426), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N116 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N148 ));
   AOI22_X1 U3960 (.ZN(n2425), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N212 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N180 ));
   INV_X1 U3961 (.ZN(n2422), 
	.A(n619));
   NAND4_X1 U3962 (.ZN(n619), 
	.A4(n2432), 
	.A3(n2431), 
	.A2(n2430), 
	.A1(n2429));
   NOR4_X1 U3963 (.ZN(n2432), 
	.A4(n2436), 
	.A3(n2435), 
	.A2(n2434), 
	.A1(n2433));
   NAND3_X1 U3964 (.ZN(n2436), 
	.A3(n6215), 
	.A2(n6213), 
	.A1(n6214));
   OAI211_X1 U3965 (.ZN(n2435), 
	.C2(n5381), 
	.C1(n5560), 
	.B(n6212), 
	.A(n6211));
   OAI222_X1 U3966 (.ZN(n2434), 
	.C2(n5349), 
	.C1(n5561), 
	.B2(n5221), 
	.B1(n5559), 
	.A2(n5253), 
	.A1(n5558));
   OAI221_X1 U3967 (.ZN(n2433), 
	.C2(n5189), 
	.C1(n5532), 
	.B2(n5157), 
	.B1(n5531), 
	.A(n2437));
   AOI22_X1 U3968 (.ZN(n2437), 
	.B2(n1926), 
	.B1(n1905), 
	.A2(n1925), 
	.A1(n1904));
   INV_X1 U3969 (.ZN(n1905), 
	.A(n4965));
   INV_X1 U3970 (.ZN(n1904), 
	.A(n4933));
   AOI211_X1 U3971 (.ZN(n2431), 
	.C2(n1927), 
	.C1(n1906), 
	.B(n2439), 
	.A(n2438));
   OAI22_X1 U3972 (.ZN(n2439), 
	.B2(n4709), 
	.B1(n5551), 
	.A2(n4805), 
	.A1(n5541));
   OAI222_X1 U3973 (.ZN(n2438), 
	.C2(n4677), 
	.C1(n5547), 
	.B2(n4613), 
	.B1(n5552), 
	.A2(n4645), 
	.A1(n5546));
   INV_X1 U3974 (.ZN(n1906), 
	.A(n4837));
   AOI221_X1 U3975 (.ZN(n2430), 
	.C2(n2440), 
	.C1(n1931), 
	.B2(n1910), 
	.B1(n1930), 
	.A(n2441));
   OAI22_X1 U3976 (.ZN(n2441), 
	.B2(n6373), 
	.B1(n5061), 
	.A2(n1934), 
	.A1(n4453));
   INV_X1 U3977 (.ZN(n2440), 
	.A(n5285));
   INV_X1 U3978 (.ZN(n1910), 
	.A(n5317));
   AOI222_X1 U3979 (.ZN(n2429), 
	.C2(n1938), 
	.C1(n1915), 
	.B2(n1914), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1913));
   INV_X1 U3980 (.ZN(n1915), 
	.A(n4485));
   INV_X1 U3981 (.ZN(n1914), 
	.A(n4421));
   INV_X1 U3982 (.ZN(n1913), 
	.A(n4517));
   AOI22_X1 U3986 (.ZN(n2443), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [8]), 
	.B1(n906), 
	.A2(\UUT/break_code[8] ), 
	.A1(n908));
   OAI21_X1 U3987 (.ZN(\UUT/break_code[8] ), 
	.B2(n2072), 
	.B1(n5897), 
	.A(n2444));
   NAND2_X1 U3988 (.ZN(n2444), 
	.A2(n2074), 
	.A1(n6222));
   INV_X1 U3989 (.ZN(n5897), 
	.A(\UUT/Mcontrol/d_sampled_finstr [8]));
   AOI222_X1 U3991 (.ZN(n5435), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[8] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n1153), 
	.A2(n5564), 
	.A1(n6190));
   NAND2_X1 U3992 (.ZN(n1153), 
	.A2(n2447), 
	.A1(n2446));
   AOI222_X1 U3993 (.ZN(n2447), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [8]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [8]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [8]));
   AOI22_X1 U3994 (.ZN(n2446), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [8]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [8]));
   NAND3_X1 U3995 (.ZN(n6190), 
	.A3(n2450), 
	.A2(n2449), 
	.A1(n2448));
   AOI222_X1 U3996 (.ZN(n2450), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[8] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[8] ), 
	.A2(n2451), 
	.A1(n1208));
   INV_X1 U3997 (.ZN(n2451), 
	.A(\UUT/Mpath/the_alu/N67 ));
   AOI22_X1 U3998 (.ZN(n2449), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N117 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N149 ));
   AOI22_X1 U3999 (.ZN(n2448), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N213 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N181 ));
   INV_X1 U4000 (.ZN(n2445), 
	.A(n640));
   NAND4_X1 U4001 (.ZN(n640), 
	.A4(FE_OFN94_n2455), 
	.A3(n2454), 
	.A2(n2453), 
	.A1(n2452));
   NOR4_X1 U4002 (.ZN(n2455), 
	.A4(n2459), 
	.A3(n2458), 
	.A2(n2457), 
	.A1(n2456));
   NAND3_X1 U4003 (.ZN(n2459), 
	.A3(n6221), 
	.A2(n6219), 
	.A1(n6220));
   OAI211_X1 U4004 (.ZN(n2458), 
	.C2(n5382), 
	.C1(n5560), 
	.B(n6218), 
	.A(n6217));
   OAI222_X1 U4005 (.ZN(n2457), 
	.C2(n5350), 
	.C1(n5561), 
	.B2(n5222), 
	.B1(n5559), 
	.A2(n5254), 
	.A1(n5558));
   OAI221_X1 U4006 (.ZN(n2456), 
	.C2(n5190), 
	.C1(n5532), 
	.B2(n5158), 
	.B1(n5531), 
	.A(n2460));
   AOI22_X1 U4007 (.ZN(n2460), 
	.B2(n1926), 
	.B1(n1885), 
	.A2(n1925), 
	.A1(n1884));
   INV_X1 U4008 (.ZN(n1885), 
	.A(n4966));
   INV_X1 U4009 (.ZN(n1884), 
	.A(n4934));
   AOI211_X1 U4010 (.ZN(n2454), 
	.C2(n1927), 
	.C1(n1886), 
	.B(n2462), 
	.A(n2461));
   OAI22_X1 U4011 (.ZN(n2462), 
	.B2(n4710), 
	.B1(n5551), 
	.A2(n4806), 
	.A1(n5541));
   OAI222_X1 U4012 (.ZN(n2461), 
	.C2(n4678), 
	.C1(n5547), 
	.B2(n4614), 
	.B1(n5552), 
	.A2(n4646), 
	.A1(n5546));
   INV_X1 U4013 (.ZN(n1886), 
	.A(n4838));
   AOI221_X1 U4014 (.ZN(n2453), 
	.C2(n2463), 
	.C1(n1931), 
	.B2(n1890), 
	.B1(n1930), 
	.A(n2464));
   OAI22_X1 U4015 (.ZN(n2464), 
	.B2(n6373), 
	.B1(n5062), 
	.A2(n1934), 
	.A1(n4454));
   INV_X1 U4016 (.ZN(n2463), 
	.A(n5286));
   INV_X1 U4017 (.ZN(n1890), 
	.A(n5318));
   AOI222_X1 U4018 (.ZN(n2452), 
	.C2(n1938), 
	.C1(n1894), 
	.B2(n1893), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1892));
   INV_X1 U4019 (.ZN(n1894), 
	.A(n4486));
   INV_X1 U4020 (.ZN(n1893), 
	.A(n4422));
   INV_X1 U4021 (.ZN(n1892), 
	.A(n4518));
   AOI22_X1 U4025 (.ZN(n2466), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [7]), 
	.B1(n906), 
	.A2(\UUT/break_code[7] ), 
	.A1(n908));
   OAI21_X1 U4026 (.ZN(\UUT/break_code[7] ), 
	.B2(n2072), 
	.B1(n6094), 
	.A(n2467));
   NAND2_X1 U4027 (.ZN(n2467), 
	.A2(n2074), 
	.A1(n6228));
   INV_X1 U4028 (.ZN(n6094), 
	.A(\UUT/Mcontrol/d_sampled_finstr [7]));
   AOI222_X1 U4030 (.ZN(n5438), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[7] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n664), 
	.A2(n5564), 
	.A1(n6191));
   NAND2_X1 U4031 (.ZN(n664), 
	.A2(n2470), 
	.A1(n2469));
   AOI222_X1 U4032 (.ZN(n2470), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [7]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [7]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [7]));
   AOI22_X1 U4033 (.ZN(n2469), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [7]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [7]));
   NAND3_X1 U4034 (.ZN(n6191), 
	.A3(n2473), 
	.A2(n2472), 
	.A1(n2471));
   AOI222_X1 U4035 (.ZN(n2473), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[7] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[7] ), 
	.A2(n2474), 
	.A1(n1208));
   INV_X1 U4036 (.ZN(n2474), 
	.A(\UUT/Mpath/the_alu/N69 ));
   AOI22_X1 U4037 (.ZN(n2472), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N118 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N150 ));
   AOI22_X1 U4038 (.ZN(n2471), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N214 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N182 ));
   INV_X1 U4039 (.ZN(n2468), 
	.A(n656));
   NAND4_X1 U4040 (.ZN(n656), 
	.A4(FE_OFN69_n2478), 
	.A3(n2477), 
	.A2(n2476), 
	.A1(n2475));
   NOR4_X1 U4041 (.ZN(n2478), 
	.A4(n2482), 
	.A3(n2481), 
	.A2(n2480), 
	.A1(n2479));
   NAND3_X1 U4042 (.ZN(n2482), 
	.A3(n6227), 
	.A2(n6225), 
	.A1(n6226));
   OAI211_X1 U4043 (.ZN(n2481), 
	.C2(n5383), 
	.C1(n5560), 
	.B(n6224), 
	.A(n6223));
   OAI222_X1 U4044 (.ZN(n2480), 
	.C2(n5351), 
	.C1(n5561), 
	.B2(n5223), 
	.B1(n5559), 
	.A2(n5255), 
	.A1(n5558));
   OAI221_X1 U4045 (.ZN(n2479), 
	.C2(n5191), 
	.C1(n5532), 
	.B2(n5159), 
	.B1(n5531), 
	.A(n2483));
   AOI22_X1 U4046 (.ZN(n2483), 
	.B2(n1926), 
	.B1(n1865), 
	.A2(n1925), 
	.A1(n1864));
   INV_X1 U4047 (.ZN(n1865), 
	.A(n4967));
   INV_X1 U4048 (.ZN(n1864), 
	.A(n4935));
   AOI211_X1 U4049 (.ZN(n2477), 
	.C2(n1927), 
	.C1(n1866), 
	.B(n2485), 
	.A(n2484));
   OAI22_X1 U4050 (.ZN(n2485), 
	.B2(n4711), 
	.B1(n5551), 
	.A2(n4807), 
	.A1(n5541));
   OAI222_X1 U4051 (.ZN(n2484), 
	.C2(n4679), 
	.C1(n5547), 
	.B2(n4615), 
	.B1(n5552), 
	.A2(n4647), 
	.A1(n5546));
   INV_X1 U4052 (.ZN(n1866), 
	.A(n4839));
   AOI221_X1 U4053 (.ZN(n2476), 
	.C2(n2486), 
	.C1(n1931), 
	.B2(n1870), 
	.B1(n1930), 
	.A(n2487));
   OAI22_X1 U4054 (.ZN(n2487), 
	.B2(n6373), 
	.B1(n5063), 
	.A2(n1934), 
	.A1(n4455));
   INV_X1 U4055 (.ZN(n2486), 
	.A(n5287));
   INV_X1 U4056 (.ZN(n1870), 
	.A(n5319));
   AOI222_X1 U4057 (.ZN(n2475), 
	.C2(n1938), 
	.C1(n1874), 
	.B2(n1873), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1872));
   INV_X1 U4058 (.ZN(n1874), 
	.A(n4487));
   INV_X1 U4059 (.ZN(n1873), 
	.A(n4423));
   INV_X1 U4060 (.ZN(n1872), 
	.A(n4519));
   AOI22_X1 U4064 (.ZN(n2489), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [6]), 
	.B1(n906), 
	.A2(\UUT/break_code[6] ), 
	.A1(n908));
   OAI21_X1 U4065 (.ZN(\UUT/break_code[6] ), 
	.B2(n2072), 
	.B1(n6143), 
	.A(n2490));
   NAND2_X1 U4066 (.ZN(n2490), 
	.A2(n2074), 
	.A1(n6234));
   INV_X1 U4067 (.ZN(n6143), 
	.A(\UUT/Mcontrol/d_sampled_finstr [6]));
   AOI222_X1 U4069 (.ZN(n5441), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[6] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n692), 
	.A2(n5564), 
	.A1(n6192));
   NAND2_X1 U4070 (.ZN(n692), 
	.A2(n2493), 
	.A1(n2492));
   AOI222_X1 U4071 (.ZN(n2493), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [6]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [6]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [6]));
   AOI22_X1 U4072 (.ZN(n2492), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [6]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [6]));
   NAND3_X1 U4073 (.ZN(n6192), 
	.A3(n2496), 
	.A2(n2495), 
	.A1(n2494));
   AOI222_X1 U4074 (.ZN(n2496), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[6] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[6] ), 
	.A2(n2497), 
	.A1(n1208));
   INV_X1 U4075 (.ZN(n2497), 
	.A(\UUT/Mpath/the_alu/N71 ));
   AOI22_X1 U4076 (.ZN(n2495), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N119 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N151 ));
   AOI22_X1 U4077 (.ZN(n2494), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N215 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N183 ));
   INV_X1 U4078 (.ZN(n2491), 
	.A(n679));
   NAND4_X1 U4079 (.ZN(n679), 
	.A4(FE_OFN71_n2501), 
	.A3(n2500), 
	.A2(n2499), 
	.A1(n2498));
   NOR4_X1 U4080 (.ZN(n2501), 
	.A4(n2505), 
	.A3(n2504), 
	.A2(n2503), 
	.A1(n2502));
   NAND3_X1 U4081 (.ZN(n2505), 
	.A3(n6233), 
	.A2(n6231), 
	.A1(n6232));
   OAI211_X1 U4082 (.ZN(n2504), 
	.C2(n5384), 
	.C1(n5560), 
	.B(n6230), 
	.A(n6229));
   OAI222_X1 U4083 (.ZN(n2503), 
	.C2(n5352), 
	.C1(n5561), 
	.B2(n5224), 
	.B1(n5559), 
	.A2(n5256), 
	.A1(n5558));
   OAI221_X1 U4084 (.ZN(n2502), 
	.C2(n5192), 
	.C1(n5532), 
	.B2(n5160), 
	.B1(n5531), 
	.A(n2506));
   AOI22_X1 U4085 (.ZN(n2506), 
	.B2(n1926), 
	.B1(n1845), 
	.A2(n1925), 
	.A1(n1844));
   INV_X1 U4086 (.ZN(n1845), 
	.A(n4968));
   INV_X1 U4087 (.ZN(n1844), 
	.A(n4936));
   AOI211_X1 U4088 (.ZN(n2500), 
	.C2(n1927), 
	.C1(n1846), 
	.B(n2508), 
	.A(n2507));
   OAI22_X1 U4089 (.ZN(n2508), 
	.B2(n4712), 
	.B1(n5551), 
	.A2(n4808), 
	.A1(n5541));
   OAI222_X1 U4090 (.ZN(n2507), 
	.C2(n4680), 
	.C1(n5547), 
	.B2(n4616), 
	.B1(n5552), 
	.A2(n4648), 
	.A1(n5546));
   INV_X1 U4091 (.ZN(n1846), 
	.A(n4840));
   AOI221_X1 U4092 (.ZN(n2499), 
	.C2(n2509), 
	.C1(n1931), 
	.B2(n1850), 
	.B1(n1930), 
	.A(n2510));
   OAI22_X1 U4093 (.ZN(n2510), 
	.B2(n6373), 
	.B1(n5064), 
	.A2(n1934), 
	.A1(n4456));
   INV_X1 U4094 (.ZN(n2509), 
	.A(n5288));
   INV_X1 U4095 (.ZN(n1850), 
	.A(n5320));
   AOI222_X1 U4096 (.ZN(n2498), 
	.C2(n1938), 
	.C1(n1854), 
	.B2(n1853), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1852));
   INV_X1 U4097 (.ZN(n1854), 
	.A(n4488));
   INV_X1 U4098 (.ZN(n1853), 
	.A(n4424));
   INV_X1 U4099 (.ZN(n1852), 
	.A(n4520));
   OAI21_X1 U4104 (.ZN(\UUT/break_code[5] ), 
	.B2(n2072), 
	.B1(n5423), 
	.A(n2513));
   NAND2_X1 U4105 (.ZN(n2513), 
	.A2(n2074), 
	.A1(n6240));
   OAI21_X1 U4107 (.ZN(n2072), 
	.B2(n2514), 
	.B1(n6170), 
	.A(n6030));
   NOR2_X1 U4108 (.ZN(n2514), 
	.A2(n445), 
	.A1(n2070));
   INV_X1 U4109 (.ZN(n445), 
	.A(n6209));
   INV_X1 U4110 (.ZN(n2070), 
	.A(n6172));
   NAND2_X1 U4111 (.ZN(n6170), 
	.A2(n929), 
	.A1(n932));
   NOR2_X1 U4112 (.ZN(n929), 
	.A2(n1219), 
	.A1(n2077));
   OAI21_X1 U4113 (.ZN(n1219), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N2071 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2066 ));
   NAND2_X1 U4114 (.ZN(n2077), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
	.A1(n915));
   INV_X1 U4115 (.ZN(n915), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2079 ));
   NOR2_X1 U4116 (.ZN(n932), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2061 ), 
	.A1(n1004));
   NAND2_X1 U4117 (.ZN(n1004), 
	.A2(n924), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2054 ));
   OR2_X1 U4118 (.ZN(n924), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2047 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   INV_X1 U4119 (.ZN(n5423), 
	.A(\UUT/Mcontrol/d_sampled_finstr [5]));
   OAI222_X1 U4120 (.ZN(\UUT/branch_rega [5]), 
	.C2(FE_OFN17_n5444), 
	.C1(n5528), 
	.B2(n2515), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5446));
   AOI222_X1 U4121 (.ZN(n5444), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[5] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n715), 
	.A2(n5564), 
	.A1(n6193));
   NAND2_X1 U4122 (.ZN(n715), 
	.A2(n2517), 
	.A1(n2516));
   AOI222_X1 U4123 (.ZN(n2517), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [5]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [5]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [5]));
   AOI22_X1 U4124 (.ZN(n2516), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [5]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [5]));
   NAND3_X1 U4125 (.ZN(n6193), 
	.A3(n2520), 
	.A2(n2519), 
	.A1(n2518));
   AOI222_X1 U4126 (.ZN(n2520), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[5] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[5] ), 
	.A2(n2521), 
	.A1(n1208));
   INV_X1 U4127 (.ZN(n2521), 
	.A(\UUT/Mpath/the_alu/N73 ));
   AOI22_X1 U4128 (.ZN(n2519), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N120 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N152 ));
   AOI22_X1 U4129 (.ZN(n2518), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N216 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N184 ));
   INV_X1 U4130 (.ZN(n2515), 
	.A(n707));
   NAND4_X1 U4131 (.ZN(n707), 
	.A4(FE_OFN74_n2525), 
	.A3(n2524), 
	.A2(n2523), 
	.A1(n2522));
   NOR4_X1 U4132 (.ZN(n2525), 
	.A4(n2529), 
	.A3(n2528), 
	.A2(n2527), 
	.A1(n2526));
   NAND3_X1 U4133 (.ZN(n2529), 
	.A3(n6239), 
	.A2(n6237), 
	.A1(n6238));
   OAI211_X1 U4134 (.ZN(n2528), 
	.C2(n5385), 
	.C1(n5560), 
	.B(n6236), 
	.A(n6235));
   OAI222_X1 U4135 (.ZN(n2527), 
	.C2(n5353), 
	.C1(n5561), 
	.B2(n5225), 
	.B1(n5559), 
	.A2(n5257), 
	.A1(n5558));
   OAI221_X1 U4136 (.ZN(n2526), 
	.C2(n5193), 
	.C1(n5532), 
	.B2(n5161), 
	.B1(n5531), 
	.A(n2530));
   AOI22_X1 U4137 (.ZN(n2530), 
	.B2(n1926), 
	.B1(n1825), 
	.A2(n1925), 
	.A1(n1824));
   INV_X1 U4138 (.ZN(n1825), 
	.A(n4969));
   INV_X1 U4139 (.ZN(n1824), 
	.A(n4937));
   AOI211_X1 U4140 (.ZN(n2524), 
	.C2(n1927), 
	.C1(n1826), 
	.B(n2532), 
	.A(n2531));
   OAI22_X1 U4141 (.ZN(n2532), 
	.B2(n4713), 
	.B1(n5551), 
	.A2(n4809), 
	.A1(n5541));
   OAI222_X1 U4142 (.ZN(n2531), 
	.C2(n4681), 
	.C1(n5547), 
	.B2(n4617), 
	.B1(n5552), 
	.A2(n4649), 
	.A1(n5546));
   INV_X1 U4143 (.ZN(n1826), 
	.A(n4841));
   AOI221_X1 U4144 (.ZN(n2523), 
	.C2(n2533), 
	.C1(n1931), 
	.B2(n1830), 
	.B1(n1930), 
	.A(n2534));
   OAI22_X1 U4145 (.ZN(n2534), 
	.B2(n6373), 
	.B1(n5065), 
	.A2(n1934), 
	.A1(n4457));
   INV_X1 U4146 (.ZN(n2533), 
	.A(n5289));
   INV_X1 U4147 (.ZN(n1830), 
	.A(n5321));
   AOI222_X1 U4148 (.ZN(n2522), 
	.C2(n1938), 
	.C1(n1834), 
	.B2(n1833), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1832));
   INV_X1 U4149 (.ZN(n1834), 
	.A(n4489));
   INV_X1 U4150 (.ZN(n1833), 
	.A(n4425));
   INV_X1 U4151 (.ZN(n1832), 
	.A(n4521));
   INV_X1 U4156 (.ZN(\UUT/break_code[4] ), 
	.A(n718));
   AOI22_X1 U4157 (.ZN(n718), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [4]), 
	.B1(n2329), 
	.A2(n2328), 
	.A1(n6247));
   OAI222_X1 U4158 (.ZN(\UUT/branch_rega [4]), 
	.C2(FE_OFN190_n5447), 
	.C1(n5528), 
	.B2(n2537), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5449));
   AOI222_X1 U4159 (.ZN(n5447), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[4] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n738), 
	.A2(n5564), 
	.A1(n6194));
   NAND2_X1 U4160 (.ZN(n738), 
	.A2(n2539), 
	.A1(n2538));
   AOI222_X1 U4161 (.ZN(n2539), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [4]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [4]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [4]));
   AOI22_X1 U4162 (.ZN(n2538), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [4]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [4]));
   NAND3_X1 U4163 (.ZN(n6194), 
	.A3(n2542), 
	.A2(n2541), 
	.A1(n2540));
   AOI222_X1 U4164 (.ZN(n2542), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[4] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[4] ), 
	.A2(n2543), 
	.A1(n1208));
   INV_X1 U4165 (.ZN(n2543), 
	.A(\UUT/Mpath/the_alu/N75 ));
   AOI22_X1 U4166 (.ZN(n2541), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N121 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N153 ));
   AOI22_X1 U4167 (.ZN(n2540), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N217 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N185 ));
   INV_X1 U4168 (.ZN(n2537), 
	.A(n730));
   NAND4_X1 U4169 (.ZN(n730), 
	.A4(FE_OFN77_n2547), 
	.A3(n2546), 
	.A2(n2545), 
	.A1(n2544));
   NOR4_X1 U4170 (.ZN(n2547), 
	.A4(n2551), 
	.A3(n2550), 
	.A2(n2549), 
	.A1(n2548));
   NAND3_X1 U4171 (.ZN(n2551), 
	.A3(n6245), 
	.A2(n6243), 
	.A1(n6244));
   OAI211_X1 U4172 (.ZN(n2550), 
	.C2(n5386), 
	.C1(n5560), 
	.B(n6242), 
	.A(n6241));
   OAI222_X1 U4173 (.ZN(n2549), 
	.C2(n5354), 
	.C1(n5561), 
	.B2(n5226), 
	.B1(n5559), 
	.A2(n5258), 
	.A1(n5558));
   OAI221_X1 U4174 (.ZN(n2548), 
	.C2(n5194), 
	.C1(n5532), 
	.B2(n5162), 
	.B1(n5531), 
	.A(n2552));
   AOI22_X1 U4175 (.ZN(n2552), 
	.B2(n1926), 
	.B1(n1805), 
	.A2(n1925), 
	.A1(n1804));
   INV_X1 U4176 (.ZN(n1805), 
	.A(n4970));
   INV_X1 U4177 (.ZN(n1804), 
	.A(n4938));
   AOI211_X1 U4178 (.ZN(n2546), 
	.C2(n1927), 
	.C1(n1806), 
	.B(n2554), 
	.A(n2553));
   OAI22_X1 U4179 (.ZN(n2554), 
	.B2(n4714), 
	.B1(n5551), 
	.A2(n4810), 
	.A1(n5541));
   OAI222_X1 U4180 (.ZN(n2553), 
	.C2(n4682), 
	.C1(n5547), 
	.B2(n4618), 
	.B1(n5552), 
	.A2(n4650), 
	.A1(n5546));
   INV_X1 U4181 (.ZN(n1806), 
	.A(n4842));
   AOI221_X1 U4182 (.ZN(n2545), 
	.C2(n2555), 
	.C1(n1931), 
	.B2(n1810), 
	.B1(n1930), 
	.A(n2556));
   OAI22_X1 U4183 (.ZN(n2556), 
	.B2(n6373), 
	.B1(n5066), 
	.A2(n1934), 
	.A1(n4458));
   INV_X1 U4184 (.ZN(n2555), 
	.A(n5290));
   INV_X1 U4185 (.ZN(n1810), 
	.A(n5322));
   AOI222_X1 U4186 (.ZN(n2544), 
	.C2(n1938), 
	.C1(n1814), 
	.B2(n1813), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1812));
   INV_X1 U4187 (.ZN(n1814), 
	.A(n4490));
   INV_X1 U4188 (.ZN(n1813), 
	.A(n4426));
   INV_X1 U4189 (.ZN(n1812), 
	.A(n4522));
   AOI22_X1 U4193 (.ZN(n2558), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [3]), 
	.B1(n906), 
	.A2(\UUT/break_code[3] ), 
	.A1(n908));
   INV_X1 U4195 (.ZN(n2559), 
	.A(n2561));
   INV_X1 U4196 (.ZN(\UUT/break_code[3] ), 
	.A(FE_OFN197_n741));
   AOI22_X1 U4197 (.ZN(n741), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [3]), 
	.B1(n2329), 
	.A2(n2328), 
	.A1(n6255));
   OAI21_X1 U4198 (.ZN(n2329), 
	.B2(n2562), 
	.B1(n6246), 
	.A(n2563));
   INV_X1 U4199 (.ZN(n2563), 
	.A(n6266));
   AND2_X1 U4200 (.ZN(n2328), 
	.A2(n913), 
	.A1(n6246));
   INV_X1 U4201 (.ZN(n913), 
	.A(n2562));
   NAND2_X1 U4202 (.ZN(n2562), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2084 ), 
	.A1(n6030));
   INV_X1 U4203 (.ZN(n6030), 
	.A(n933));
   NOR2_X1 U4204 (.ZN(n933), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2083 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   AND3_X1 U4205 (.ZN(n908), 
	.A3(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.A2(n2564), 
	.A1(\UUT/Mcontrol/st_logic/N65 ));
   AOI222_X1 U4207 (.ZN(n5450), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[3] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n761), 
	.A2(n5564), 
	.A1(n6195));
   NAND2_X1 U4208 (.ZN(n761), 
	.A2(n2567), 
	.A1(n2566));
   AOI222_X1 U4209 (.ZN(n2567), 
	.C2(n6199), 
	.C1(\UUT/Mpath/the_shift/sh_rol [3]), 
	.B2(\UUT/Mpath/the_shift/N118 ), 
	.B1(\UUT/Mpath/the_shift/sh_srl [3]), 
	.A2(FE_OFN88_n6201), 
	.A1(\UUT/Mpath/the_shift/sh_ror [3]));
   AOI22_X1 U4210 (.ZN(n2566), 
	.B2(n6198), 
	.B1(\UUT/Mpath/the_shift/sh_sra [3]), 
	.A2(n6200), 
	.A1(\UUT/Mpath/the_shift/sh_sll [3]));
   NAND3_X1 U4211 (.ZN(n6195), 
	.A3(n2570), 
	.A2(n2569), 
	.A1(n2568));
   AOI222_X1 U4212 (.ZN(n2570), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[3] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[3] ), 
	.A2(n2571), 
	.A1(n1208));
   INV_X1 U4214 (.ZN(n2572), 
	.A(n2047));
   INV_X1 U4215 (.ZN(n2571), 
	.A(\UUT/Mpath/the_alu/N77 ));
   INV_X1 U4217 (.ZN(n2573), 
	.A(n2574));
   AOI22_X1 U4218 (.ZN(n2569), 
	.B2(n1213), 
	.B1(\UUT/Mpath/the_alu/N122 ), 
	.A2(n1212), 
	.A1(\UUT/Mpath/the_alu/N154 ));
   INV_X1 U4220 (.ZN(\UUT/Mpath/the_alu/N492 ), 
	.A(\UUT/Mpath/the_alu/N491 ));
   NOR4_X1 U4221 (.ZN(n6348), 
	.A4(\UUT/Mpath/the_alu/N498 ), 
	.A3(n2050), 
	.A2(FE_OFN87_n1211), 
	.A1(n2047));
   INV_X1 U4222 (.ZN(n2050), 
	.A(\UUT/Mpath/the_alu/N503 ));
   INV_X1 U4224 (.ZN(n2575), 
	.A(\UUT/Mpath/the_alu/N468 ));
   NAND2_X1 U4225 (.ZN(n2047), 
	.A2(\UUT/Mpath/the_alu/N509 ), 
	.A1(\UUT/Mpath/the_alu/N515 ));
   INV_X1 U4227 (.ZN(n2576), 
	.A(\UUT/Mpath/the_alu/N486 ));
   AOI22_X1 U4228 (.ZN(n2568), 
	.B2(n1215), 
	.B1(\UUT/Mpath/the_alu/N218 ), 
	.A2(FE_OFN86_n1214), 
	.A1(\UUT/Mpath/the_alu/N186 ));
   NOR3_X1 U4230 (.ZN(n2574), 
	.A3(\UUT/Mpath/the_alu/N480 ), 
	.A2(n6349), 
	.A1(\UUT/Mpath/the_alu/N486 ));
   INV_X1 U4232 (.ZN(n2577), 
	.A(\UUT/Mpath/the_alu/N480 ));
   INV_X1 U4234 (.ZN(n2565), 
	.A(n753));
   NAND4_X1 U4235 (.ZN(n753), 
	.A4(FE_OFN80_n2581), 
	.A3(n2580), 
	.A2(n2579), 
	.A1(n2578));
   NOR4_X1 U4236 (.ZN(n2581), 
	.A4(n2585), 
	.A3(n2584), 
	.A2(n2583), 
	.A1(n2582));
   NAND3_X1 U4237 (.ZN(n2585), 
	.A3(n6254), 
	.A2(n6252), 
	.A1(n6253));
   OAI211_X1 U4238 (.ZN(n2584), 
	.C2(n5387), 
	.C1(n5560), 
	.B(n6251), 
	.A(n6250));
   OAI222_X1 U4239 (.ZN(n2583), 
	.C2(n5355), 
	.C1(n5561), 
	.B2(n5227), 
	.B1(n5559), 
	.A2(n5259), 
	.A1(n5558));
   OAI221_X1 U4240 (.ZN(n2582), 
	.C2(n5195), 
	.C1(n5532), 
	.B2(n5163), 
	.B1(n5531), 
	.A(n2586));
   AOI22_X1 U4241 (.ZN(n2586), 
	.B2(n1926), 
	.B1(n1785), 
	.A2(n1925), 
	.A1(n1784));
   INV_X1 U4243 (.ZN(n1785), 
	.A(n4971));
   INV_X1 U4245 (.ZN(n1784), 
	.A(n4939));
   AOI211_X1 U4246 (.ZN(n2580), 
	.C2(n1927), 
	.C1(n1786), 
	.B(n2588), 
	.A(n2587));
   OAI22_X1 U4247 (.ZN(n2588), 
	.B2(n4715), 
	.B1(n5551), 
	.A2(n4811), 
	.A1(n5541));
   OAI222_X1 U4248 (.ZN(n2587), 
	.C2(n4683), 
	.C1(n5547), 
	.B2(n4619), 
	.B1(n5552), 
	.A2(n4651), 
	.A1(n5546));
   INV_X1 U4250 (.ZN(n1786), 
	.A(n4843));
   AOI221_X1 U4251 (.ZN(n2579), 
	.C2(n2589), 
	.C1(n1931), 
	.B2(n1790), 
	.B1(n1930), 
	.A(n2590));
   OAI22_X1 U4252 (.ZN(n2590), 
	.B2(n6373), 
	.B1(n5067), 
	.A2(n1934), 
	.A1(n4459));
   INV_X1 U4255 (.ZN(n2589), 
	.A(n5291));
   INV_X1 U4257 (.ZN(n1790), 
	.A(n5323));
   INV_X1 U4259 (.ZN(n2591), 
	.A(n6318));
   AOI222_X1 U4260 (.ZN(n2578), 
	.C2(n1938), 
	.C1(n1794), 
	.B2(n1793), 
	.B1(n1937), 
	.A2(n1936), 
	.A1(n1792));
   INV_X1 U4262 (.ZN(n1794), 
	.A(n4491));
   INV_X1 U4263 (.ZN(n1793), 
	.A(n4427));
   INV_X1 U4266 (.ZN(n1792), 
	.A(n4523));
   INV_X1 U4269 (.ZN(n2592), 
	.A(n6303));
   INV_X1 U4271 (.ZN(\UUT/byp_controlA[0] ), 
	.A(\UUT/Mcontrol/st_logic/N47 ));
   NAND2_X1 U4272 (.ZN(\UUT/Mcontrol/st_logic/N47 ), 
	.A2(n2594), 
	.A1(\UUT/Mcontrol/bp_logicA/memory_main ));
   INV_X1 U4273 (.ZN(n2594), 
	.A(\UUT/Mcontrol/bp_logicA/exec_main ));
   AOI21_X1 U4276 (.ZN(n2561), 
	.B2(\UUT/Mcontrol/st_logic/N65 ), 
	.B1(n2564), 
	.A(\UUT/Mcontrol/st_logic/N109 ));
   INV_X1 U4278 (.ZN(n2564), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N116 ));
   INV_X1 U4279 (.ZN(n2560), 
	.A(\UUT/Mcontrol/st_logic/N103 ));
   INV_X1 U4280 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2085 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2084 ));
   NOR2_X1 U4281 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2079 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2071 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   INV_X1 U4282 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2061 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2060 ));
   NOR2_X1 U4283 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2043 ), 
	.A2(\UUT/Mcontrol/d_instr [26]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2041 ));
   NOR2_X1 U4284 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2023 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   NOR2_X1 U4285 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1993 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   NOR2_X1 U4286 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2007 ), 
	.A2(\UUT/Mcontrol/d_instr [26]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2005 ));
   NOR2_X1 U4287 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2001 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1974 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1922 ));
   INV_X1 U4288 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1995 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1994 ));
   INV_X1 U4289 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1976 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1975 ));
   INV_X1 U4290 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1922 ), 
	.A(\UUT/Mcontrol/d_instr [26]));
   INV_X1 U4300 (.ZN(n4339), 
	.A(\localbus/N338 ));
   INV_X1 U4303 (.ZN(n4340), 
	.A(\localbus/N62 ));
   NOR2_X1 U4304 (.ZN(\localbus/c1_op[OP][1] ), 
	.A2(n4343), 
	.A1(\localbus/c1_op[OP][0] ));
   INV_X1 U4305 (.ZN(n4343), 
	.A(\localbus/N46 ));
   NOR2_X1 U4306 (.ZN(\localbus/c1_op[MASTER] ), 
	.A2(\localbus/N46 ), 
	.A1(\localbus/c1_op[OP][0] ));
   INV_X1 U4315 (.ZN(\localbus/c1_addr_outbus[30] ), 
	.A(n4352));
   INV_X1 U4317 (.ZN(\localbus/c1_addr_outbus[29] ), 
	.A(n4354));
   INV_X1 U4318 (.ZN(\localbus/c1_addr_outbus[28] ), 
	.A(n4355));
   INV_X1 U4319 (.ZN(\localbus/c1_addr_outbus[27] ), 
	.A(n4356));
   INV_X1 U4320 (.ZN(\localbus/c1_addr_outbus[26] ), 
	.A(n4357));
   INV_X1 U4321 (.ZN(\localbus/c1_addr_outbus[25] ), 
	.A(n4358));
   INV_X1 U4322 (.ZN(\localbus/c1_addr_outbus[24] ), 
	.A(n4359));
   INV_X1 U4323 (.ZN(\localbus/c1_addr_outbus[23] ), 
	.A(n4360));
   INV_X1 U4324 (.ZN(\localbus/c1_addr_outbus[22] ), 
	.A(n4361));
   INV_X1 U4325 (.ZN(\localbus/c1_addr_outbus[21] ), 
	.A(n4362));
   INV_X1 U4326 (.ZN(\localbus/c1_addr_outbus[20] ), 
	.A(n4363));
   INV_X1 U4328 (.ZN(\localbus/c1_addr_outbus[19] ), 
	.A(n4365));
   INV_X1 U4329 (.ZN(\localbus/c1_addr_outbus[18] ), 
	.A(n4366));
   INV_X1 U4330 (.ZN(\localbus/c1_addr_outbus[17] ), 
	.A(n4367));
   INV_X1 U4331 (.ZN(\localbus/c1_addr_outbus[16] ), 
	.A(n4368));
   INV_X1 U4332 (.ZN(\localbus/c1_addr_outbus[15] ), 
	.A(n4369));
   INV_X1 U4333 (.ZN(\localbus/c1_addr_outbus[14] ), 
	.A(n4370));
   INV_X1 U4334 (.ZN(\localbus/c1_addr_outbus[13] ), 
	.A(n4371));
   INV_X1 U4339 (.ZN(dram_mw), 
	.A(\localbus/N89 ));
   INV_X1 U4340 (.ZN(dram_mr), 
	.A(\localbus/N85 ));
   NOR2_X1 U4341 (.ZN(dram_data_outbus[9]), 
	.A2(n4377), 
	.A1(n4376));
   NOR2_X1 U4342 (.ZN(dram_data_outbus[8]), 
	.A2(n4377), 
	.A1(n4378));
   NOR2_X1 U4343 (.ZN(dram_data_outbus[7]), 
	.A2(n4380), 
	.A1(n4379));
   NOR2_X1 U4344 (.ZN(dram_data_outbus[6]), 
	.A2(n4381), 
	.A1(n4379));
   NOR2_X1 U4345 (.ZN(dram_data_outbus[5]), 
	.A2(n4382), 
	.A1(n4379));
   NOR2_X1 U4346 (.ZN(dram_data_outbus[4]), 
	.A2(n4383), 
	.A1(n4379));
   NOR2_X1 U4347 (.ZN(dram_data_outbus[3]), 
	.A2(n4384), 
	.A1(n4379));
   NOR2_X1 U4348 (.ZN(dram_data_outbus[31]), 
	.A2(n4377), 
	.A1(n4385));
   NOR2_X1 U4349 (.ZN(dram_data_outbus[30]), 
	.A2(n4377), 
	.A1(n4386));
   NOR2_X1 U4350 (.ZN(dram_data_outbus[2]), 
	.A2(n4387), 
	.A1(n4379));
   NOR2_X1 U4351 (.ZN(dram_data_outbus[29]), 
	.A2(n4377), 
	.A1(n4388));
   NOR2_X1 U4352 (.ZN(dram_data_outbus[28]), 
	.A2(n4377), 
	.A1(n4389));
   NOR2_X1 U4353 (.ZN(dram_data_outbus[27]), 
	.A2(n4377), 
	.A1(n4390));
   NOR2_X1 U4354 (.ZN(dram_data_outbus[26]), 
	.A2(n4377), 
	.A1(n4391));
   NOR2_X1 U4355 (.ZN(dram_data_outbus[25]), 
	.A2(n4377), 
	.A1(n4392));
   NOR2_X1 U4356 (.ZN(dram_data_outbus[24]), 
	.A2(n4377), 
	.A1(n4393));
   NOR2_X1 U4357 (.ZN(dram_data_outbus[23]), 
	.A2(n4377), 
	.A1(n4394));
   NOR2_X1 U4358 (.ZN(dram_data_outbus[22]), 
	.A2(n4377), 
	.A1(n4395));
   NOR2_X1 U4359 (.ZN(dram_data_outbus[21]), 
	.A2(n4377), 
	.A1(n4396));
   NOR2_X1 U4360 (.ZN(dram_data_outbus[20]), 
	.A2(n4377), 
	.A1(n4397));
   NOR2_X1 U4361 (.ZN(dram_data_outbus[1]), 
	.A2(n4379), 
	.A1(n4398));
   NOR2_X1 U4362 (.ZN(dram_data_outbus[19]), 
	.A2(n4377), 
	.A1(n4399));
   NOR2_X1 U4363 (.ZN(dram_data_outbus[18]), 
	.A2(n4377), 
	.A1(n4400));
   NOR2_X1 U4364 (.ZN(dram_data_outbus[17]), 
	.A2(n4377), 
	.A1(n4401));
   NOR2_X1 U4365 (.ZN(dram_data_outbus[16]), 
	.A2(n4377), 
	.A1(n4402));
   NOR2_X1 U4366 (.ZN(dram_data_outbus[15]), 
	.A2(n4377), 
	.A1(n4403));
   NOR2_X1 U4367 (.ZN(dram_data_outbus[14]), 
	.A2(n4377), 
	.A1(n4404));
   NOR2_X1 U4368 (.ZN(dram_data_outbus[13]), 
	.A2(n4377), 
	.A1(n4405));
   NOR2_X1 U4369 (.ZN(dram_data_outbus[12]), 
	.A2(n4377), 
	.A1(n4406));
   NOR2_X1 U4370 (.ZN(dram_data_outbus[11]), 
	.A2(n4377), 
	.A1(n4407));
   NOR2_X1 U4371 (.ZN(dram_data_outbus[10]), 
	.A2(n4377), 
	.A1(n4408));
   INV_X1 U4372 (.ZN(n4377), 
	.A(\localbus/N218 ));
   NOR2_X1 U4373 (.ZN(dram_data_outbus[0]), 
	.A2(n4379), 
	.A1(n4409));
   NAND2_X1 U4374 (.ZN(n4379), 
	.A2(\localbus/N51 ), 
	.A1(\localbus/N218 ));
   NOR2_X1 U4375 (.ZN(dram_addr_outbus[9]), 
	.A2(\localbus/N214 ), 
	.A1(n4344));
   NOR2_X1 U4376 (.ZN(dram_addr_outbus[8]), 
	.A2(n4345), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4377 (.ZN(dram_addr_outbus[7]), 
	.A2(n4346), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4378 (.ZN(dram_addr_outbus[6]), 
	.A2(n4347), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4379 (.ZN(dram_addr_outbus[5]), 
	.A2(n4348), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4380 (.ZN(dram_addr_outbus[4]), 
	.A2(n4349), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4381 (.ZN(dram_addr_outbus[3]), 
	.A2(n4350), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4382 (.ZN(dram_addr_outbus[2]), 
	.A2(n4353), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4383 (.ZN(dram_addr_outbus[12]), 
	.A2(n4372), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4384 (.ZN(dram_addr_outbus[11]), 
	.A2(n4373), 
	.A1(\localbus/N214 ));
   NOR2_X1 U4385 (.ZN(dram_addr_outbus[10]), 
	.A2(n4374), 
	.A1(\localbus/N214 ));
   AND4_X1 U4387 (.ZN(d_select[31]), 
	.A4(n4414), 
	.A3(n4413), 
	.A2(n4412), 
	.A1(n4411));
   NAND2_X1 U4388 (.ZN(n4411), 
	.A2(n4416), 
	.A1(n4415));
   INV_X1 U4389 (.ZN(n4416), 
	.A(N35));
   AND3_X1 U4390 (.ZN(d_select[23]), 
	.A3(n4417), 
	.A2(n4413), 
	.A1(n4412));
   OAI21_X1 U4391 (.ZN(n4417), 
	.B2(n4415), 
	.B1(N35), 
	.A(n4414));
   INV_X1 U4392 (.ZN(n4414), 
	.A(N31));
   NOR2_X1 U4393 (.ZN(n4415), 
	.A2(N42), 
	.A1(N43));
   INV_X1 U4394 (.ZN(n4413), 
	.A(N27));
   INV_X1 U4395 (.ZN(n4412), 
	.A(N22));
   OAI21_X1 U4396 (.ZN(d_select[9]), 
	.B2(n4418), 
	.B1(N43), 
	.A(n4419));
   INV_X1 U4397 (.ZN(n4418), 
	.A(N42));
   NAND2_X1 U4398 (.ZN(d_select[7]), 
	.A2(n4420), 
	.A1(n4419));
   INV_X1 U4399 (.ZN(n4420), 
	.A(N43));
   NOR4_X1 U4400 (.ZN(n4419), 
	.A4(N35), 
	.A3(N31), 
	.A2(N27), 
	.A1(N22));
   OR2_X1 U4401 (.ZN(dmem_write), 
	.A2(\UUT/x_we ), 
	.A1(\UUT/Mcontrol/x_sampled_dmem_command[MW] ));
   AND2_X1 U4402 (.ZN(\UUT/regfile/N358 ), 
	.A2(n5413), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[4] ));
   AND2_X1 U4403 (.ZN(\UUT/rd_addr [3]), 
	.A2(n5413), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[3] ));
   AND2_X1 U4404 (.ZN(\UUT/rd_addr [2]), 
	.A2(n5413), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[2] ));
   AND2_X1 U4405 (.ZN(\UUT/rd_addr [1]), 
	.A2(n5413), 
	.A1(\UUT/Mcontrol/m_sampled_xrd[1] ));
   OR2_X1 U4406 (.ZN(\UUT/byp_controlB[2] ), 
	.A2(\UUT/Mcontrol/bp_logicB/exec_main ), 
	.A1(\UUT/Mcontrol/bp_logicB/memory_main ));
   OR2_X1 U4407 (.ZN(\UUT/byp_controlA[2] ), 
	.A2(\UUT/Mcontrol/bp_logicA/exec_main ), 
	.A1(\UUT/Mcontrol/bp_logicA/memory_main ));
   OAI222_X1 U4408 (.ZN(\UUT/branch_regb [9]), 
	.C2(n5434), 
	.C1(n5433), 
	.B2(n5432), 
	.B1(n5431), 
	.A2(n5430), 
	.A1(FE_OFN194_n5429));
   OAI222_X1 U4409 (.ZN(\UUT/branch_regb [8]), 
	.C2(n5434), 
	.C1(n5437), 
	.B2(n5432), 
	.B1(n5436), 
	.A2(n5430), 
	.A1(FE_OFN191_n5435));
   OAI222_X1 U4410 (.ZN(\UUT/branch_regb [7]), 
	.C2(n5434), 
	.C1(n5440), 
	.B2(n5432), 
	.B1(n5439), 
	.A2(n5430), 
	.A1(FE_OFN195_n5438));
   OAI222_X1 U4411 (.ZN(\UUT/branch_regb [6]), 
	.C2(n5434), 
	.C1(n5443), 
	.B2(n5432), 
	.B1(n5442), 
	.A2(n5430), 
	.A1(FE_OFN18_n5441));
   OAI222_X1 U4412 (.ZN(\UUT/branch_regb [5]), 
	.C2(n5434), 
	.C1(n5446), 
	.B2(n5432), 
	.B1(n5445), 
	.A2(n5430), 
	.A1(FE_OFN17_n5444));
   OAI222_X1 U4413 (.ZN(\UUT/branch_regb [4]), 
	.C2(n5434), 
	.C1(n5449), 
	.B2(n5432), 
	.B1(n5448), 
	.A2(n5430), 
	.A1(FE_OFN190_n5447));
   OAI222_X1 U4414 (.ZN(\UUT/branch_regb [3]), 
	.C2(n5434), 
	.C1(n5452), 
	.B2(n5432), 
	.B1(n5451), 
	.A2(n5430), 
	.A1(FE_OFN30_n5450));
   OAI222_X1 U4416 (.ZN(\UUT/branch_regb [30]), 
	.C2(n5434), 
	.C1(n5458), 
	.B2(n5432), 
	.B1(n5457), 
	.A2(n5430), 
	.A1(n5456));
   OAI222_X1 U4417 (.ZN(\UUT/branch_regb [2]), 
	.C2(n5434), 
	.C1(n5461), 
	.B2(n5432), 
	.B1(n5460), 
	.A2(n5430), 
	.A1(FE_OFN189_n5459));
   OAI222_X1 U4419 (.ZN(\UUT/branch_regb [28]), 
	.C2(n5434), 
	.C1(n5467), 
	.B2(n5432), 
	.B1(n5466), 
	.A2(n5430), 
	.A1(n5465));
   OAI222_X1 U4422 (.ZN(\UUT/branch_regb [25]), 
	.C2(n5434), 
	.C1(n5476), 
	.B2(n5432), 
	.B1(n5475), 
	.A2(n5430), 
	.A1(n5474));
   OAI222_X1 U4423 (.ZN(\UUT/branch_regb [24]), 
	.C2(n5434), 
	.C1(n5479), 
	.B2(n5432), 
	.B1(n5478), 
	.A2(n5430), 
	.A1(n5477));
   OAI222_X1 U4424 (.ZN(\UUT/branch_regb [23]), 
	.C2(n5434), 
	.C1(n5482), 
	.B2(n5432), 
	.B1(n5481), 
	.A2(n5430), 
	.A1(n5480));
   OAI222_X1 U4425 (.ZN(\UUT/branch_regb [22]), 
	.C2(n5434), 
	.C1(n5485), 
	.B2(n5432), 
	.B1(n5484), 
	.A2(n5430), 
	.A1(n5483));
   OAI222_X1 U4426 (.ZN(\UUT/branch_regb [21]), 
	.C2(n5434), 
	.C1(n5488), 
	.B2(n5432), 
	.B1(n5487), 
	.A2(n5430), 
	.A1(n5486));
   OAI222_X1 U4427 (.ZN(\UUT/branch_regb [20]), 
	.C2(n5434), 
	.C1(n5491), 
	.B2(n5432), 
	.B1(n5490), 
	.A2(n5430), 
	.A1(n5489));
   OAI222_X1 U4428 (.ZN(\UUT/branch_regb [1]), 
	.C2(n5434), 
	.C1(n5494), 
	.B2(n5432), 
	.B1(n5493), 
	.A2(n5430), 
	.A1(FE_OFN188_n5492));
   OAI222_X1 U4429 (.ZN(\UUT/branch_regb [19]), 
	.C2(n5434), 
	.C1(n5497), 
	.B2(n5432), 
	.B1(n5496), 
	.A2(n5430), 
	.A1(n5495));
   OAI222_X1 U4430 (.ZN(\UUT/branch_regb [18]), 
	.C2(n5434), 
	.C1(n5500), 
	.B2(n5432), 
	.B1(n5499), 
	.A2(n5430), 
	.A1(n5498));
   OAI222_X1 U4431 (.ZN(\UUT/branch_regb [17]), 
	.C2(n5434), 
	.C1(n5503), 
	.B2(n5432), 
	.B1(n5502), 
	.A2(n5430), 
	.A1(n5501));
   OAI222_X1 U4432 (.ZN(\UUT/branch_regb [16]), 
	.C2(n5434), 
	.C1(n5506), 
	.B2(n5432), 
	.B1(n5505), 
	.A2(n5430), 
	.A1(n5504));
   OAI222_X1 U4433 (.ZN(\UUT/branch_regb [15]), 
	.C2(n5434), 
	.C1(n5509), 
	.B2(n5432), 
	.B1(n5508), 
	.A2(n5430), 
	.A1(n5507));
   OAI222_X1 U4434 (.ZN(\UUT/branch_regb [14]), 
	.C2(n5434), 
	.C1(n5512), 
	.B2(n5432), 
	.B1(n5511), 
	.A2(n5430), 
	.A1(n5510));
   OAI222_X1 U4435 (.ZN(\UUT/branch_regb [13]), 
	.C2(n5434), 
	.C1(n5515), 
	.B2(n5432), 
	.B1(n5514), 
	.A2(n5430), 
	.A1(n5513));
   OAI222_X1 U4436 (.ZN(\UUT/branch_regb [12]), 
	.C2(n5434), 
	.C1(n5518), 
	.B2(n5432), 
	.B1(n5517), 
	.A2(n5430), 
	.A1(n5516));
   OAI222_X1 U4437 (.ZN(\UUT/branch_regb [11]), 
	.C2(n5434), 
	.C1(n5521), 
	.B2(n5432), 
	.B1(n5520), 
	.A2(n5430), 
	.A1(n5519));
   OAI222_X1 U4438 (.ZN(\UUT/branch_regb [10]), 
	.C2(n5434), 
	.C1(n5524), 
	.B2(n5432), 
	.B1(n5523), 
	.A2(n5430), 
	.A1(FE_OFN193_n5522));
   OAI222_X1 U4439 (.ZN(\UUT/branch_regb [0]), 
	.C2(n5434), 
	.C1(n5527), 
	.B2(n5432), 
	.B1(n5526), 
	.A2(n5430), 
	.A1(n5525));
   AOI22_X1 U4444 (.ZN(n5533), 
	.B2(\UUT/regfile/reg_out[18][30] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][30] ), 
	.A1(n5534));
   AOI22_X1 U4445 (.ZN(n5538), 
	.B2(\UUT/regfile/reg_out[20][30] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][30] ), 
	.A1(n5539));
   AOI22_X1 U4446 (.ZN(n5543), 
	.B2(\UUT/regfile/reg_out[24][30] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][30] ), 
	.A1(n5544));
   AOI22_X1 U4447 (.ZN(n5548), 
	.B2(\UUT/regfile/reg_out[28][30] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][30] ), 
	.A1(n5549));
   AOI22_X1 U4448 (.ZN(n5555), 
	.B2(\UUT/regfile/reg_out[4][30] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][30] ), 
	.A1(n6376));
   AOI22_X1 U4451 (.ZN(n5565), 
	.B2(\UUT/regfile/reg_out[18][29] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][29] ), 
	.A1(n5534));
   AOI22_X1 U4452 (.ZN(n5566), 
	.B2(\UUT/regfile/reg_out[20][29] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][29] ), 
	.A1(n5539));
   AOI22_X1 U4453 (.ZN(n5567), 
	.B2(\UUT/regfile/reg_out[24][29] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][29] ), 
	.A1(n5544));
   AOI22_X1 U4454 (.ZN(n5568), 
	.B2(\UUT/regfile/reg_out[28][29] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][29] ), 
	.A1(n5549));
   AOI22_X1 U4455 (.ZN(n5569), 
	.B2(\UUT/regfile/reg_out[4][29] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][29] ), 
	.A1(n6376));
   AOI22_X1 U4458 (.ZN(n5572), 
	.B2(\UUT/regfile/reg_out[18][28] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][28] ), 
	.A1(n5534));
   AOI22_X1 U4459 (.ZN(n5573), 
	.B2(\UUT/regfile/reg_out[20][28] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][28] ), 
	.A1(n5539));
   AOI22_X1 U4460 (.ZN(n5574), 
	.B2(\UUT/regfile/reg_out[24][28] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][28] ), 
	.A1(n5544));
   AOI22_X1 U4461 (.ZN(n5575), 
	.B2(\UUT/regfile/reg_out[28][28] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][28] ), 
	.A1(n5549));
   AOI22_X1 U4462 (.ZN(n5576), 
	.B2(\UUT/regfile/reg_out[4][28] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][28] ), 
	.A1(n6375));
   AOI22_X1 U4465 (.ZN(n5579), 
	.B2(\UUT/regfile/reg_out[18][27] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][27] ), 
	.A1(n5534));
   AOI22_X1 U4466 (.ZN(n5580), 
	.B2(\UUT/regfile/reg_out[20][27] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][27] ), 
	.A1(n5539));
   AOI22_X1 U4467 (.ZN(n5581), 
	.B2(\UUT/regfile/reg_out[24][27] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][27] ), 
	.A1(n5544));
   AOI22_X1 U4468 (.ZN(n5582), 
	.B2(\UUT/regfile/reg_out[28][27] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][27] ), 
	.A1(n5549));
   AOI22_X1 U4469 (.ZN(n5583), 
	.B2(\UUT/regfile/reg_out[4][27] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][27] ), 
	.A1(n6375));
   AOI22_X1 U4472 (.ZN(n5586), 
	.B2(\UUT/regfile/reg_out[18][26] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][26] ), 
	.A1(n5534));
   AOI22_X1 U4473 (.ZN(n5587), 
	.B2(\UUT/regfile/reg_out[20][26] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][26] ), 
	.A1(n5539));
   AOI22_X1 U4474 (.ZN(n5588), 
	.B2(\UUT/regfile/reg_out[24][26] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][26] ), 
	.A1(n5544));
   AOI22_X1 U4475 (.ZN(n5589), 
	.B2(\UUT/regfile/reg_out[28][26] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][26] ), 
	.A1(n5549));
   AOI22_X1 U4476 (.ZN(n5590), 
	.B2(\UUT/regfile/reg_out[4][26] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][26] ), 
	.A1(n6376));
   AOI22_X1 U4479 (.ZN(n5593), 
	.B2(\UUT/regfile/reg_out[18][25] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][25] ), 
	.A1(n5534));
   AOI22_X1 U4480 (.ZN(n5594), 
	.B2(\UUT/regfile/reg_out[20][25] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][25] ), 
	.A1(n5539));
   AOI22_X1 U4481 (.ZN(n5595), 
	.B2(\UUT/regfile/reg_out[24][25] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][25] ), 
	.A1(n5544));
   AOI22_X1 U4482 (.ZN(n5596), 
	.B2(\UUT/regfile/reg_out[28][25] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][25] ), 
	.A1(n5549));
   AOI22_X1 U4483 (.ZN(n5597), 
	.B2(\UUT/regfile/reg_out[4][25] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][25] ), 
	.A1(n6375));
   AOI22_X1 U4484 (.ZN(n5474), 
	.B2(n5564), 
	.B1(n5599), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5598));
   AOI22_X1 U4486 (.ZN(n5600), 
	.B2(\UUT/regfile/reg_out[18][24] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][24] ), 
	.A1(n5534));
   AOI22_X1 U4487 (.ZN(n5601), 
	.B2(\UUT/regfile/reg_out[20][24] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][24] ), 
	.A1(n5539));
   AOI22_X1 U4488 (.ZN(n5602), 
	.B2(\UUT/regfile/reg_out[24][24] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][24] ), 
	.A1(n5544));
   AOI22_X1 U4489 (.ZN(n5603), 
	.B2(\UUT/regfile/reg_out[28][24] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][24] ), 
	.A1(n5549));
   AOI22_X1 U4490 (.ZN(n5604), 
	.B2(\UUT/regfile/reg_out[4][24] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][24] ), 
	.A1(n6376));
   AOI22_X1 U4491 (.ZN(n5477), 
	.B2(n5564), 
	.B1(n5606), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5605));
   OAI222_X1 U4492 (.ZN(\UUT/branch_rega [0]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5527), 
	.B2(FE_OFN97_n5529), 
	.B1(n5422), 
	.A2(n5528), 
	.A1(n5525));
   AOI22_X1 U4493 (.ZN(n5607), 
	.B2(\UUT/regfile/reg_out[18][0] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][0] ), 
	.A1(n5534));
   AOI22_X1 U4494 (.ZN(n5608), 
	.B2(\UUT/regfile/reg_out[20][0] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][0] ), 
	.A1(n5539));
   AOI22_X1 U4495 (.ZN(n5609), 
	.B2(\UUT/regfile/reg_out[24][0] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][0] ), 
	.A1(n5544));
   AOI22_X1 U4496 (.ZN(n5610), 
	.B2(\UUT/regfile/reg_out[28][0] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][0] ), 
	.A1(n5549));
   AOI22_X1 U4497 (.ZN(n5611), 
	.B2(\UUT/regfile/reg_out[4][0] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][0] ), 
	.A1(n6375));
   AOI222_X1 U4498 (.ZN(n5525), 
	.C2(\UUT/Mpath/N119 ), 
	.C1(n5613), 
	.B2(n5612), 
	.B1(\UUT/Mpath/out_jar[0] ), 
	.A2(n5564), 
	.A1(\UUT/daddr_out [0]));
   AOI22_X1 U4499 (.ZN(n5718), 
	.B2(\UUT/regfile/reg_out[18][9] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][9] ), 
	.A1(n5719));
   AOI22_X1 U4500 (.ZN(n5723), 
	.B2(\UUT/regfile/reg_out[20][9] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][9] ), 
	.A1(n5724));
   AOI22_X1 U4501 (.ZN(n5728), 
	.B2(\UUT/regfile/reg_out[24][9] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][9] ), 
	.A1(n5729));
   AOI22_X1 U4502 (.ZN(n5733), 
	.B2(\UUT/regfile/reg_out[28][9] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][9] ), 
	.A1(n5734));
   AOI22_X1 U4503 (.ZN(n5740), 
	.B2(\UUT/regfile/reg_out[4][9] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][9] ), 
	.A1(n5741));
   AOI22_X1 U4504 (.ZN(n5749), 
	.B2(\UUT/regfile/reg_out[18][8] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][8] ), 
	.A1(n5719));
   AOI22_X1 U4505 (.ZN(n5750), 
	.B2(\UUT/regfile/reg_out[20][8] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][8] ), 
	.A1(n5724));
   AOI22_X1 U4506 (.ZN(n5751), 
	.B2(\UUT/regfile/reg_out[24][8] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][8] ), 
	.A1(n5729));
   AOI22_X1 U4507 (.ZN(n5752), 
	.B2(\UUT/regfile/reg_out[28][8] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][8] ), 
	.A1(n5734));
   AOI22_X1 U4508 (.ZN(n5753), 
	.B2(\UUT/regfile/reg_out[4][8] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][8] ), 
	.A1(n5741));
   OAI22_X1 U4509 (.ZN(n5759), 
	.B2(n5763), 
	.B1(n5762), 
	.A2(n5761), 
	.A1(n5760));
   AOI22_X1 U4510 (.ZN(n5764), 
	.B2(\UUT/regfile/reg_out[18][7] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][7] ), 
	.A1(n5719));
   AOI22_X1 U4511 (.ZN(n5765), 
	.B2(\UUT/regfile/reg_out[20][7] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][7] ), 
	.A1(n5724));
   AOI22_X1 U4512 (.ZN(n5766), 
	.B2(\UUT/regfile/reg_out[24][7] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][7] ), 
	.A1(n5729));
   AOI22_X1 U4513 (.ZN(n5767), 
	.B2(\UUT/regfile/reg_out[28][7] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][7] ), 
	.A1(n5734));
   AOI22_X1 U4514 (.ZN(n5768), 
	.B2(\UUT/regfile/reg_out[4][7] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][7] ), 
	.A1(n5741));
   OAI22_X1 U4515 (.ZN(n5771), 
	.B2(n5773), 
	.B1(n5763), 
	.A2(n5772), 
	.A1(n5761));
   OAI22_X1 U4516 (.ZN(n5775), 
	.B2(n5778), 
	.B1(n5773), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5776));
   AOI22_X1 U4517 (.ZN(n5773), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[6]), 
	.A2(n5779), 
	.A1(dram_data_inbus[6]));
   INV_X1 U4518 (.ZN(n5774), 
	.A(n5772));
   AOI22_X1 U4519 (.ZN(n5781), 
	.B2(\UUT/regfile/reg_out[18][6] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][6] ), 
	.A1(n5719));
   AOI22_X1 U4520 (.ZN(n5782), 
	.B2(\UUT/regfile/reg_out[20][6] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][6] ), 
	.A1(n5724));
   AOI22_X1 U4521 (.ZN(n5783), 
	.B2(\UUT/regfile/reg_out[24][6] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][6] ), 
	.A1(n5729));
   AOI22_X1 U4522 (.ZN(n5784), 
	.B2(\UUT/regfile/reg_out[28][6] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][6] ), 
	.A1(n5734));
   AOI22_X1 U4523 (.ZN(n5785), 
	.B2(\UUT/regfile/reg_out[4][6] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][6] ), 
	.A1(n5741));
   OAI22_X1 U4524 (.ZN(n5788), 
	.B2(n5790), 
	.B1(n5763), 
	.A2(n5789), 
	.A1(n5761));
   OAI22_X1 U4525 (.ZN(n5792), 
	.B2(n5778), 
	.B1(n5790), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5793));
   AOI22_X1 U4526 (.ZN(n5790), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[5]), 
	.A2(n5779), 
	.A1(dram_data_inbus[5]));
   INV_X1 U4527 (.ZN(n5791), 
	.A(n5789));
   AOI22_X1 U4528 (.ZN(n5794), 
	.B2(\UUT/regfile/reg_out[18][5] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][5] ), 
	.A1(n5719));
   AOI22_X1 U4529 (.ZN(n5795), 
	.B2(\UUT/regfile/reg_out[20][5] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][5] ), 
	.A1(n5724));
   AOI22_X1 U4530 (.ZN(n5796), 
	.B2(\UUT/regfile/reg_out[24][5] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][5] ), 
	.A1(n5729));
   AOI22_X1 U4531 (.ZN(n5797), 
	.B2(\UUT/regfile/reg_out[28][5] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][5] ), 
	.A1(n5734));
   AOI22_X1 U4532 (.ZN(n5798), 
	.B2(\UUT/regfile/reg_out[4][5] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][5] ), 
	.A1(n5741));
   OAI22_X1 U4533 (.ZN(n5801), 
	.B2(n5803), 
	.B1(n5763), 
	.A2(n5802), 
	.A1(n5761));
   OAI22_X1 U4534 (.ZN(n5805), 
	.B2(n5778), 
	.B1(n5803), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5806));
   AOI22_X1 U4535 (.ZN(n5803), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[4]), 
	.A2(n5779), 
	.A1(dram_data_inbus[4]));
   INV_X1 U4536 (.ZN(n5804), 
	.A(n5802));
   AOI22_X1 U4537 (.ZN(n5807), 
	.B2(\UUT/regfile/reg_out[18][4] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][4] ), 
	.A1(n5719));
   AOI22_X1 U4538 (.ZN(n5808), 
	.B2(\UUT/regfile/reg_out[20][4] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][4] ), 
	.A1(n5724));
   AOI22_X1 U4539 (.ZN(n5809), 
	.B2(\UUT/regfile/reg_out[24][4] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][4] ), 
	.A1(n5729));
   AOI22_X1 U4540 (.ZN(n5810), 
	.B2(\UUT/regfile/reg_out[28][4] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][4] ), 
	.A1(n5734));
   AOI22_X1 U4541 (.ZN(n5811), 
	.B2(\UUT/regfile/reg_out[4][4] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][4] ), 
	.A1(n5741));
   OAI22_X1 U4542 (.ZN(n5814), 
	.B2(n5816), 
	.B1(n5763), 
	.A2(n5815), 
	.A1(n5761));
   OAI22_X1 U4543 (.ZN(n5818), 
	.B2(n5778), 
	.B1(n5816), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5819));
   AOI22_X1 U4544 (.ZN(n5816), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[3]), 
	.A2(n5779), 
	.A1(dram_data_inbus[3]));
   INV_X1 U4545 (.ZN(n5817), 
	.A(n5815));
   AOI22_X1 U4546 (.ZN(n5820), 
	.B2(\UUT/regfile/reg_out[18][3] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][3] ), 
	.A1(n5719));
   AOI22_X1 U4547 (.ZN(n5821), 
	.B2(\UUT/regfile/reg_out[20][3] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][3] ), 
	.A1(n5724));
   AOI22_X1 U4548 (.ZN(n5822), 
	.B2(\UUT/regfile/reg_out[24][3] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][3] ), 
	.A1(n5729));
   AOI22_X1 U4549 (.ZN(n5823), 
	.B2(\UUT/regfile/reg_out[28][3] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][3] ), 
	.A1(n5734));
   AOI22_X1 U4550 (.ZN(n5824), 
	.B2(\UUT/regfile/reg_out[4][3] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][3] ), 
	.A1(n5741));
   AOI22_X1 U4551 (.ZN(n5826), 
	.B2(\UUT/regfile/reg_out[18][31] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][31] ), 
	.A1(n5719));
   AOI22_X1 U4552 (.ZN(n5827), 
	.B2(\UUT/regfile/reg_out[20][31] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][31] ), 
	.A1(n5724));
   AOI22_X1 U4553 (.ZN(n5828), 
	.B2(\UUT/regfile/reg_out[24][31] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][31] ), 
	.A1(n5729));
   AOI22_X1 U4554 (.ZN(n5829), 
	.B2(\UUT/regfile/reg_out[28][31] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][31] ), 
	.A1(n5734));
   AOI22_X1 U4555 (.ZN(n5830), 
	.B2(\UUT/regfile/reg_out[4][31] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][31] ), 
	.A1(n5741));
   AOI22_X1 U4556 (.ZN(n5833), 
	.B2(\UUT/regfile/reg_out[18][30] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][30] ), 
	.A1(n5719));
   AOI22_X1 U4557 (.ZN(n5834), 
	.B2(\UUT/regfile/reg_out[20][30] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][30] ), 
	.A1(n5724));
   AOI22_X1 U4558 (.ZN(n5835), 
	.B2(\UUT/regfile/reg_out[24][30] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][30] ), 
	.A1(n5729));
   AOI22_X1 U4559 (.ZN(n5836), 
	.B2(\UUT/regfile/reg_out[28][30] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][30] ), 
	.A1(n5734));
   AOI22_X1 U4560 (.ZN(n5837), 
	.B2(\UUT/regfile/reg_out[4][30] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][30] ), 
	.A1(n5741));
   OAI22_X1 U4561 (.ZN(n5840), 
	.B2(n5842), 
	.B1(n5763), 
	.A2(n5841), 
	.A1(n5761));
   OAI22_X1 U4562 (.ZN(n5844), 
	.B2(n5778), 
	.B1(n5842), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5845));
   AOI22_X1 U4563 (.ZN(n5842), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[2]), 
	.A2(n5779), 
	.A1(dram_data_inbus[2]));
   INV_X1 U4564 (.ZN(n5843), 
	.A(n5841));
   AOI22_X1 U4565 (.ZN(n5846), 
	.B2(\UUT/regfile/reg_out[18][2] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][2] ), 
	.A1(n5719));
   AOI22_X1 U4566 (.ZN(n5847), 
	.B2(\UUT/regfile/reg_out[20][2] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][2] ), 
	.A1(n5724));
   AOI22_X1 U4567 (.ZN(n5848), 
	.B2(\UUT/regfile/reg_out[24][2] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][2] ), 
	.A1(n5729));
   AOI22_X1 U4568 (.ZN(n5849), 
	.B2(\UUT/regfile/reg_out[28][2] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][2] ), 
	.A1(n5734));
   AOI22_X1 U4569 (.ZN(n5850), 
	.B2(\UUT/regfile/reg_out[4][2] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][2] ), 
	.A1(n5741));
   AOI22_X1 U4570 (.ZN(n5852), 
	.B2(\UUT/regfile/reg_out[18][29] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][29] ), 
	.A1(n5719));
   AOI22_X1 U4571 (.ZN(n5853), 
	.B2(\UUT/regfile/reg_out[20][29] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][29] ), 
	.A1(n5724));
   AOI22_X1 U4572 (.ZN(n5854), 
	.B2(\UUT/regfile/reg_out[24][29] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][29] ), 
	.A1(n5729));
   AOI22_X1 U4573 (.ZN(n5855), 
	.B2(\UUT/regfile/reg_out[28][29] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][29] ), 
	.A1(n5734));
   AOI22_X1 U4574 (.ZN(n5856), 
	.B2(\UUT/regfile/reg_out[4][29] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][29] ), 
	.A1(n5741));
   AOI22_X1 U4575 (.ZN(n5858), 
	.B2(\UUT/regfile/reg_out[18][28] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][28] ), 
	.A1(n5719));
   AOI22_X1 U4576 (.ZN(n5859), 
	.B2(\UUT/regfile/reg_out[20][28] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][28] ), 
	.A1(n5724));
   AOI22_X1 U4577 (.ZN(n5860), 
	.B2(\UUT/regfile/reg_out[24][28] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][28] ), 
	.A1(n5729));
   AOI22_X1 U4578 (.ZN(n5861), 
	.B2(\UUT/regfile/reg_out[28][28] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][28] ), 
	.A1(n5734));
   AOI22_X1 U4579 (.ZN(n5862), 
	.B2(\UUT/regfile/reg_out[4][28] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][28] ), 
	.A1(n5741));
   AOI22_X1 U4580 (.ZN(n5864), 
	.B2(\UUT/regfile/reg_out[18][27] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][27] ), 
	.A1(n5719));
   AOI22_X1 U4581 (.ZN(n5865), 
	.B2(\UUT/regfile/reg_out[20][27] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][27] ), 
	.A1(n5724));
   AOI22_X1 U4582 (.ZN(n5866), 
	.B2(\UUT/regfile/reg_out[24][27] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][27] ), 
	.A1(n5729));
   AOI22_X1 U4583 (.ZN(n5867), 
	.B2(\UUT/regfile/reg_out[28][27] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][27] ), 
	.A1(n5734));
   AOI22_X1 U4584 (.ZN(n5868), 
	.B2(\UUT/regfile/reg_out[4][27] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][27] ), 
	.A1(n5741));
   NOR2_X1 U4585 (.ZN(n5869), 
	.A2(n5872), 
	.A1(n5871));
   AOI22_X1 U4586 (.ZN(n5874), 
	.B2(\UUT/regfile/reg_out[18][26] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][26] ), 
	.A1(n5719));
   AOI22_X1 U4587 (.ZN(n5875), 
	.B2(\UUT/regfile/reg_out[20][26] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][26] ), 
	.A1(n5724));
   AOI22_X1 U4588 (.ZN(n5876), 
	.B2(\UUT/regfile/reg_out[24][26] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][26] ), 
	.A1(n5729));
   AOI22_X1 U4589 (.ZN(n5877), 
	.B2(\UUT/regfile/reg_out[28][26] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][26] ), 
	.A1(n5734));
   AOI22_X1 U4590 (.ZN(n5878), 
	.B2(\UUT/regfile/reg_out[4][26] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][26] ), 
	.A1(n5741));
   AOI22_X1 U4591 (.ZN(n5883), 
	.B2(\UUT/regfile/reg_out[18][25] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][25] ), 
	.A1(n5719));
   AOI22_X1 U4592 (.ZN(n5884), 
	.B2(\UUT/regfile/reg_out[20][25] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][25] ), 
	.A1(n5724));
   AOI22_X1 U4593 (.ZN(n5885), 
	.B2(\UUT/regfile/reg_out[24][25] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][25] ), 
	.A1(n5729));
   AOI22_X1 U4594 (.ZN(n5886), 
	.B2(\UUT/regfile/reg_out[28][25] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][25] ), 
	.A1(n5734));
   AOI22_X1 U4595 (.ZN(n5887), 
	.B2(\UUT/regfile/reg_out[4][25] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][25] ), 
	.A1(n5741));
   AOI22_X1 U4596 (.ZN(n5891), 
	.B2(\UUT/regfile/reg_out[18][24] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][24] ), 
	.A1(n5719));
   AOI22_X1 U4597 (.ZN(n5892), 
	.B2(\UUT/regfile/reg_out[20][24] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][24] ), 
	.A1(n5724));
   AOI22_X1 U4598 (.ZN(n5893), 
	.B2(\UUT/regfile/reg_out[24][24] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][24] ), 
	.A1(n5729));
   AOI22_X1 U4599 (.ZN(n5894), 
	.B2(\UUT/regfile/reg_out[28][24] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][24] ), 
	.A1(n5734));
   AOI22_X1 U4600 (.ZN(n5895), 
	.B2(\UUT/regfile/reg_out[4][24] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][24] ), 
	.A1(n5741));
   AOI22_X1 U4601 (.ZN(n5898), 
	.B2(\UUT/regfile/reg_out[18][23] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][23] ), 
	.A1(n5719));
   AOI22_X1 U4602 (.ZN(n5899), 
	.B2(\UUT/regfile/reg_out[20][23] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][23] ), 
	.A1(n5724));
   AOI22_X1 U4603 (.ZN(n5900), 
	.B2(\UUT/regfile/reg_out[24][23] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][23] ), 
	.A1(n5729));
   AOI22_X1 U4604 (.ZN(n5901), 
	.B2(\UUT/regfile/reg_out[28][23] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][23] ), 
	.A1(n5734));
   AOI22_X1 U4605 (.ZN(n5902), 
	.B2(\UUT/regfile/reg_out[4][23] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][23] ), 
	.A1(n5741));
   AOI22_X1 U4606 (.ZN(n5903), 
	.B2(\UUT/regfile/reg_out[18][22] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][22] ), 
	.A1(n5719));
   AOI22_X1 U4607 (.ZN(n5904), 
	.B2(\UUT/regfile/reg_out[20][22] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][22] ), 
	.A1(n5724));
   AOI22_X1 U4608 (.ZN(n5905), 
	.B2(\UUT/regfile/reg_out[24][22] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][22] ), 
	.A1(n5729));
   AOI22_X1 U4609 (.ZN(n5906), 
	.B2(\UUT/regfile/reg_out[28][22] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][22] ), 
	.A1(n5734));
   AOI22_X1 U4610 (.ZN(n5907), 
	.B2(\UUT/regfile/reg_out[4][22] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][22] ), 
	.A1(n5741));
   AOI22_X1 U4611 (.ZN(n5908), 
	.B2(\UUT/regfile/reg_out[18][21] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][21] ), 
	.A1(n5719));
   AOI22_X1 U4612 (.ZN(n5909), 
	.B2(\UUT/regfile/reg_out[20][21] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][21] ), 
	.A1(n5724));
   AOI22_X1 U4613 (.ZN(n5910), 
	.B2(\UUT/regfile/reg_out[24][21] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][21] ), 
	.A1(n5729));
   AOI22_X1 U4614 (.ZN(n5911), 
	.B2(\UUT/regfile/reg_out[28][21] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][21] ), 
	.A1(n5734));
   AOI22_X1 U4615 (.ZN(n5912), 
	.B2(\UUT/regfile/reg_out[4][21] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][21] ), 
	.A1(n5741));
   AOI22_X1 U4616 (.ZN(n5913), 
	.B2(\UUT/regfile/reg_out[18][20] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][20] ), 
	.A1(n5719));
   AOI22_X1 U4617 (.ZN(n5914), 
	.B2(\UUT/regfile/reg_out[20][20] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][20] ), 
	.A1(n5724));
   AOI22_X1 U4618 (.ZN(n5915), 
	.B2(\UUT/regfile/reg_out[24][20] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][20] ), 
	.A1(n5729));
   AOI22_X1 U4619 (.ZN(n5916), 
	.B2(\UUT/regfile/reg_out[28][20] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][20] ), 
	.A1(n5734));
   AOI22_X1 U4620 (.ZN(n5917), 
	.B2(\UUT/regfile/reg_out[4][20] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][20] ), 
	.A1(n5741));
   OAI22_X1 U4621 (.ZN(n5918), 
	.B2(n5920), 
	.B1(n5763), 
	.A2(n5919), 
	.A1(n5761));
   OAI22_X1 U4623 (.ZN(n5923), 
	.B2(n5778), 
	.B1(n5920), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5921));
   AOI22_X1 U4624 (.ZN(n5920), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[1]), 
	.A2(n5779), 
	.A1(dram_data_inbus[1]));
   AOI22_X1 U4625 (.ZN(n5921), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[9]), 
	.A2(n5779), 
	.A1(dram_data_inbus[9]));
   INV_X1 U4626 (.ZN(n5712), 
	.A(n5882));
   INV_X1 U4627 (.ZN(n5922), 
	.A(n5919));
   AOI22_X1 U4628 (.ZN(n5924), 
	.B2(\UUT/regfile/reg_out[18][1] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][1] ), 
	.A1(n5719));
   AOI22_X1 U4629 (.ZN(n5925), 
	.B2(\UUT/regfile/reg_out[20][1] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][1] ), 
	.A1(n5724));
   AOI22_X1 U4630 (.ZN(n5926), 
	.B2(\UUT/regfile/reg_out[24][1] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][1] ), 
	.A1(n5729));
   AOI22_X1 U4631 (.ZN(n5927), 
	.B2(\UUT/regfile/reg_out[28][1] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][1] ), 
	.A1(n5734));
   AOI22_X1 U4632 (.ZN(n5928), 
	.B2(\UUT/regfile/reg_out[4][1] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][1] ), 
	.A1(n5741));
   AOI22_X1 U4633 (.ZN(n5929), 
	.B2(\UUT/regfile/reg_out[18][19] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][19] ), 
	.A1(n5719));
   AOI22_X1 U4634 (.ZN(n5930), 
	.B2(\UUT/regfile/reg_out[20][19] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][19] ), 
	.A1(n5724));
   AOI22_X1 U4635 (.ZN(n5931), 
	.B2(\UUT/regfile/reg_out[24][19] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][19] ), 
	.A1(n5729));
   AOI22_X1 U4636 (.ZN(n5932), 
	.B2(\UUT/regfile/reg_out[28][19] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][19] ), 
	.A1(n5734));
   AOI22_X1 U4637 (.ZN(n5933), 
	.B2(\UUT/regfile/reg_out[4][19] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][19] ), 
	.A1(n5741));
   AOI22_X1 U4638 (.ZN(n5934), 
	.B2(\UUT/regfile/reg_out[18][18] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][18] ), 
	.A1(n5719));
   AOI22_X1 U4639 (.ZN(n5935), 
	.B2(\UUT/regfile/reg_out[20][18] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][18] ), 
	.A1(n5724));
   AOI22_X1 U4640 (.ZN(n5936), 
	.B2(\UUT/regfile/reg_out[24][18] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][18] ), 
	.A1(n5729));
   AOI22_X1 U4641 (.ZN(n5937), 
	.B2(\UUT/regfile/reg_out[28][18] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][18] ), 
	.A1(n5734));
   AOI22_X1 U4642 (.ZN(n5938), 
	.B2(\UUT/regfile/reg_out[4][18] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][18] ), 
	.A1(n5741));
   AOI22_X1 U4643 (.ZN(n5939), 
	.B2(\UUT/regfile/reg_out[18][17] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][17] ), 
	.A1(n5719));
   AOI22_X1 U4644 (.ZN(n5940), 
	.B2(\UUT/regfile/reg_out[20][17] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][17] ), 
	.A1(n5724));
   AOI22_X1 U4645 (.ZN(n5941), 
	.B2(\UUT/regfile/reg_out[24][17] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][17] ), 
	.A1(n5729));
   AOI22_X1 U4646 (.ZN(n5942), 
	.B2(\UUT/regfile/reg_out[28][17] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][17] ), 
	.A1(n5734));
   AOI22_X1 U4647 (.ZN(n5943), 
	.B2(\UUT/regfile/reg_out[4][17] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][17] ), 
	.A1(n5741));
   NOR3_X1 U4648 (.ZN(n5945), 
	.A3(n5948), 
	.A2(n5947), 
	.A1(n5946));
   AOI22_X1 U4649 (.ZN(n5947), 
	.B2(n5756), 
	.B1(\UUT/Mpath/the_memhandle/N239 ), 
	.A2(n5949), 
	.A1(n487));
   INV_X1 U4650 (.ZN(n5946), 
	.A(\UUT/Mpath/the_memhandle/N86 ));
   AOI22_X1 U4651 (.ZN(n5952), 
	.B2(\UUT/regfile/reg_out[18][16] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][16] ), 
	.A1(n5719));
   AOI22_X1 U4652 (.ZN(n5953), 
	.B2(\UUT/regfile/reg_out[20][16] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][16] ), 
	.A1(n5724));
   AOI22_X1 U4653 (.ZN(n5954), 
	.B2(\UUT/regfile/reg_out[24][16] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][16] ), 
	.A1(n5729));
   AOI22_X1 U4654 (.ZN(n5955), 
	.B2(\UUT/regfile/reg_out[28][16] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][16] ), 
	.A1(n5734));
   AOI22_X1 U4655 (.ZN(n5956), 
	.B2(\UUT/regfile/reg_out[4][16] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][16] ), 
	.A1(n5741));
   INV_X1 U4657 (.ZN(n5756), 
	.A(n5825));
   AOI22_X1 U4658 (.ZN(n5958), 
	.B2(\UUT/regfile/reg_out[18][15] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][15] ), 
	.A1(n5719));
   AOI22_X1 U4659 (.ZN(n5959), 
	.B2(\UUT/regfile/reg_out[20][15] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][15] ), 
	.A1(n5724));
   AOI22_X1 U4660 (.ZN(n5960), 
	.B2(\UUT/regfile/reg_out[24][15] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][15] ), 
	.A1(n5729));
   AOI22_X1 U4661 (.ZN(n5961), 
	.B2(\UUT/regfile/reg_out[28][15] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][15] ), 
	.A1(n5734));
   AOI22_X1 U4662 (.ZN(n5962), 
	.B2(\UUT/regfile/reg_out[4][15] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][15] ), 
	.A1(n5741));
   AOI22_X1 U4664 (.ZN(n5776), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[14]), 
	.A2(n5779), 
	.A1(dram_data_inbus[14]));
   INV_X1 U4665 (.ZN(n5769), 
	.A(n5832));
   AOI22_X1 U4666 (.ZN(n5963), 
	.B2(\UUT/regfile/reg_out[18][14] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][14] ), 
	.A1(n5719));
   AOI22_X1 U4667 (.ZN(n5964), 
	.B2(\UUT/regfile/reg_out[20][14] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][14] ), 
	.A1(n5724));
   AOI22_X1 U4668 (.ZN(n5965), 
	.B2(\UUT/regfile/reg_out[24][14] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][14] ), 
	.A1(n5729));
   AOI22_X1 U4669 (.ZN(n5966), 
	.B2(\UUT/regfile/reg_out[28][14] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][14] ), 
	.A1(n5734));
   AOI22_X1 U4670 (.ZN(n5967), 
	.B2(\UUT/regfile/reg_out[4][14] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][14] ), 
	.A1(n5741));
   AOI22_X1 U4672 (.ZN(n5793), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[13]), 
	.A2(n5779), 
	.A1(dram_data_inbus[13]));
   INV_X1 U4673 (.ZN(n5786), 
	.A(n5851));
   AOI22_X1 U4674 (.ZN(n5968), 
	.B2(\UUT/regfile/reg_out[18][13] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][13] ), 
	.A1(n5719));
   AOI22_X1 U4675 (.ZN(n5969), 
	.B2(\UUT/regfile/reg_out[20][13] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][13] ), 
	.A1(n5724));
   AOI22_X1 U4676 (.ZN(n5970), 
	.B2(\UUT/regfile/reg_out[24][13] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][13] ), 
	.A1(n5729));
   AOI22_X1 U4677 (.ZN(n5971), 
	.B2(\UUT/regfile/reg_out[28][13] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][13] ), 
	.A1(n5734));
   AOI22_X1 U4678 (.ZN(n5972), 
	.B2(\UUT/regfile/reg_out[4][13] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][13] ), 
	.A1(n5741));
   AOI22_X1 U4680 (.ZN(n5806), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[12]), 
	.A2(n5779), 
	.A1(dram_data_inbus[12]));
   INV_X1 U4681 (.ZN(n5799), 
	.A(n5857));
   AOI22_X1 U4682 (.ZN(n5973), 
	.B2(\UUT/regfile/reg_out[18][12] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][12] ), 
	.A1(n5719));
   AOI22_X1 U4683 (.ZN(n5974), 
	.B2(\UUT/regfile/reg_out[20][12] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][12] ), 
	.A1(n5724));
   AOI22_X1 U4684 (.ZN(n5975), 
	.B2(\UUT/regfile/reg_out[24][12] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][12] ), 
	.A1(n5729));
   AOI22_X1 U4685 (.ZN(n5976), 
	.B2(\UUT/regfile/reg_out[28][12] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][12] ), 
	.A1(n5734));
   AOI22_X1 U4686 (.ZN(n5977), 
	.B2(\UUT/regfile/reg_out[4][12] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][12] ), 
	.A1(n5741));
   AOI22_X1 U4688 (.ZN(n5819), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[11]), 
	.A2(n5779), 
	.A1(dram_data_inbus[11]));
   INV_X1 U4689 (.ZN(n5812), 
	.A(n5863));
   AOI22_X1 U4690 (.ZN(n5978), 
	.B2(\UUT/regfile/reg_out[18][11] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][11] ), 
	.A1(n5719));
   AOI22_X1 U4691 (.ZN(n5979), 
	.B2(\UUT/regfile/reg_out[20][11] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][11] ), 
	.A1(n5724));
   AOI22_X1 U4692 (.ZN(n5980), 
	.B2(\UUT/regfile/reg_out[24][11] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][11] ), 
	.A1(n5729));
   AOI22_X1 U4693 (.ZN(n5981), 
	.B2(\UUT/regfile/reg_out[28][11] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][11] ), 
	.A1(n5734));
   AOI22_X1 U4694 (.ZN(n5982), 
	.B2(\UUT/regfile/reg_out[4][11] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][11] ), 
	.A1(n5741));
   INV_X1 U4695 (.ZN(n5715), 
	.A(n5754));
   OAI22_X1 U4696 (.ZN(n5984), 
	.B2(n5986), 
	.B1(n5760), 
	.A2(n5985), 
	.A1(n5825));
   INV_X1 U4697 (.ZN(n5986), 
	.A(\UUT/Mpath/the_memhandle/N37 ));
   INV_X1 U4698 (.ZN(n5985), 
	.A(\UUT/Mpath/the_memhandle/N36 ));
   OAI22_X1 U4699 (.ZN(n5983), 
	.B2(n5778), 
	.B1(n5762), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5957));
   AOI22_X1 U4700 (.ZN(n5762), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[7]), 
	.A2(n5779), 
	.A1(dram_data_inbus[7]));
   AOI22_X1 U4701 (.ZN(n5957), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[15]), 
	.A2(n5779), 
	.A1(dram_data_inbus[15]));
   AOI22_X1 U4703 (.ZN(n5845), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[10]), 
	.A2(n5779), 
	.A1(dram_data_inbus[10]));
   NOR2_X1 U4704 (.ZN(n5713), 
	.A2(n5987), 
	.A1(n5948));
   INV_X1 U4705 (.ZN(n5838), 
	.A(n5873));
   NOR2_X1 U4706 (.ZN(n5711), 
	.A2(n5948), 
	.A1(n5988));
   INV_X1 U4707 (.ZN(n5948), 
	.A(n5950));
   NOR2_X1 U4708 (.ZN(n5950), 
	.A2(\UUT/Mpath/the_memhandle/N72 ), 
	.A1(\UUT/Mpath/the_memhandle/N34 ));
   AOI22_X1 U4709 (.ZN(n5989), 
	.B2(\UUT/regfile/reg_out[18][10] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][10] ), 
	.A1(n5719));
   AOI22_X1 U4710 (.ZN(n5990), 
	.B2(\UUT/regfile/reg_out[20][10] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][10] ), 
	.A1(n5724));
   AOI22_X1 U4711 (.ZN(n5991), 
	.B2(\UUT/regfile/reg_out[24][10] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][10] ), 
	.A1(n5729));
   AOI22_X1 U4712 (.ZN(n5992), 
	.B2(\UUT/regfile/reg_out[28][10] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][10] ), 
	.A1(n5734));
   AOI22_X1 U4713 (.ZN(n5993), 
	.B2(\UUT/regfile/reg_out[4][10] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][10] ), 
	.A1(n5741));
   OAI22_X1 U4714 (.ZN(n5994), 
	.B2(n5995), 
	.B1(n5763), 
	.A2(n5944), 
	.A1(n5761));
   AOI21_X1 U4715 (.ZN(n5763), 
	.B2(n5988), 
	.B1(n5996), 
	.A(n5997));
   AND2_X1 U4716 (.ZN(n5997), 
	.A2(\UUT/Mpath/the_memhandle/N72 ), 
	.A1(\UUT/Mpath/the_memhandle/N39 ));
   INV_X1 U4717 (.ZN(n5761), 
	.A(n5998));
   OAI22_X1 U4718 (.ZN(n5998), 
	.B2(n5988), 
	.B1(\UUT/Mpath/the_memhandle/N72 ), 
	.A2(\UUT/Mpath/the_memhandle/N241 ), 
	.A1(n5996));
   INV_X1 U4719 (.ZN(n5988), 
	.A(n5987));
   NOR2_X1 U4720 (.ZN(n5987), 
	.A2(n5951), 
	.A1(n5949));
   NOR2_X1 U4721 (.ZN(n5951), 
	.A2(\UUT/Mpath/the_memhandle/N86 ), 
	.A1(\UUT/Mpath/the_memhandle/N120 ));
   INV_X1 U4722 (.ZN(n5949), 
	.A(\UUT/Mpath/the_memhandle/N239 ));
   INV_X1 U4723 (.ZN(n5996), 
	.A(\UUT/Mpath/the_memhandle/N72 ));
   AND2_X1 U4725 (.ZN(n5757), 
	.A2(\UUT/Mpath/the_memhandle/N72 ), 
	.A1(\UUT/Mpath/the_memhandle/N76 ));
   AND2_X1 U4726 (.ZN(n5755), 
	.A2(\UUT/Mpath/the_memhandle/N72 ), 
	.A1(\UUT/Mpath/the_memhandle/N36 ));
   OAI22_X1 U4727 (.ZN(n6001), 
	.B2(n5778), 
	.B1(n5995), 
	.A2(\UUT/Mpath/the_memhandle/N242 ), 
	.A1(n5999));
   INV_X1 U4728 (.ZN(n5778), 
	.A(\UUT/Mpath/the_memhandle/N39 ));
   AOI22_X1 U4729 (.ZN(n5995), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[0]), 
	.A2(n5779), 
	.A1(dram_data_inbus[0]));
   AOI22_X1 U4731 (.ZN(n5999), 
	.B2(FE_OFN92_n5780), 
	.B1(BUS_DATA_INBUS[8]), 
	.A2(n5779), 
	.A1(dram_data_inbus[8]));
   INV_X1 U4732 (.ZN(n5747), 
	.A(n5890));
   INV_X1 U4733 (.ZN(n6000), 
	.A(n5944));
   NOR3_X1 U4734 (.ZN(n5780), 
	.A3(n6002), 
	.A2(\localbus/c2_op[MASTER] ), 
	.A1(\localbus/N93 ));
   INV_X1 U4735 (.ZN(n6002), 
	.A(\localbus/N95 ));
   INV_X1 U4737 (.ZN(n6003), 
	.A(\localbus/N93 ));
   AOI22_X1 U4738 (.ZN(n6004), 
	.B2(\UUT/regfile/reg_out[18][0] ), 
	.B1(n5720), 
	.A2(\UUT/regfile/reg_out[19][0] ), 
	.A1(n5719));
   AND2_X1 U4743 (.ZN(n6005), 
	.A2(n6010), 
	.A1(n6009));
   AOI22_X1 U4744 (.ZN(n6011), 
	.B2(\UUT/regfile/reg_out[20][0] ), 
	.B1(n5725), 
	.A2(\UUT/regfile/reg_out[21][0] ), 
	.A1(n5724));
   NAND3_X1 U4747 (.ZN(n5722), 
	.A3(n6009), 
	.A2(\UUT/rs2_addr [2]), 
	.A1(n6006));
   NAND4_X1 U4748 (.ZN(n5721), 
	.A4(\UUT/rs2_addr [2]), 
	.A3(\UUT/rs2_addr [0]), 
	.A2(\UUT/rs2_addr [1]), 
	.A1(n6009));
   NOR2_X1 U4749 (.ZN(n6009), 
	.A2(\UUT/rs2_addr [3]), 
	.A1(n6014));
   AOI22_X1 U4750 (.ZN(n6015), 
	.B2(\UUT/regfile/reg_out[24][0] ), 
	.B1(n5730), 
	.A2(\UUT/regfile/reg_out[25][0] ), 
	.A1(n5729));
   NAND3_X1 U4753 (.ZN(n5727), 
	.A3(n6018), 
	.A2(\UUT/rs2_addr [4]), 
	.A1(n6006));
   AOI22_X1 U4755 (.ZN(n6019), 
	.B2(\UUT/regfile/reg_out[28][0] ), 
	.B1(n5735), 
	.A2(\UUT/regfile/reg_out[29][0] ), 
	.A1(n5734));
   NOR2_X1 U4760 (.ZN(n6017), 
	.A2(n6007), 
	.A1(n6014));
   AOI22_X1 U4763 (.ZN(n6024), 
	.B2(\UUT/regfile/reg_out[4][0] ), 
	.B1(n5742), 
	.A2(\UUT/regfile/reg_out[5][0] ), 
	.A1(n5741));
   NAND3_X1 U4766 (.ZN(n5739), 
	.A3(n6023), 
	.A2(n6022), 
	.A1(\UUT/rs2_addr [2]));
   NAND3_X1 U4767 (.ZN(n5738), 
	.A3(n6021), 
	.A2(\UUT/rs2_addr [2]), 
	.A1(\UUT/rs2_addr [1]));
   AND2_X1 U4768 (.ZN(n6021), 
	.A2(n6022), 
	.A1(n6025));
   NOR2_X1 U4771 (.ZN(n6020), 
	.A2(n6010), 
	.A1(n6022));
   AND2_X1 U4772 (.ZN(n6012), 
	.A2(n6007), 
	.A1(n6013));
   INV_X1 U4773 (.ZN(\UUT/rs2_addr [3]), 
	.A(n6022));
   NOR2_X1 U4774 (.ZN(n6013), 
	.A2(\UUT/rs2_addr [1]), 
	.A1(n6010));
   INV_X1 U4775 (.ZN(n6010), 
	.A(\UUT/rs2_addr [2]));
   INV_X1 U4777 (.ZN(\UUT/rs2_addr [1]), 
	.A(n6008));
   AND2_X1 U4779 (.ZN(n6023), 
	.A2(n6014), 
	.A1(n6006));
   NOR2_X1 U4780 (.ZN(n6006), 
	.A2(\UUT/rs2_addr [0]), 
	.A1(n6008));
   AND2_X1 U4781 (.ZN(n6016), 
	.A2(n6008), 
	.A1(n6018));
   NAND2_X1 U4782 (.ZN(n6008), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1871 ), 
	.A1(\UUT/Mcontrol/d_sampled_finstr [17]));
   NOR2_X1 U4783 (.ZN(n6018), 
	.A2(\UUT/rs2_addr [2]), 
	.A1(n6022));
   NAND2_X1 U4784 (.ZN(\UUT/rs2_addr [2]), 
	.A2(n6026), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1871 ));
   NAND2_X1 U4785 (.ZN(n6022), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1871 ), 
	.A1(\UUT/Mcontrol/d_sampled_finstr [19]));
   NOR2_X1 U4786 (.ZN(n6025), 
	.A2(\UUT/rs2_addr [4]), 
	.A1(n6007));
   INV_X1 U4787 (.ZN(\UUT/rs2_addr [4]), 
	.A(n6014));
   NAND2_X1 U4788 (.ZN(n6014), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [20]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1871 ));
   INV_X1 U4789 (.ZN(n6007), 
	.A(\UUT/rs2_addr [0]));
   NAND2_X1 U4790 (.ZN(\UUT/rs2_addr [0]), 
	.A2(n6027), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1871 ));
   AOI21_X1 U4799 (.ZN(n6038), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N1952 ), 
	.B1(n6040), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1964 ));
   NAND4_X1 U4800 (.ZN(n6041), 
	.A4(n6045), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N89 ), 
	.A2(n6044), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1907 ));
   NOR3_X1 U4801 (.ZN(n6044), 
	.A3(n6039), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1970 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1958 ));
   NOR4_X1 U4802 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N255 ), 
	.A4(n6054), 
	.A3(n6053), 
	.A2(n6029), 
	.A1(n6052));
   AOI21_X1 U4803 (.ZN(n6052), 
	.B2(n6046), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N1928 ), 
	.A(n1008));
   OAI21_X1 U4804 (.ZN(\UUT/Mcontrol/d_jump_type[2] ), 
	.B2(n6053), 
	.B1(n6055), 
	.A(n6056));
   AOI21_X1 U4805 (.ZN(n6055), 
	.B2(n6057), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [18]), 
	.A(n6058));
   AOI21_X1 U4806 (.ZN(n6058), 
	.B2(n6060), 
	.B1(n6059), 
	.A(n1008));
   OAI21_X1 U4807 (.ZN(\UUT/Mcontrol/d_jump_type[1] ), 
	.B2(n6053), 
	.B1(n6061), 
	.A(n6056));
   AOI21_X1 U4808 (.ZN(n6061), 
	.B2(n6062), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [17]), 
	.A(n6045));
   OAI21_X1 U4809 (.ZN(\UUT/Mcontrol/d_jump_type[0] ), 
	.B2(n6064), 
	.B1(n6063), 
	.A(n6056));
   AOI221_X1 U4810 (.ZN(n6063), 
	.C2(\UUT/Mcontrol/d_sampled_finstr [16]), 
	.C1(n1008), 
	.B2(n6060), 
	.B1(n6065), 
	.A(n6066));
   INV_X1 U4811 (.ZN(n6060), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1940 ));
   OAI22_X1 U4812 (.ZN(n6065), 
	.B2(n6059), 
	.B1(n1008), 
	.A2(n6067), 
	.A1(n6027));
   NOR2_X1 U4813 (.ZN(n6059), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1934 ), 
	.A1(n6068));
   AOI21_X1 U4814 (.ZN(n6068), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N89 ), 
	.B1(\UUT/Mcontrol/Operation_decoding32/N62 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1928 ));
   INV_X1 U4821 (.ZN(n6075), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2061 ));
   OAI211_X1 U4822 (.ZN(n6077), 
	.C2(n6039), 
	.C1(n6076), 
	.B(n6078), 
	.A(n6051));
   AOI22_X1 U4823 (.ZN(n6080), 
	.B2(\UUT/regfile/reg_out[18][1] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][1] ), 
	.A1(n5534));
   AOI22_X1 U4824 (.ZN(n6081), 
	.B2(\UUT/regfile/reg_out[20][1] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][1] ), 
	.A1(n5539));
   AOI22_X1 U4825 (.ZN(n6082), 
	.B2(\UUT/regfile/reg_out[24][1] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][1] ), 
	.A1(n5544));
   AOI22_X1 U4826 (.ZN(n6083), 
	.B2(\UUT/regfile/reg_out[28][1] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][1] ), 
	.A1(n5549));
   AOI22_X1 U4827 (.ZN(n6084), 
	.B2(\UUT/regfile/reg_out[4][1] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][1] ), 
	.A1(n6376));
   INV_X1 U4828 (.ZN(\UUT/Mcontrol/d_instr [1]), 
	.A(n5427));
   AOI22_X1 U4829 (.ZN(n6087), 
	.B2(\UUT/regfile/reg_out[18][23] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][23] ), 
	.A1(n5534));
   AOI22_X1 U4830 (.ZN(n6088), 
	.B2(\UUT/regfile/reg_out[20][23] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][23] ), 
	.A1(n5539));
   AOI22_X1 U4831 (.ZN(n6089), 
	.B2(\UUT/regfile/reg_out[24][23] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][23] ), 
	.A1(n5544));
   AOI22_X1 U4832 (.ZN(n6090), 
	.B2(\UUT/regfile/reg_out[28][23] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][23] ), 
	.A1(n5549));
   AOI22_X1 U4833 (.ZN(n6091), 
	.B2(\UUT/regfile/reg_out[4][23] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][23] ), 
	.A1(n6375));
   OAI21_X1 U4834 (.ZN(n6093), 
	.B2(n5872), 
	.B1(n6037), 
	.A(n5880));
   INV_X1 U4835 (.ZN(\UUT/Mcontrol/d_instr [7]), 
	.A(n6094));
   AOI22_X1 U4836 (.ZN(n6095), 
	.B2(\UUT/regfile/reg_out[18][22] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][22] ), 
	.A1(n5534));
   AOI22_X1 U4837 (.ZN(n6096), 
	.B2(\UUT/regfile/reg_out[20][22] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][22] ), 
	.A1(n5539));
   AOI22_X1 U4838 (.ZN(n6097), 
	.B2(\UUT/regfile/reg_out[24][22] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][22] ), 
	.A1(n5544));
   AOI22_X1 U4839 (.ZN(n6098), 
	.B2(\UUT/regfile/reg_out[28][22] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][22] ), 
	.A1(n5549));
   AOI22_X1 U4840 (.ZN(n6099), 
	.B2(\UUT/regfile/reg_out[4][22] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][22] ), 
	.A1(n6376));
   OAI21_X1 U4841 (.ZN(n6101), 
	.B2(n5872), 
	.B1(n6029), 
	.A(n5880));
   AOI22_X1 U4842 (.ZN(n6102), 
	.B2(\UUT/regfile/reg_out[18][21] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][21] ), 
	.A1(n5534));
   AOI22_X1 U4843 (.ZN(n6103), 
	.B2(\UUT/regfile/reg_out[20][21] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][21] ), 
	.A1(n5539));
   AOI22_X1 U4844 (.ZN(n6104), 
	.B2(\UUT/regfile/reg_out[24][21] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][21] ), 
	.A1(n5544));
   AOI22_X1 U4845 (.ZN(n6105), 
	.B2(\UUT/regfile/reg_out[28][21] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][21] ), 
	.A1(n5549));
   AOI22_X1 U4846 (.ZN(n6106), 
	.B2(\UUT/regfile/reg_out[4][21] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][21] ), 
	.A1(n6376));
   OAI21_X1 U4847 (.ZN(n6108), 
	.B2(n5872), 
	.B1(n6031), 
	.A(n5880));
   INV_X1 U4848 (.ZN(\UUT/Mcontrol/d_instr [5]), 
	.A(n5423));
   AOI22_X1 U4849 (.ZN(n6109), 
	.B2(\UUT/regfile/reg_out[18][20] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][20] ), 
	.A1(n5534));
   AOI22_X1 U4850 (.ZN(n6110), 
	.B2(\UUT/regfile/reg_out[20][20] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][20] ), 
	.A1(n5539));
   AOI22_X1 U4851 (.ZN(n6111), 
	.B2(\UUT/regfile/reg_out[24][20] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][20] ), 
	.A1(n5544));
   AOI22_X1 U4852 (.ZN(n6112), 
	.B2(\UUT/regfile/reg_out[28][20] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][20] ), 
	.A1(n5549));
   AOI22_X1 U4853 (.ZN(n6113), 
	.B2(\UUT/regfile/reg_out[4][20] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][20] ), 
	.A1(n6376));
   OAI21_X1 U4854 (.ZN(n6115), 
	.B2(n6026), 
	.B1(n5872), 
	.A(n5880));
   OAI21_X1 U4855 (.ZN(n5870), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.B1(n5831), 
	.A(n6117));
   AOI22_X1 U4856 (.ZN(n6119), 
	.B2(\UUT/regfile/reg_out[18][19] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][19] ), 
	.A1(n5534));
   AOI22_X1 U4857 (.ZN(n6120), 
	.B2(\UUT/regfile/reg_out[20][19] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][19] ), 
	.A1(n5539));
   AOI22_X1 U4858 (.ZN(n6121), 
	.B2(\UUT/regfile/reg_out[24][19] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][19] ), 
	.A1(n5544));
   AOI22_X1 U4859 (.ZN(n6122), 
	.B2(\UUT/regfile/reg_out[28][19] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][19] ), 
	.A1(n5549));
   AOI22_X1 U4860 (.ZN(n6123), 
	.B2(\UUT/regfile/reg_out[4][19] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][19] ), 
	.A1(n6375));
   OAI221_X1 U4861 (.ZN(n6126), 
	.C2(n6128), 
	.C1(n5871), 
	.B2(n6118), 
	.B1(n6034), 
	.A(n6117));
   AOI22_X1 U4862 (.ZN(n6129), 
	.B2(\UUT/regfile/reg_out[18][18] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][18] ), 
	.A1(n5534));
   AOI22_X1 U4863 (.ZN(n6130), 
	.B2(\UUT/regfile/reg_out[20][18] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][18] ), 
	.A1(n5539));
   AOI22_X1 U4864 (.ZN(n6131), 
	.B2(\UUT/regfile/reg_out[24][18] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][18] ), 
	.A1(n5544));
   AOI22_X1 U4865 (.ZN(n6132), 
	.B2(\UUT/regfile/reg_out[28][18] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][18] ), 
	.A1(n5549));
   AOI22_X1 U4866 (.ZN(n6133), 
	.B2(\UUT/regfile/reg_out[4][18] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][18] ), 
	.A1(n6376));
   OAI221_X1 U4867 (.ZN(n6135), 
	.C2(n6128), 
	.C1(n5879), 
	.B2(n6027), 
	.B1(n6118), 
	.A(n6117));
   AND2_X1 U4868 (.ZN(n6117), 
	.A2(n6137), 
	.A1(n6136));
   OR3_X1 U4869 (.ZN(n6137), 
	.A3(n5831), 
	.A2(n6045), 
	.A1(n6053));
   NAND2_X1 U4870 (.ZN(n6118), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A1(n6064));
   OAI21_X1 U4871 (.ZN(n6086), 
	.B2(n6138), 
	.B1(n6073), 
	.A(n6139));
   NAND3_X1 U4872 (.ZN(n6139), 
	.A3(n6142), 
	.A2(n6141), 
	.A1(n6140));
   INV_X1 U4873 (.ZN(n6141), 
	.A(n6128));
   INV_X1 U4874 (.ZN(\UUT/Mcontrol/d_instr [6]), 
	.A(n6143));
   OAI21_X1 U4875 (.ZN(n6085), 
	.B2(n6145), 
	.B1(n6144), 
	.A(n6146));
   AOI21_X1 U4876 (.ZN(n6146), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
	.B1(n6078), 
	.A(n6073));
   INV_X1 U4877 (.ZN(n6145), 
	.A(n6142));
   NOR3_X1 U4878 (.ZN(n6142), 
	.A3(n6073), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2019 ), 
	.A1(n6048));
   INV_X1 U4879 (.ZN(n6144), 
	.A(n6039));
   NAND2_X1 U4880 (.ZN(n6039), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A1(n6140));
   AND4_X1 U4881 (.ZN(n6140), 
	.A4(n6042), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1987 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A1(n6043));
   NOR3_X1 U4882 (.ZN(n6043), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N1995 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2007 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2001 ));
   INV_X1 U4883 (.ZN(\UUT/Mcontrol/d_instr [0]), 
	.A(n5428));
   AOI22_X1 U4884 (.ZN(n6147), 
	.B2(\UUT/regfile/reg_out[18][17] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][17] ), 
	.A1(n5534));
   AOI22_X1 U4885 (.ZN(n6148), 
	.B2(\UUT/regfile/reg_out[20][17] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][17] ), 
	.A1(n5539));
   AOI22_X1 U4886 (.ZN(n6149), 
	.B2(\UUT/regfile/reg_out[24][17] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][17] ), 
	.A1(n5544));
   AOI22_X1 U4887 (.ZN(n6150), 
	.B2(\UUT/regfile/reg_out[28][17] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][17] ), 
	.A1(n5549));
   AOI22_X1 U4888 (.ZN(n6151), 
	.B2(\UUT/regfile/reg_out[4][17] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][17] ), 
	.A1(n6376));
   OAI221_X1 U4889 (.ZN(n6153), 
	.C2(n5831), 
	.C1(n6154), 
	.B2(n5888), 
	.B1(n6128), 
	.A(n6136));
   INV_X1 U4890 (.ZN(n6154), 
	.A(n6155));
   AOI22_X1 U4891 (.ZN(n6156), 
	.B2(\UUT/regfile/reg_out[18][16] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][16] ), 
	.A1(n5534));
   AOI22_X1 U4892 (.ZN(n6157), 
	.B2(\UUT/regfile/reg_out[20][16] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][16] ), 
	.A1(n5539));
   AOI22_X1 U4893 (.ZN(n6158), 
	.B2(\UUT/regfile/reg_out[24][16] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][16] ), 
	.A1(n5544));
   AOI22_X1 U4894 (.ZN(n6159), 
	.B2(\UUT/regfile/reg_out[28][16] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][16] ), 
	.A1(n5549));
   AOI22_X1 U4895 (.ZN(n6160), 
	.B2(\UUT/regfile/reg_out[4][16] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][16] ), 
	.A1(n6375));
   OAI221_X1 U4896 (.ZN(n6162), 
	.C2(n6128), 
	.C1(n5896), 
	.B2(n6032), 
	.B1(n6163), 
	.A(n6136));
   AOI22_X1 U4897 (.ZN(n6164), 
	.B2(\UUT/regfile/reg_out[18][15] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][15] ), 
	.A1(n5534));
   AOI22_X1 U4898 (.ZN(n6165), 
	.B2(\UUT/regfile/reg_out[20][15] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][15] ), 
	.A1(n5539));
   AOI22_X1 U4899 (.ZN(n6166), 
	.B2(\UUT/regfile/reg_out[24][15] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][15] ), 
	.A1(n5544));
   AOI22_X1 U4900 (.ZN(n6167), 
	.B2(\UUT/regfile/reg_out[28][15] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][15] ), 
	.A1(n5549));
   AOI22_X1 U4901 (.ZN(n6168), 
	.B2(\UUT/regfile/reg_out[4][15] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][15] ), 
	.A1(n6376));
   AOI21_X1 U4903 (.ZN(n6173), 
	.B2(n6174), 
	.B1(n445), 
	.A(n6127));
   NOR2_X1 U4904 (.ZN(n6127), 
	.A2(n445), 
	.A1(n5831));
   OAI221_X1 U4905 (.ZN(n6174), 
	.C2(n6128), 
	.C1(n6037), 
	.B2(n6033), 
	.B1(n6163), 
	.A(n6136));
   NAND2_X1 U4906 (.ZN(n6136), 
	.A2(\UUT/Mcontrol/d_sampled_finstr [15]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1976 ));
   AOI22_X1 U4907 (.ZN(n6175), 
	.B2(\UUT/regfile/reg_out[18][14] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][14] ), 
	.A1(n5534));
   AOI22_X1 U4908 (.ZN(n6176), 
	.B2(\UUT/regfile/reg_out[20][14] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][14] ), 
	.A1(n5539));
   AOI22_X1 U4909 (.ZN(n6177), 
	.B2(\UUT/regfile/reg_out[24][14] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][14] ), 
	.A1(n5544));
   AOI22_X1 U4910 (.ZN(n6178), 
	.B2(\UUT/regfile/reg_out[28][14] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][14] ), 
	.A1(n5549));
   AOI22_X1 U4911 (.ZN(n6179), 
	.B2(\UUT/regfile/reg_out[4][14] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][14] ), 
	.A1(n6375));
   AOI22_X1 U4913 (.ZN(n6182), 
	.B2(\UUT/regfile/reg_out[18][13] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][13] ), 
	.A1(n5534));
   AOI22_X1 U4914 (.ZN(n6183), 
	.B2(\UUT/regfile/reg_out[20][13] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][13] ), 
	.A1(n5539));
   AOI22_X1 U4915 (.ZN(n6184), 
	.B2(\UUT/regfile/reg_out[24][13] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][13] ), 
	.A1(n5544));
   AOI22_X1 U4916 (.ZN(n6185), 
	.B2(\UUT/regfile/reg_out[28][13] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][13] ), 
	.A1(n5549));
   AOI22_X1 U4917 (.ZN(n6186), 
	.B2(\UUT/regfile/reg_out[4][13] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][13] ), 
	.A1(n6375));
   AOI21_X1 U4919 (.ZN(n6206), 
	.B2(\UUT/Mcontrol/Operation_decoding32/N2036 ), 
	.B1(n6207), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2043 ));
   OAI21_X1 U4920 (.ZN(n6207), 
	.B2(n6074), 
	.B1(n6208), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2030 ));
   AOI211_X1 U4921 (.ZN(n6208), 
	.C2(\UUT/Mcontrol/Operation_decoding32/N1945 ), 
	.C1(n6046), 
	.B(n6064), 
	.A(n6066));
   INV_X1 U4922 (.ZN(n6064), 
	.A(n6210));
   AOI22_X1 U4923 (.ZN(n6211), 
	.B2(\UUT/regfile/reg_out[18][9] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][9] ), 
	.A1(n5534));
   AOI22_X1 U4924 (.ZN(n6212), 
	.B2(\UUT/regfile/reg_out[20][9] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][9] ), 
	.A1(n5539));
   AOI22_X1 U4925 (.ZN(n6213), 
	.B2(\UUT/regfile/reg_out[24][9] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][9] ), 
	.A1(n5544));
   AOI22_X1 U4926 (.ZN(n6214), 
	.B2(\UUT/regfile/reg_out[28][9] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][9] ), 
	.A1(n5549));
   AOI22_X1 U4927 (.ZN(n6215), 
	.B2(\UUT/regfile/reg_out[4][9] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][9] ), 
	.A1(n6376));
   OAI222_X1 U4928 (.ZN(n6216), 
	.C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.C1(n5889), 
	.B2(n6094), 
	.B1(n6163), 
	.A2(n5831), 
	.A1(n6128));
   AOI22_X1 U4929 (.ZN(n6217), 
	.B2(\UUT/regfile/reg_out[18][8] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][8] ), 
	.A1(n5534));
   AOI22_X1 U4930 (.ZN(n6218), 
	.B2(\UUT/regfile/reg_out[20][8] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][8] ), 
	.A1(n5539));
   AOI22_X1 U4931 (.ZN(n6219), 
	.B2(\UUT/regfile/reg_out[24][8] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][8] ), 
	.A1(n5544));
   AOI22_X1 U4932 (.ZN(n6220), 
	.B2(\UUT/regfile/reg_out[28][8] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][8] ), 
	.A1(n5549));
   AOI22_X1 U4933 (.ZN(n6221), 
	.B2(\UUT/regfile/reg_out[4][8] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][8] ), 
	.A1(n6375));
   OAI222_X1 U4934 (.ZN(n6222), 
	.C2(n5897), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n6143), 
	.B1(n6163), 
	.A2(n6032), 
	.A1(n6128));
   AOI22_X1 U4935 (.ZN(n6223), 
	.B2(\UUT/regfile/reg_out[18][7] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][7] ), 
	.A1(n5534));
   AOI22_X1 U4936 (.ZN(n6224), 
	.B2(\UUT/regfile/reg_out[20][7] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][7] ), 
	.A1(n5539));
   AOI22_X1 U4937 (.ZN(n6225), 
	.B2(\UUT/regfile/reg_out[24][7] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][7] ), 
	.A1(n5544));
   AOI22_X1 U4938 (.ZN(n6226), 
	.B2(\UUT/regfile/reg_out[28][7] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][7] ), 
	.A1(n5549));
   AOI22_X1 U4939 (.ZN(n6227), 
	.B2(\UUT/regfile/reg_out[4][7] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][7] ), 
	.A1(n6375));
   OAI222_X1 U4940 (.ZN(n6228), 
	.C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.C1(n6094), 
	.B2(n6163), 
	.B1(n5423), 
	.A2(n6033), 
	.A1(n6128));
   AOI22_X1 U4941 (.ZN(n6229), 
	.B2(\UUT/regfile/reg_out[18][6] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][6] ), 
	.A1(n5534));
   AOI22_X1 U4942 (.ZN(n6230), 
	.B2(\UUT/regfile/reg_out[20][6] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][6] ), 
	.A1(n5539));
   AOI22_X1 U4943 (.ZN(n6231), 
	.B2(\UUT/regfile/reg_out[24][6] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][6] ), 
	.A1(n5544));
   AOI22_X1 U4944 (.ZN(n6232), 
	.B2(\UUT/regfile/reg_out[28][6] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][6] ), 
	.A1(n5549));
   AOI22_X1 U4945 (.ZN(n6233), 
	.B2(\UUT/regfile/reg_out[4][6] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][6] ), 
	.A1(n6375));
   OAI222_X1 U4946 (.ZN(n6234), 
	.C2(n6143), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n6163), 
	.B1(n5424), 
	.A2(n6035), 
	.A1(n6128));
   AOI22_X1 U4947 (.ZN(n6235), 
	.B2(\UUT/regfile/reg_out[18][5] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][5] ), 
	.A1(n5534));
   AOI22_X1 U4948 (.ZN(n6236), 
	.B2(\UUT/regfile/reg_out[20][5] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][5] ), 
	.A1(n5539));
   AOI22_X1 U4949 (.ZN(n6237), 
	.B2(\UUT/regfile/reg_out[24][5] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][5] ), 
	.A1(n5544));
   AOI22_X1 U4950 (.ZN(n6238), 
	.B2(\UUT/regfile/reg_out[28][5] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][5] ), 
	.A1(n5549));
   AOI22_X1 U4951 (.ZN(n6239), 
	.B2(\UUT/regfile/reg_out[4][5] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][5] ), 
	.A1(n6376));
   OAI222_X1 U4952 (.ZN(n6240), 
	.C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.C1(n5423), 
	.B2(n5425), 
	.B1(n6163), 
	.A2(n6036), 
	.A1(n6128));
   AOI22_X1 U4953 (.ZN(n6241), 
	.B2(\UUT/regfile/reg_out[18][4] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][4] ), 
	.A1(n5534));
   AOI22_X1 U4954 (.ZN(n6242), 
	.B2(\UUT/regfile/reg_out[20][4] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][4] ), 
	.A1(n5539));
   AOI22_X1 U4955 (.ZN(n6243), 
	.B2(\UUT/regfile/reg_out[24][4] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][4] ), 
	.A1(n5544));
   AOI22_X1 U4956 (.ZN(n6244), 
	.B2(\UUT/regfile/reg_out[28][4] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][4] ), 
	.A1(n5549));
   AOI22_X1 U4957 (.ZN(n6245), 
	.B2(\UUT/regfile/reg_out[4][4] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][4] ), 
	.A1(n6375));
   OAI22_X1 U4958 (.ZN(n6247), 
	.B2(n6048), 
	.B1(n6248), 
	.A2(n6138), 
	.A1(n5881));
   AOI22_X1 U4959 (.ZN(n6248), 
	.B2(n6209), 
	.B1(\UUT/Mcontrol/d_instr [4]), 
	.A2(n6249), 
	.A1(n445));
   INV_X1 U4960 (.ZN(\UUT/Mcontrol/d_instr [4]), 
	.A(n5424));
   OAI222_X1 U4961 (.ZN(n6249), 
	.C2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.C1(n5424), 
	.B2(n5426), 
	.B1(n6163), 
	.A2(n5881), 
	.A1(n6128));
   AOI22_X1 U4962 (.ZN(n6250), 
	.B2(\UUT/regfile/reg_out[18][3] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][3] ), 
	.A1(n5534));
   AOI22_X1 U4963 (.ZN(n6251), 
	.B2(\UUT/regfile/reg_out[20][3] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][3] ), 
	.A1(n5539));
   AOI22_X1 U4964 (.ZN(n6252), 
	.B2(\UUT/regfile/reg_out[24][3] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][3] ), 
	.A1(n5544));
   AOI22_X1 U4965 (.ZN(n6253), 
	.B2(\UUT/regfile/reg_out[28][3] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][3] ), 
	.A1(n5549));
   AOI22_X1 U4966 (.ZN(n6254), 
	.B2(\UUT/regfile/reg_out[4][3] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][3] ), 
	.A1(n6376));
   OAI22_X1 U4967 (.ZN(n6255), 
	.B2(n6048), 
	.B1(n6256), 
	.A2(n6138), 
	.A1(n5889));
   AOI22_X1 U4968 (.ZN(n6256), 
	.B2(n6209), 
	.B1(\UUT/Mcontrol/d_instr [3]), 
	.A2(n6257), 
	.A1(n445));
   INV_X1 U4969 (.ZN(\UUT/Mcontrol/d_instr [3]), 
	.A(n5425));
   OAI222_X1 U4970 (.ZN(n6257), 
	.C2(n5425), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n5427), 
	.B1(n6163), 
	.A2(n5889), 
	.A1(n6128));
   AOI22_X1 U4971 (.ZN(n6258), 
	.B2(\UUT/regfile/reg_out[18][2] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][2] ), 
	.A1(n5534));
   AOI22_X1 U4972 (.ZN(n6259), 
	.B2(\UUT/regfile/reg_out[20][2] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][2] ), 
	.A1(n5539));
   AOI22_X1 U4973 (.ZN(n6260), 
	.B2(\UUT/regfile/reg_out[24][2] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][2] ), 
	.A1(n5544));
   AOI22_X1 U4974 (.ZN(n6261), 
	.B2(\UUT/regfile/reg_out[28][2] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][2] ), 
	.A1(n5549));
   AOI22_X1 U4975 (.ZN(n6262), 
	.B2(\UUT/regfile/reg_out[4][2] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][2] ), 
	.A1(n6375));
   OAI22_X1 U4976 (.ZN(n6263), 
	.B2(n6048), 
	.B1(n6264), 
	.A2(n6138), 
	.A1(n5897));
   AOI22_X1 U4977 (.ZN(n6264), 
	.B2(n6209), 
	.B1(\UUT/Mcontrol/d_instr [2]), 
	.A2(n6265), 
	.A1(n445));
   INV_X1 U4978 (.ZN(\UUT/Mcontrol/d_instr [2]), 
	.A(n5426));
   OAI222_X1 U4979 (.ZN(n6265), 
	.C2(n5426), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n5428), 
	.B1(n6163), 
	.A2(n5897), 
	.A1(n6128));
   NAND2_X1 U4980 (.ZN(n6138), 
	.A2(n6028), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2037 ));
   AND2_X1 U4981 (.ZN(n6266), 
	.A2(n6030), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N2085 ));
   NOR2_X1 U4982 (.ZN(n6246), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2079 ), 
	.A1(n6073));
   AOI22_X1 U4983 (.ZN(n6267), 
	.B2(\UUT/regfile/reg_out[18][12] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][12] ), 
	.A1(n5534));
   AOI22_X1 U4984 (.ZN(n6268), 
	.B2(\UUT/regfile/reg_out[20][12] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][12] ), 
	.A1(n5539));
   AOI22_X1 U4985 (.ZN(n6269), 
	.B2(\UUT/regfile/reg_out[24][12] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][12] ), 
	.A1(n5544));
   AOI22_X1 U4986 (.ZN(n6270), 
	.B2(\UUT/regfile/reg_out[28][12] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][12] ), 
	.A1(n5549));
   AOI22_X1 U4987 (.ZN(n6271), 
	.B2(\UUT/regfile/reg_out[4][12] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][12] ), 
	.A1(n6375));
   AOI22_X1 U4989 (.ZN(n6273), 
	.B2(\UUT/regfile/reg_out[18][11] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][11] ), 
	.A1(n5534));
   AOI22_X1 U4990 (.ZN(n6274), 
	.B2(\UUT/regfile/reg_out[20][11] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][11] ), 
	.A1(n5539));
   AOI22_X1 U4991 (.ZN(n6275), 
	.B2(\UUT/regfile/reg_out[24][11] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][11] ), 
	.A1(n5544));
   AOI22_X1 U4992 (.ZN(n6276), 
	.B2(\UUT/regfile/reg_out[28][11] ), 
	.B1(n6370), 
	.A2(\UUT/regfile/reg_out[29][11] ), 
	.A1(n5549));
   AOI22_X1 U4993 (.ZN(n6277), 
	.B2(\UUT/regfile/reg_out[4][11] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][11] ), 
	.A1(n6375));
   AOI22_X1 U4995 (.ZN(n6279), 
	.B2(\UUT/regfile/reg_out[18][10] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][10] ), 
	.A1(n5534));
   AOI22_X1 U4996 (.ZN(n6280), 
	.B2(\UUT/regfile/reg_out[20][10] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][10] ), 
	.A1(n5539));
   AOI22_X1 U4997 (.ZN(n6281), 
	.B2(\UUT/regfile/reg_out[24][10] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][10] ), 
	.A1(n5544));
   AOI22_X1 U4998 (.ZN(n6282), 
	.B2(\UUT/regfile/reg_out[28][10] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][10] ), 
	.A1(n5549));
   AOI22_X1 U4999 (.ZN(n6283), 
	.B2(\UUT/regfile/reg_out[4][10] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][10] ), 
	.A1(n6376));
   INV_X1 U5001 (.ZN(n6284), 
	.A(\UUT/Mpath/N115 ));
   NAND3_X1 U5002 (.ZN(\UUT/Mcontrol/d_jump_type[3] ), 
	.A3(n6286), 
	.A2(n6285), 
	.A1(n6056));
   AOI21_X1 U5003 (.ZN(n6286), 
	.B2(n6062), 
	.B1(\UUT/Mcontrol/d_sampled_finstr [19]), 
	.A(n6045));
   NAND2_X1 U5004 (.ZN(n6062), 
	.A2(n6079), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1945 ));
   INV_X1 U5005 (.ZN(n6056), 
	.A(n6054));
   NAND3_X1 U5006 (.ZN(n6054), 
	.A3(n6050), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A1(n445));
   NOR2_X1 U5009 (.ZN(n6291), 
	.A2(\UUT/Mcontrol/st_logic/N70 ), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N25 ));
   AOI21_X1 U5012 (.ZN(n6293), 
	.B2(n6294), 
	.B1(\UUT/Mcontrol/Nextpc_decoding/N247 ), 
	.A(n6296));
   INV_X1 U5018 (.ZN(n6297), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N242 ));
   AOI22_X1 U5020 (.ZN(n6300), 
	.B2(\UUT/regfile/reg_out[18][31] ), 
	.B1(n5535), 
	.A2(\UUT/regfile/reg_out[19][31] ), 
	.A1(n5534));
   AND2_X1 U5025 (.ZN(n6301), 
	.A2(n6306), 
	.A1(n6305));
   AOI22_X1 U5026 (.ZN(n6307), 
	.B2(\UUT/regfile/reg_out[20][31] ), 
	.B1(n5540), 
	.A2(\UUT/regfile/reg_out[21][31] ), 
	.A1(n5539));
   NAND3_X1 U5029 (.ZN(n5537), 
	.A3(n6305), 
	.A2(\UUT/rs1_addr [2]), 
	.A1(n6302));
   NAND4_X1 U5030 (.ZN(n5536), 
	.A4(\UUT/rs1_addr [2]), 
	.A3(\UUT/rs1_addr [0]), 
	.A2(FE_OFN98_UUT_rs1_addr_1_), 
	.A1(n6305));
   NOR2_X1 U5031 (.ZN(n6305), 
	.A2(FE_OFCN199_UUT_rs1_addr_3_), 
	.A1(n6310));
   AOI22_X1 U5032 (.ZN(n6311), 
	.B2(\UUT/regfile/reg_out[24][31] ), 
	.B1(n5545), 
	.A2(\UUT/regfile/reg_out[25][31] ), 
	.A1(n5544));
   AND3_X2 U5033 (.ZN(n5545), 
	.A3(n6312), 
	.A2(n6303), 
	.A1(\UUT/rs1_addr [4]));
   NAND3_X1 U5035 (.ZN(n5542), 
	.A3(n6314), 
	.A2(\UUT/rs1_addr [4]), 
	.A1(n6302));
   AOI22_X1 U5037 (.ZN(n6315), 
	.B2(\UUT/regfile/reg_out[28][31] ), 
	.B1(n6371), 
	.A2(\UUT/regfile/reg_out[29][31] ), 
	.A1(n5549));
   NOR2_X1 U5042 (.ZN(n6313), 
	.A2(n6303), 
	.A1(n6310));
   AOI22_X1 U5045 (.ZN(n6320), 
	.B2(\UUT/regfile/reg_out[4][31] ), 
	.B1(n5557), 
	.A2(\UUT/regfile/reg_out[5][31] ), 
	.A1(n6376));
   NAND3_X1 U5048 (.ZN(n5554), 
	.A3(n6319), 
	.A2(n6318), 
	.A1(\UUT/rs1_addr [2]));
   NAND3_X1 U5049 (.ZN(n5553), 
	.A3(n6317), 
	.A2(\UUT/rs1_addr [2]), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   AND2_X1 U5050 (.ZN(n6317), 
	.A2(n6318), 
	.A1(n6321));
   NOR2_X1 U5053 (.ZN(n6316), 
	.A2(n6306), 
	.A1(n6318));
   NOR2_X1 U5055 (.ZN(n6309), 
	.A2(FE_OFN98_UUT_rs1_addr_1_), 
	.A1(n6306));
   AND2_X1 U5059 (.ZN(n6319), 
	.A2(n6310), 
	.A1(n6302));
   INV_X1 U5061 (.ZN(n6310), 
	.A(\UUT/rs1_addr [4]));
   AND2_X1 U5062 (.ZN(n6312), 
	.A2(n6304), 
	.A1(n6314));
   INV_X1 U5063 (.ZN(n6304), 
	.A(FE_OFN98_UUT_rs1_addr_1_));
   NOR2_X1 U5065 (.ZN(n6314), 
	.A2(\UUT/rs1_addr [2]), 
	.A1(n6318));
   NAND2_X1 U5066 (.ZN(\UUT/rs1_addr [2]), 
	.A2(n5888), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1871 ));
   INV_X1 U5067 (.ZN(n6318), 
	.A(FE_OFCN199_UUT_rs1_addr_3_));
   NOR2_X1 U5068 (.ZN(\UUT/rs1_addr [3]), 
	.A2(n6322), 
	.A1(n5879));
   NOR2_X1 U5069 (.ZN(n6321), 
	.A2(\UUT/rs1_addr [4]), 
	.A1(n6303));
   NOR2_X2 U5070 (.ZN(\UUT/rs1_addr [4]), 
	.A2(n5871), 
	.A1(n6322));
   INV_X1 U5071 (.ZN(n6303), 
	.A(\UUT/rs1_addr [0]));
   NOR2_X2 U5072 (.ZN(\UUT/rs1_addr [0]), 
	.A2(n6322), 
	.A1(n6037));
   INV_X1 U5073 (.ZN(n6322), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1871 ));
   INV_X1 U5077 (.ZN(n6323), 
	.A(n6324));
   NOR3_X1 U5079 (.ZN(n6324), 
	.A3(\UUT/Mpath/the_shift/N111 ), 
	.A2(\UUT/Mpath/the_shift/N118 ), 
	.A1(\UUT/Mpath/the_shift/N115 ));
   INV_X1 U5081 (.ZN(n6325), 
	.A(\UUT/Mpath/the_shift/N115 ));
   NOR3_X1 U5082 (.ZN(n6201), 
	.A3(n6326), 
	.A2(\UUT/Mpath/the_shift/N118 ), 
	.A1(\UUT/Mpath/the_shift/N115 ));
   INV_X1 U5083 (.ZN(n6326), 
	.A(\UUT/Mpath/the_shift/N111 ));
   INV_X1 U5084 (.ZN(n6292), 
	.A(\UUT/Mcontrol/st_logic/N89 ));
   INV_X1 U5085 (.ZN(n6287), 
	.A(\UUT/Mcontrol/Nextpc_decoding/N266 ));
   OAI222_X1 U5086 (.ZN(n6327), 
	.C2(n5881), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n5897), 
	.B1(n6163), 
	.A2(n6027), 
	.A1(n6128));
   OAI21_X1 U5088 (.ZN(n6155), 
	.B2(n6066), 
	.B1(n6045), 
	.A(n6210));
   NAND2_X1 U5089 (.ZN(n6066), 
	.A2(n6040), 
	.A1(n6328));
   INV_X1 U5093 (.ZN(n6067), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1928 ));
   NOR2_X1 U5096 (.ZN(n6046), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1940 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1934 ));
   INV_X1 U5097 (.ZN(n6285), 
	.A(n6053));
   INV_X1 U5100 (.ZN(n6040), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1958 ));
   INV_X1 U5101 (.ZN(n6328), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1952 ));
   NAND2_X1 U5103 (.ZN(n6209), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1981 ), 
	.A1(n6116));
   NOR2_X1 U5104 (.ZN(n6172), 
	.A2(n6170), 
	.A1(n6048));
   NOR2_X1 U5105 (.ZN(n6078), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2025 ), 
	.A1(n6587));
   INV_X1 U5106 (.ZN(BUS_MW), 
	.A(\localbus/N90 ));
   INV_X1 U5107 (.ZN(BUS_MR), 
	.A(\localbus/N86 ));
   NOR2_X1 U5108 (.ZN(BUS_DATA_OUTBUS[9]), 
	.A2(n6329), 
	.A1(n4376));
   AOI22_X1 U5109 (.ZN(n4376), 
	.B2(D_DATA_OUTBUS[1]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[9] ), 
	.A1(n6330));
   NOR2_X1 U5110 (.ZN(BUS_DATA_OUTBUS[8]), 
	.A2(n6329), 
	.A1(n4378));
   AOI22_X1 U5111 (.ZN(n4378), 
	.B2(D_DATA_OUTBUS[0]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[8] ), 
	.A1(n6330));
   NOR2_X1 U5112 (.ZN(BUS_DATA_OUTBUS[7]), 
	.A2(n6332), 
	.A1(n4380));
   NOR2_X1 U5113 (.ZN(BUS_DATA_OUTBUS[6]), 
	.A2(n6332), 
	.A1(n4381));
   NOR2_X1 U5114 (.ZN(BUS_DATA_OUTBUS[5]), 
	.A2(n6332), 
	.A1(n4382));
   NOR2_X1 U5115 (.ZN(BUS_DATA_OUTBUS[4]), 
	.A2(n6332), 
	.A1(n4383));
   NOR2_X1 U5116 (.ZN(BUS_DATA_OUTBUS[3]), 
	.A2(n6332), 
	.A1(n4384));
   NOR2_X1 U5117 (.ZN(BUS_DATA_OUTBUS[31]), 
	.A2(n6329), 
	.A1(n4385));
   AOI221_X1 U5118 (.ZN(n4385), 
	.C2(D_DATA_OUTBUS[7]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
	.B1(n6333), 
	.A(n6334));
   AND2_X1 U5119 (.ZN(n6334), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[31] ));
   NOR2_X1 U5120 (.ZN(BUS_DATA_OUTBUS[30]), 
	.A2(n6329), 
	.A1(n4386));
   AOI221_X1 U5121 (.ZN(n4386), 
	.C2(D_DATA_OUTBUS[6]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
	.B1(n6333), 
	.A(n6336));
   AND2_X1 U5122 (.ZN(n6336), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[30] ));
   NOR2_X1 U5123 (.ZN(BUS_DATA_OUTBUS[2]), 
	.A2(n6332), 
	.A1(n4387));
   NOR2_X1 U5124 (.ZN(BUS_DATA_OUTBUS[29]), 
	.A2(n6329), 
	.A1(n4388));
   AOI221_X1 U5125 (.ZN(n4388), 
	.C2(D_DATA_OUTBUS[5]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
	.B1(n6333), 
	.A(n6337));
   AND2_X1 U5126 (.ZN(n6337), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[29] ));
   NOR2_X1 U5127 (.ZN(BUS_DATA_OUTBUS[28]), 
	.A2(n6329), 
	.A1(n4389));
   AOI221_X1 U5128 (.ZN(n4389), 
	.C2(D_DATA_OUTBUS[4]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
	.B1(n6333), 
	.A(n6338));
   AND2_X1 U5129 (.ZN(n6338), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[28] ));
   NOR2_X1 U5130 (.ZN(BUS_DATA_OUTBUS[27]), 
	.A2(n6329), 
	.A1(n4390));
   AOI221_X1 U5131 (.ZN(n4390), 
	.C2(D_DATA_OUTBUS[3]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
	.B1(n6333), 
	.A(n6339));
   AND2_X1 U5132 (.ZN(n6339), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[27] ));
   NOR2_X1 U5133 (.ZN(BUS_DATA_OUTBUS[26]), 
	.A2(n6329), 
	.A1(n4391));
   AOI221_X1 U5134 (.ZN(n4391), 
	.C2(D_DATA_OUTBUS[2]), 
	.C1(n6331), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
	.B1(n6333), 
	.A(n6340));
   AND2_X1 U5135 (.ZN(n6340), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[26] ));
   NOR2_X1 U5136 (.ZN(BUS_DATA_OUTBUS[25]), 
	.A2(n6329), 
	.A1(n4392));
   AOI221_X1 U5137 (.ZN(n4392), 
	.C2(D_DATA_OUTBUS[1]), 
	.C1(n6331), 
	.B2(n6333), 
	.B1(\UUT/Mpath/the_memhandle/smdr_out[9] ), 
	.A(n6341));
   AND2_X1 U5138 (.ZN(n6341), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[25] ));
   NOR2_X1 U5139 (.ZN(BUS_DATA_OUTBUS[24]), 
	.A2(n6329), 
	.A1(n4393));
   AOI221_X1 U5140 (.ZN(n4393), 
	.C2(D_DATA_OUTBUS[0]), 
	.C1(n6331), 
	.B2(n6333), 
	.B1(\UUT/Mpath/the_memhandle/smdr_out[8] ), 
	.A(n6342));
   AND2_X1 U5141 (.ZN(n6342), 
	.A2(n6335), 
	.A1(\UUT/Mpath/the_memhandle/smdr_out[24] ));
   INV_X1 U5142 (.ZN(n6333), 
	.A(n6343));
   NOR2_X1 U5143 (.ZN(BUS_DATA_OUTBUS[23]), 
	.A2(n6329), 
	.A1(n4394));
   AOI22_X1 U5144 (.ZN(n4394), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[23] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[7]), 
	.A1(n6344));
   NOR2_X1 U5145 (.ZN(BUS_DATA_OUTBUS[22]), 
	.A2(n6329), 
	.A1(n4395));
   AOI22_X1 U5146 (.ZN(n4395), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[22] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[6]), 
	.A1(n6344));
   NOR2_X1 U5147 (.ZN(BUS_DATA_OUTBUS[21]), 
	.A2(n6329), 
	.A1(n4396));
   AOI22_X1 U5148 (.ZN(n4396), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[21] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[5]), 
	.A1(n6344));
   NOR2_X1 U5149 (.ZN(BUS_DATA_OUTBUS[20]), 
	.A2(n6329), 
	.A1(n4397));
   AOI22_X1 U5150 (.ZN(n4397), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[20] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[4]), 
	.A1(n6344));
   NOR2_X1 U5151 (.ZN(BUS_DATA_OUTBUS[1]), 
	.A2(n6332), 
	.A1(n4398));
   NOR2_X1 U5152 (.ZN(BUS_DATA_OUTBUS[19]), 
	.A2(n6329), 
	.A1(n4399));
   AOI22_X1 U5153 (.ZN(n4399), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[19] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[3]), 
	.A1(n6344));
   NOR2_X1 U5154 (.ZN(BUS_DATA_OUTBUS[18]), 
	.A2(n6329), 
	.A1(n4400));
   AOI22_X1 U5155 (.ZN(n4400), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[18] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[2]), 
	.A1(n6344));
   NOR2_X1 U5156 (.ZN(BUS_DATA_OUTBUS[17]), 
	.A2(n6329), 
	.A1(n4401));
   AOI22_X1 U5157 (.ZN(n4401), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[17] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[1]), 
	.A1(n6344));
   NOR2_X1 U5158 (.ZN(BUS_DATA_OUTBUS[16]), 
	.A2(n6329), 
	.A1(n4402));
   AOI22_X1 U5159 (.ZN(n4402), 
	.B2(\UUT/Mpath/the_memhandle/smdr_out[16] ), 
	.B1(n6335), 
	.A2(D_DATA_OUTBUS[0]), 
	.A1(n6344));
   AND2_X1 U5160 (.ZN(n6335), 
	.A2(dmem_ishalf), 
	.A1(n6330));
   NAND2_X1 U5161 (.ZN(n6344), 
	.A2(n6343), 
	.A1(n6345));
   NAND2_X1 U5162 (.ZN(n6343), 
	.A2(n6330), 
	.A1(\UUT/Mpath/the_memhandle/N237 ));
   NOR2_X1 U5163 (.ZN(BUS_DATA_OUTBUS[15]), 
	.A2(n6329), 
	.A1(n4403));
   AOI22_X1 U5164 (.ZN(n4403), 
	.B2(D_DATA_OUTBUS[7]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[15] ), 
	.A1(n6330));
   NOR2_X1 U5165 (.ZN(BUS_DATA_OUTBUS[14]), 
	.A2(n6329), 
	.A1(n4404));
   AOI22_X1 U5166 (.ZN(n4404), 
	.B2(D_DATA_OUTBUS[6]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[14] ), 
	.A1(n6330));
   NOR2_X1 U5167 (.ZN(BUS_DATA_OUTBUS[13]), 
	.A2(n6329), 
	.A1(n4405));
   AOI22_X1 U5168 (.ZN(n4405), 
	.B2(D_DATA_OUTBUS[5]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[13] ), 
	.A1(n6330));
   NOR2_X1 U5169 (.ZN(BUS_DATA_OUTBUS[12]), 
	.A2(n6329), 
	.A1(n4406));
   AOI22_X1 U5170 (.ZN(n4406), 
	.B2(D_DATA_OUTBUS[4]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[12] ), 
	.A1(n6330));
   NOR2_X1 U5171 (.ZN(BUS_DATA_OUTBUS[11]), 
	.A2(n6329), 
	.A1(n4407));
   AOI22_X1 U5172 (.ZN(n4407), 
	.B2(D_DATA_OUTBUS[3]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[11] ), 
	.A1(n6330));
   NOR2_X1 U5173 (.ZN(BUS_DATA_OUTBUS[10]), 
	.A2(n6329), 
	.A1(n4408));
   INV_X1 U5174 (.ZN(n6329), 
	.A(\localbus/N229 ));
   AOI22_X1 U5175 (.ZN(n4408), 
	.B2(D_DATA_OUTBUS[2]), 
	.B1(n6331), 
	.A2(\UUT/Mpath/the_memhandle/smdr_out[10] ), 
	.A1(n6330));
   INV_X1 U5176 (.ZN(n6331), 
	.A(n6345));
   NAND2_X1 U5177 (.ZN(n6345), 
	.A2(\UUT/Mpath/the_memhandle/N234 ), 
	.A1(\localbus/N51 ));
   AND2_X1 U5178 (.ZN(n6330), 
	.A2(dmem_isbyte), 
	.A1(\localbus/N51 ));
   NOR2_X1 U5179 (.ZN(BUS_DATA_OUTBUS[0]), 
	.A2(n6332), 
	.A1(n4409));
   NAND2_X1 U5180 (.ZN(n6332), 
	.A2(\localbus/N51 ), 
	.A1(\localbus/N229 ));
   NOR2_X1 U5181 (.ZN(BUS_ADDR_OUTBUS[9]), 
	.A2(\localbus/N225 ), 
	.A1(n4344));
   NAND2_X1 U5182 (.ZN(n4344), 
	.A2(n6189), 
	.A1(n6347));
   NOR2_X1 U5183 (.ZN(BUS_ADDR_OUTBUS[8]), 
	.A2(\localbus/N225 ), 
	.A1(n4345));
   NAND2_X1 U5184 (.ZN(n4345), 
	.A2(n6190), 
	.A1(n6347));
   NOR2_X1 U5185 (.ZN(BUS_ADDR_OUTBUS[7]), 
	.A2(\localbus/N225 ), 
	.A1(n4346));
   NAND2_X1 U5186 (.ZN(n4346), 
	.A2(n6191), 
	.A1(n6347));
   NOR2_X1 U5187 (.ZN(BUS_ADDR_OUTBUS[6]), 
	.A2(\localbus/N225 ), 
	.A1(n4347));
   NAND2_X1 U5188 (.ZN(n4347), 
	.A2(n6192), 
	.A1(n6347));
   NOR2_X1 U5189 (.ZN(BUS_ADDR_OUTBUS[5]), 
	.A2(\localbus/N225 ), 
	.A1(n4348));
   NAND2_X1 U5190 (.ZN(n4348), 
	.A2(n6193), 
	.A1(n6347));
   NOR2_X1 U5191 (.ZN(BUS_ADDR_OUTBUS[4]), 
	.A2(\localbus/N225 ), 
	.A1(n4349));
   NAND2_X1 U5192 (.ZN(n4349), 
	.A2(n6194), 
	.A1(n6347));
   NOR2_X1 U5193 (.ZN(BUS_ADDR_OUTBUS[3]), 
	.A2(\localbus/N225 ), 
	.A1(n4350));
   NAND2_X1 U5194 (.ZN(n4350), 
	.A2(n6195), 
	.A1(n6347));
   NOR2_X1 U5195 (.ZN(BUS_ADDR_OUTBUS[31]), 
	.A2(n6425), 
	.A1(\localbus/N225 ));
   NOR2_X1 U5197 (.ZN(BUS_ADDR_OUTBUS[30]), 
	.A2(n4352), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5198 (.ZN(n4352), 
	.A2(n5563), 
	.A1(n6347));
   NOR2_X1 U5199 (.ZN(BUS_ADDR_OUTBUS[2]), 
	.A2(\localbus/N225 ), 
	.A1(n4353));
   NAND2_X1 U5200 (.ZN(n4353), 
	.A2(n6202), 
	.A1(n6347));
   NOR2_X1 U5201 (.ZN(BUS_ADDR_OUTBUS[29]), 
	.A2(n4354), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5202 (.ZN(n4354), 
	.A2(n5571), 
	.A1(n6347));
   NOR2_X1 U5203 (.ZN(BUS_ADDR_OUTBUS[28]), 
	.A2(n4355), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5204 (.ZN(n4355), 
	.A2(n5578), 
	.A1(n6347));
   NOR2_X1 U5205 (.ZN(BUS_ADDR_OUTBUS[27]), 
	.A2(n4356), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5206 (.ZN(n4356), 
	.A2(n5585), 
	.A1(n6347));
   NOR2_X1 U5207 (.ZN(BUS_ADDR_OUTBUS[26]), 
	.A2(n4357), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5208 (.ZN(n4357), 
	.A2(n5592), 
	.A1(n6347));
   NOR2_X1 U5209 (.ZN(BUS_ADDR_OUTBUS[25]), 
	.A2(n4358), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5210 (.ZN(n4358), 
	.A2(n5599), 
	.A1(n6347));
   NOR2_X1 U5211 (.ZN(BUS_ADDR_OUTBUS[24]), 
	.A2(n4359), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5212 (.ZN(n4359), 
	.A2(n5606), 
	.A1(n6347));
   NOR2_X1 U5213 (.ZN(BUS_ADDR_OUTBUS[23]), 
	.A2(n4360), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5214 (.ZN(n4360), 
	.A2(n6092), 
	.A1(n6347));
   NOR2_X1 U5215 (.ZN(BUS_ADDR_OUTBUS[22]), 
	.A2(n4361), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5216 (.ZN(n4361), 
	.A2(n6100), 
	.A1(n6347));
   NOR2_X1 U5217 (.ZN(BUS_ADDR_OUTBUS[21]), 
	.A2(n4362), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5218 (.ZN(n4362), 
	.A2(n6107), 
	.A1(n6347));
   NOR2_X1 U5219 (.ZN(BUS_ADDR_OUTBUS[20]), 
	.A2(n4363), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5220 (.ZN(n4363), 
	.A2(n6114), 
	.A1(n6347));
   NOR2_X1 U5221 (.ZN(BUS_ADDR_OUTBUS[1]), 
	.A2(n4364), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5222 (.ZN(n4364), 
	.A2(\localbus/N50 ), 
	.A1(D_ADDR_OUTBUS[1]));
   AND2_X1 U5223 (.ZN(D_ADDR_OUTBUS[1]), 
	.A2(\UUT/daddr_out [1]), 
	.A1(\UUT/N3 ));
   NOR2_X1 U5224 (.ZN(BUS_ADDR_OUTBUS[19]), 
	.A2(n4365), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5225 (.ZN(n4365), 
	.A2(n6124), 
	.A1(n6347));
   NOR2_X1 U5226 (.ZN(BUS_ADDR_OUTBUS[18]), 
	.A2(n4366), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5227 (.ZN(n4366), 
	.A2(n6134), 
	.A1(n6347));
   NOR2_X1 U5228 (.ZN(BUS_ADDR_OUTBUS[17]), 
	.A2(n4367), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5229 (.ZN(n4367), 
	.A2(n6152), 
	.A1(n6347));
   NOR2_X1 U5230 (.ZN(BUS_ADDR_OUTBUS[16]), 
	.A2(n4368), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5231 (.ZN(n4368), 
	.A2(n6161), 
	.A1(n6347));
   NOR2_X1 U5232 (.ZN(BUS_ADDR_OUTBUS[15]), 
	.A2(n4369), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5233 (.ZN(n4369), 
	.A2(n6169), 
	.A1(n6347));
   NOR2_X1 U5234 (.ZN(BUS_ADDR_OUTBUS[14]), 
	.A2(n4370), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5235 (.ZN(n4370), 
	.A2(n6180), 
	.A1(n6347));
   NOR2_X1 U5236 (.ZN(BUS_ADDR_OUTBUS[13]), 
	.A2(n4371), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5237 (.ZN(n4371), 
	.A2(n6187), 
	.A1(n6347));
   NOR2_X1 U5238 (.ZN(BUS_ADDR_OUTBUS[12]), 
	.A2(\localbus/N225 ), 
	.A1(n4372));
   NAND2_X1 U5239 (.ZN(n4372), 
	.A2(n6203), 
	.A1(n6347));
   NOR2_X1 U5240 (.ZN(BUS_ADDR_OUTBUS[11]), 
	.A2(\localbus/N225 ), 
	.A1(n4373));
   NAND2_X1 U5241 (.ZN(n4373), 
	.A2(n6204), 
	.A1(n6347));
   NOR2_X1 U5242 (.ZN(BUS_ADDR_OUTBUS[10]), 
	.A2(\localbus/N225 ), 
	.A1(n4374));
   NAND2_X1 U5243 (.ZN(n4374), 
	.A2(n6205), 
	.A1(n6347));
   NAND2_X1 U5244 (.ZN(n6349), 
	.A2(n6350), 
	.A1(n6348));
   INV_X1 U5245 (.ZN(n6350), 
	.A(\UUT/Mpath/the_alu/N492 ));
   NOR2_X1 U5247 (.ZN(BUS_ADDR_OUTBUS[0]), 
	.A2(n4375), 
	.A1(\localbus/N225 ));
   NAND2_X1 U5248 (.ZN(n4375), 
	.A2(\localbus/N50 ), 
	.A1(D_ADDR_OUTBUS[0]));
   AND2_X1 U5249 (.ZN(D_ADDR_OUTBUS[0]), 
	.A2(\UUT/daddr_out [0]), 
	.A1(\UUT/N3 ));
   OAI21_X1 U5250 (.ZN(n6351), 
	.B2(n6352), 
	.B1(\UUT/Mpath/the_alu/N492 ), 
	.A(n6353));
   NAND2_X1 U5251 (.ZN(n6353), 
	.A2(\UUT/Mpath/the_alu/N492 ), 
	.A1(\UUT/Mpath/the_alu/N125 ));
   AOI22_X1 U5252 (.ZN(n6352), 
	.B2(\UUT/Mpath/the_alu/N486 ), 
	.B1(\UUT/Mpath/the_alu/N157 ), 
	.A2(\UUT/Mpath/the_alu/N485 ), 
	.A1(n6354));
   OAI21_X1 U5253 (.ZN(n6354), 
	.B2(n6355), 
	.B1(\UUT/Mpath/the_alu/N480 ), 
	.A(n6356));
   NAND2_X1 U5254 (.ZN(n6356), 
	.A2(\UUT/Mpath/the_alu/N480 ), 
	.A1(\UUT/Mpath/the_alu/N189 ));
   AOI22_X1 U5255 (.ZN(n6355), 
	.B2(FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_), 
	.B1(\UUT/Mpath/the_alu/N473 ), 
	.A2(\UUT/Mpath/the_alu/N474 ), 
	.A1(\UUT/Mpath/the_alu/N221 ));
   up_island_DW01_add_0 \UUT/Mpath/the_mult/accumulate/add_391  (.A({ 1'b0,
		\UUT/Mpath/the_mult/acc_out[63] ,
		\UUT/Mpath/the_mult/acc_out[62] ,
		\UUT/Mpath/the_mult/acc_out[61] ,
		\UUT/Mpath/the_mult/acc_out[60] ,
		\UUT/Mpath/the_mult/acc_out[59] ,
		\UUT/Mpath/the_mult/acc_out[58] ,
		\UUT/Mpath/the_mult/acc_out[57] ,
		\UUT/Mpath/the_mult/acc_out[56] ,
		\UUT/Mpath/the_mult/acc_out[55] ,
		\UUT/Mpath/the_mult/acc_out[54] ,
		\UUT/Mpath/the_mult/acc_out[53] ,
		\UUT/Mpath/the_mult/acc_out[52] ,
		\UUT/Mpath/the_mult/acc_out[51] ,
		\UUT/Mpath/the_mult/acc_out[50] ,
		\UUT/Mpath/the_mult/acc_out[49] ,
		\UUT/Mpath/the_mult/acc_out[48] ,
		\UUT/Mpath/the_mult/acc_out[47] ,
		\UUT/Mpath/the_mult/acc_out[46] ,
		\UUT/Mpath/the_mult/acc_out[45] ,
		\UUT/Mpath/the_mult/acc_out[44] ,
		\UUT/Mpath/the_mult/acc_out[43] ,
		\UUT/Mpath/the_mult/acc_out[42] ,
		\UUT/Mpath/the_mult/acc_out[41] ,
		\UUT/Mpath/the_mult/acc_out[40] ,
		\UUT/Mpath/the_mult/acc_out[39] ,
		\UUT/Mpath/the_mult/acc_out[38] ,
		\UUT/Mpath/the_mult/acc_out[37] ,
		\UUT/Mpath/the_mult/acc_out[36] ,
		\UUT/Mpath/the_mult/acc_out[35] ,
		\UUT/Mpath/the_mult/acc_out[34] ,
		\UUT/Mpath/the_mult/acc_out[33] ,
		\UUT/Mpath/the_mult/acc_out[32] ,
		\UUT/Mpath/the_mult/acc_out[31] ,
		\UUT/Mpath/the_mult/acc_out[30] ,
		\UUT/Mpath/the_mult/acc_out[29] ,
		\UUT/Mpath/the_mult/acc_out[28] ,
		\UUT/Mpath/the_mult/acc_out[27] ,
		\UUT/Mpath/the_mult/acc_out[26] ,
		\UUT/Mpath/the_mult/acc_out[25] ,
		\UUT/Mpath/the_mult/acc_out[24] ,
		\UUT/Mpath/the_mult/acc_out[23] ,
		\UUT/Mpath/the_mult/acc_out[22] ,
		\UUT/Mpath/the_mult/acc_out[21] ,
		\UUT/Mpath/the_mult/acc_out[20] ,
		\UUT/Mpath/the_mult/acc_out[19] ,
		\UUT/Mpath/the_mult/acc_out[18] ,
		\UUT/Mpath/the_mult/acc_out[17] ,
		\UUT/Mpath/the_mult/acc_out[16] ,
		\UUT/Mpath/the_mult/acc_out[15] ,
		\UUT/Mpath/the_mult/acc_out[14] ,
		\UUT/Mpath/the_mult/acc_out[13] ,
		\UUT/Mpath/the_mult/acc_out[12] ,
		\UUT/Mpath/the_mult/acc_out[11] ,
		\UUT/Mpath/the_mult/acc_out[10] ,
		\UUT/Mpath/the_mult/acc_out[9] ,
		\UUT/Mpath/the_mult/acc_out[8] ,
		\UUT/Mpath/the_mult/acc_out[7] ,
		\UUT/Mpath/the_mult/acc_out[6] ,
		\UUT/Mpath/the_mult/acc_out[5] ,
		\UUT/Mpath/the_mult/acc_out[4] ,
		\UUT/Mpath/the_mult/acc_out[3] ,
		\UUT/Mpath/the_mult/acc_out[2] ,
		\UUT/Mpath/the_mult/acc_out[1] ,
		\UUT/Mpath/the_mult/acc_out[0]  }), 
	.B({ 1'b0,
		\UUT/Mpath/the_mult/Mult_out[63] ,
		\UUT/Mpath/the_mult/Mult_out[62] ,
		\UUT/Mpath/the_mult/Mult_out[61] ,
		\UUT/Mpath/the_mult/Mult_out[60] ,
		\UUT/Mpath/the_mult/Mult_out[59] ,
		\UUT/Mpath/the_mult/Mult_out[58] ,
		\UUT/Mpath/the_mult/Mult_out[57] ,
		\UUT/Mpath/the_mult/Mult_out[56] ,
		\UUT/Mpath/the_mult/Mult_out[55] ,
		\UUT/Mpath/the_mult/Mult_out[54] ,
		\UUT/Mpath/the_mult/Mult_out[53] ,
		\UUT/Mpath/the_mult/Mult_out[52] ,
		\UUT/Mpath/the_mult/Mult_out[51] ,
		\UUT/Mpath/the_mult/Mult_out[50] ,
		\UUT/Mpath/the_mult/Mult_out[49] ,
		\UUT/Mpath/the_mult/Mult_out[48] ,
		\UUT/Mpath/the_mult/Mult_out[47] ,
		\UUT/Mpath/the_mult/Mult_out[46] ,
		\UUT/Mpath/the_mult/Mult_out[45] ,
		\UUT/Mpath/the_mult/Mult_out[44] ,
		\UUT/Mpath/the_mult/Mult_out[43] ,
		\UUT/Mpath/the_mult/Mult_out[42] ,
		\UUT/Mpath/the_mult/Mult_out[41] ,
		\UUT/Mpath/the_mult/Mult_out[40] ,
		\UUT/Mpath/the_mult/Mult_out[39] ,
		\UUT/Mpath/the_mult/Mult_out[38] ,
		\UUT/Mpath/the_mult/Mult_out[37] ,
		\UUT/Mpath/the_mult/Mult_out[36] ,
		\UUT/Mpath/the_mult/Mult_out[35] ,
		\UUT/Mpath/the_mult/Mult_out[34] ,
		\UUT/Mpath/the_mult/Mult_out[33] ,
		\UUT/Mpath/the_mult/Mult_out[32] ,
		\UUT/Mpath/the_mult/Mult_out[31] ,
		\UUT/Mpath/the_mult/Mult_out[30] ,
		\UUT/Mpath/the_mult/Mult_out[29] ,
		\UUT/Mpath/the_mult/Mult_out[28] ,
		\UUT/Mpath/the_mult/Mult_out[27] ,
		\UUT/Mpath/the_mult/Mult_out[26] ,
		\UUT/Mpath/the_mult/Mult_out[25] ,
		\UUT/Mpath/the_mult/Mult_out[24] ,
		\UUT/Mpath/the_mult/Mult_out[23] ,
		\UUT/Mpath/the_mult/Mult_out[22] ,
		\UUT/Mpath/the_mult/Mult_out[21] ,
		\UUT/Mpath/the_mult/Mult_out[20] ,
		\UUT/Mpath/the_mult/Mult_out[19] ,
		\UUT/Mpath/the_mult/Mult_out[18] ,
		\UUT/Mpath/the_mult/Mult_out[17] ,
		\UUT/Mpath/the_mult/Mult_out[16] ,
		\UUT/Mpath/the_mult/Mult_out[15] ,
		\UUT/Mpath/the_mult/Mult_out[14] ,
		\UUT/Mpath/the_mult/Mult_out[13] ,
		\UUT/Mpath/the_mult/Mult_out[12] ,
		\UUT/Mpath/the_mult/Mult_out[11] ,
		\UUT/Mpath/the_mult/Mult_out[10] ,
		\UUT/Mpath/the_mult/Mult_out[9] ,
		\UUT/Mpath/the_mult/Mult_out[8] ,
		\UUT/Mpath/the_mult/Mult_out[7] ,
		\UUT/Mpath/the_mult/Mult_out[6] ,
		\UUT/Mpath/the_mult/Mult_out[5] ,
		\UUT/Mpath/the_mult/Mult_out[4] ,
		\UUT/Mpath/the_mult/Mult_out[3] ,
		\UUT/Mpath/the_mult/Mult_out[2] ,
		\UUT/Mpath/the_mult/Mult_out[1] ,
		\UUT/Mpath/the_mult/Mult_out[0]  }), 
	.CI(1'b0), 
	.SUM({ SYNOPSYS_UNCONNECTED__0,
		\UUT/Mpath/the_mult/Mad_out  }), 
	.FE_PT1_n380(n380), 
	.n806(n806), 
	.n769(n769), 
	.n555(n555), 
	.n529(n529), 
	.n746(n746), 
	.n402(n402), 
	.n632(n632), 
	.n454(n454), 
	.n580(n580), 
	.n599(n599), 
	.n577(n577), 
	.FE_PT1_n213(n213), 
	.n615(n615), 
	.n552(n552), 
	.n424(n424), 
	.n794(n794), 
	.n772(n772), 
	.n723(n723), 
	.n700(n700), 
	.n946(n946), 
	.n635(n635), 
	.n861(n861));
   up_island_DW01_add_1 \UUT/Mcontrol/Nextpc_decoding/bta_calc/add_391  (.A({ 1'b0,
		\UUT/Mcontrol/f_currpc  }), 
	.B({ 1'b0,
		\UUT/break_code[23] ,
		\UUT/break_code[22] ,
		\UUT/break_code[21] ,
		\UUT/break_code[20] ,
		\UUT/break_code[19] ,
		\UUT/break_code[18] ,
		\UUT/break_code[17] ,
		\UUT/break_code[16] ,
		\UUT/break_code[15] ,
		\UUT/break_code[14] ,
		\UUT/break_code[13] ,
		\UUT/break_code[12] ,
		\UUT/break_code[11] ,
		\UUT/break_code[10] ,
		\UUT/break_code[9] ,
		\UUT/break_code[8] ,
		\UUT/break_code[7] ,
		\UUT/break_code[6] ,
		\UUT/break_code[5] ,
		\UUT/break_code[4] ,
		\UUT/break_code[3] ,
		\UUT/break_code[2] ,
		\UUT/break_code[1] ,
		\UUT/break_code[0]  }), 
	.CI(1'b0), 
	.SUM({ SYNOPSYS_UNCONNECTED__1,
		\UUT/Mcontrol/Nextpc_decoding/Bta  }));
   up_island_DW01_add_2 \UUT/Mcontrol/Nextpc_decoding/incr/add_391  (.A({ 1'b0,
		\UUT/Mcontrol/f_currpc  }), 
	.B({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b1,
		1'b0,
		1'b0 }), 
	.CI(1'b0), 
	.SUM({ SYNOPSYS_UNCONNECTED__2,
		\UUT/jar_in  }));
   up_island_DW01_cmp6_0 r771 (.A({ n6488,
		\UUT/branch_rega [30],
		\UUT/branch_rega [29],
		\UUT/branch_rega [28],
		\UUT/branch_rega [27],
		\UUT/branch_rega [26],
		\UUT/branch_rega [25],
		\UUT/branch_rega [24],
		\UUT/branch_rega [23],
		\UUT/branch_rega [22],
		\UUT/branch_rega [21],
		\UUT/branch_rega [20],
		\UUT/branch_rega [19],
		\UUT/branch_rega [18],
		\UUT/branch_rega [17],
		\UUT/branch_rega [16],
		\UUT/branch_rega [15],
		\UUT/branch_rega [14],
		\UUT/branch_rega [13],
		\UUT/branch_rega [12],
		\UUT/branch_rega [11],
		\UUT/branch_rega [10],
		\UUT/branch_rega [9],
		\UUT/branch_rega [8],
		\UUT/branch_rega [7],
		\UUT/branch_rega [6],
		\UUT/branch_rega [5],
		\UUT/branch_rega [4],
		\UUT/branch_rega [3],
		\UUT/branch_rega [2],
		FE_OFN187_UUT_branch_rega_1_,
		\UUT/branch_rega [0] }), 
	.B(\UUT/branch_regb ), 
	.TC(1'b0), 
	.EQ(\UUT/Mcontrol/Nextpc_decoding/N22 ), 
	.NE(\UUT/Mcontrol/Nextpc_decoding/N25 ), 
	.n6832(n6832));
   up_island_DW01_sub_0 \UUT/Mpath/the_alu/sub_96  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.B({ \UUT/Mpath/out_regB[31] ,
		\UUT/Mpath/out_regB[30] ,
		\UUT/Mpath/out_regB[29] ,
		\UUT/Mpath/out_regB[28] ,
		\UUT/Mpath/out_regB[27] ,
		\UUT/Mpath/out_regB[26] ,
		\UUT/Mpath/out_regB[25] ,
		\UUT/Mpath/out_regB[24] ,
		\UUT/Mpath/out_regB[23] ,
		\UUT/Mpath/out_regB[22] ,
		\UUT/Mpath/out_regB[21] ,
		\UUT/Mpath/out_regB[20] ,
		\UUT/Mpath/out_regB[19] ,
		\UUT/Mpath/out_regB[18] ,
		\UUT/Mpath/out_regB[17] ,
		\UUT/Mpath/out_regB[16] ,
		\UUT/Mpath/out_regB[15] ,
		\UUT/Mpath/out_regB[14] ,
		\UUT/Mpath/out_regB[13] ,
		\UUT/Mpath/out_regB[12] ,
		\UUT/Mpath/out_regB[11] ,
		\UUT/Mpath/out_regB[10] ,
		\UUT/Mpath/out_regB[9] ,
		\UUT/Mpath/out_regB[8] ,
		\UUT/Mpath/out_regB[7] ,
		\UUT/Mpath/out_regB[6] ,
		\UUT/Mpath/out_regB[5] ,
		FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		\UUT/Mpath/out_regB[1] ,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.CI(1'b0), 
	.DIFF({ \UUT/Mpath/the_alu/diff[31] ,
		\UUT/Mpath/the_alu/diff[30] ,
		\UUT/Mpath/the_alu/diff[29] ,
		\UUT/Mpath/the_alu/diff[28] ,
		\UUT/Mpath/the_alu/diff[27] ,
		\UUT/Mpath/the_alu/diff[26] ,
		\UUT/Mpath/the_alu/diff[25] ,
		\UUT/Mpath/the_alu/diff[24] ,
		\UUT/Mpath/the_alu/diff[23] ,
		\UUT/Mpath/the_alu/diff[22] ,
		\UUT/Mpath/the_alu/diff[21] ,
		\UUT/Mpath/the_alu/diff[20] ,
		\UUT/Mpath/the_alu/diff[19] ,
		\UUT/Mpath/the_alu/diff[18] ,
		\UUT/Mpath/the_alu/diff[17] ,
		\UUT/Mpath/the_alu/diff[16] ,
		\UUT/Mpath/the_alu/diff[15] ,
		\UUT/Mpath/the_alu/diff[14] ,
		\UUT/Mpath/the_alu/diff[13] ,
		\UUT/Mpath/the_alu/diff[12] ,
		\UUT/Mpath/the_alu/diff[11] ,
		\UUT/Mpath/the_alu/diff[10] ,
		\UUT/Mpath/the_alu/diff[9] ,
		\UUT/Mpath/the_alu/diff[8] ,
		\UUT/Mpath/the_alu/diff[7] ,
		\UUT/Mpath/the_alu/diff[6] ,
		\UUT/Mpath/the_alu/diff[5] ,
		\UUT/Mpath/the_alu/diff[4] ,
		\UUT/Mpath/the_alu/diff[3] ,
		\UUT/Mpath/the_alu/diff[2] ,
		\UUT/Mpath/the_alu/diff[1] ,
		\UUT/Mpath/the_alu/diff[0]  }));
   up_island_DW01_add_3 \UUT/Mpath/the_alu/add_95  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.B({ \UUT/Mpath/out_regB[31] ,
		\UUT/Mpath/out_regB[30] ,
		\UUT/Mpath/out_regB[29] ,
		\UUT/Mpath/out_regB[28] ,
		\UUT/Mpath/out_regB[27] ,
		\UUT/Mpath/out_regB[26] ,
		\UUT/Mpath/out_regB[25] ,
		\UUT/Mpath/out_regB[24] ,
		\UUT/Mpath/out_regB[23] ,
		\UUT/Mpath/out_regB[22] ,
		\UUT/Mpath/out_regB[21] ,
		\UUT/Mpath/out_regB[20] ,
		\UUT/Mpath/out_regB[19] ,
		\UUT/Mpath/out_regB[18] ,
		\UUT/Mpath/out_regB[17] ,
		\UUT/Mpath/out_regB[16] ,
		\UUT/Mpath/out_regB[15] ,
		\UUT/Mpath/out_regB[14] ,
		\UUT/Mpath/out_regB[13] ,
		\UUT/Mpath/out_regB[12] ,
		\UUT/Mpath/out_regB[11] ,
		\UUT/Mpath/out_regB[10] ,
		\UUT/Mpath/out_regB[9] ,
		\UUT/Mpath/out_regB[8] ,
		\UUT/Mpath/out_regB[7] ,
		\UUT/Mpath/out_regB[6] ,
		\UUT/Mpath/out_regB[5] ,
		FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		FE_OFN175_UUT_Mpath_out_regB_1_,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.CI(1'b0), 
	.SUM({ \UUT/Mpath/the_alu/sum[31] ,
		\UUT/Mpath/the_alu/sum[30] ,
		\UUT/Mpath/the_alu/sum[29] ,
		\UUT/Mpath/the_alu/sum[28] ,
		\UUT/Mpath/the_alu/sum[27] ,
		\UUT/Mpath/the_alu/sum[26] ,
		\UUT/Mpath/the_alu/sum[25] ,
		\UUT/Mpath/the_alu/sum[24] ,
		\UUT/Mpath/the_alu/sum[23] ,
		\UUT/Mpath/the_alu/sum[22] ,
		\UUT/Mpath/the_alu/sum[21] ,
		\UUT/Mpath/the_alu/sum[20] ,
		\UUT/Mpath/the_alu/sum[19] ,
		\UUT/Mpath/the_alu/sum[18] ,
		\UUT/Mpath/the_alu/sum[17] ,
		\UUT/Mpath/the_alu/sum[16] ,
		\UUT/Mpath/the_alu/sum[15] ,
		\UUT/Mpath/the_alu/sum[14] ,
		\UUT/Mpath/the_alu/sum[13] ,
		\UUT/Mpath/the_alu/sum[12] ,
		\UUT/Mpath/the_alu/sum[11] ,
		\UUT/Mpath/the_alu/sum[10] ,
		\UUT/Mpath/the_alu/sum[9] ,
		\UUT/Mpath/the_alu/sum[8] ,
		\UUT/Mpath/the_alu/sum[7] ,
		\UUT/Mpath/the_alu/sum[6] ,
		\UUT/Mpath/the_alu/sum[5] ,
		\UUT/Mpath/the_alu/sum[4] ,
		\UUT/Mpath/the_alu/sum[3] ,
		\UUT/Mpath/the_alu/sum[2] ,
		\UUT/Mpath/the_alu/sum[1] ,
		\UUT/Mpath/the_alu/sum[0]  }), 
	.FE_PT1__UUT_Mpath_the_alu_N182_(\UUT/Mpath/the_alu/N182 ), 
	.FE_PT1__UUT_Mpath_the_alu_N183_(\UUT/Mpath/the_alu/N183 ), 
	.FE_PT1__UUT_Mpath_the_alu_N169_(\UUT/Mpath/the_alu/N169 ), 
	.FE_PT1__UUT_Mpath_the_alu_N170_(\UUT/Mpath/the_alu/N170 ), 
	.FE_PT1__UUT_Mpath_the_alu_N164_(\UUT/Mpath/the_alu/N164 ), 
	.FE_PT1__UUT_Mpath_the_alu_N165_(\UUT/Mpath/the_alu/N165 ), 
	.FE_PT1__UUT_Mpath_the_alu_N162_(\UUT/Mpath/the_alu/N162 ), 
	.FE_PT1__UUT_Mpath_the_alu_N171_(\UUT/Mpath/the_alu/N171 ), 
	.FE_PT1__UUT_Mpath_the_alu_N184_(\UUT/Mpath/the_alu/N184 ), 
	.FE_PT1__UUT_Mpath_the_alu_N163_(\UUT/Mpath/the_alu/N163 ), 
	.FE_PT1__UUT_Mpath_the_alu_N172_(\UUT/Mpath/the_alu/N172 ), 
	.FE_PT1__UUT_Mpath_the_alu_N166_(\UUT/Mpath/the_alu/N166 ), 
	.FE_PT1__UUT_Mpath_the_alu_N173_(\UUT/Mpath/the_alu/N173 ), 
	.FE_PT1__UUT_Mpath_the_alu_N167_(\UUT/Mpath/the_alu/N167 ), 
	.FE_PT1__UUT_Mpath_the_alu_N174_(\UUT/Mpath/the_alu/N174 ), 
	.FE_PT1__UUT_Mpath_the_alu_N168_(\UUT/Mpath/the_alu/N168 ), 
	.FE_PT1__UUT_Mpath_the_alu_N175_(\UUT/Mpath/the_alu/N175 ), 
	.FE_PT1__UUT_Mpath_the_alu_N159_(\UUT/Mpath/the_alu/N159 ), 
	.FE_PT1__UUT_Mpath_the_alu_N176_(\UUT/Mpath/the_alu/N176 ), 
	.FE_PT1__UUT_Mpath_the_alu_N177_(\UUT/Mpath/the_alu/N177 ), 
	.FE_PT1__UUT_Mpath_the_alu_N178_(\UUT/Mpath/the_alu/N178 ), 
	.FE_OFN181_UUT_Mpath_out_regB_0_(FE_OFN185_UUT_Mpath_out_regB_0_));
   up_island_DW_mult_tc_1 \UUT/Mpath/the_mult/mult_186  (.a({ FE_OFN177_UUT_Mpath_the_mult_x_operand1_31_,
		\UUT/Mpath/the_mult/x_operand1[30] ,
		FE_OFN113_UUT_Mpath_the_mult_x_operand1_29_,
		\UUT/Mpath/the_mult/x_operand1[28] ,
		FE_OFN117_UUT_Mpath_the_mult_x_operand1_27_,
		\UUT/Mpath/the_mult/x_operand1[26] ,
		FE_OFN121_UUT_Mpath_the_mult_x_operand1_25_,
		\UUT/Mpath/the_mult/x_operand1[24] ,
		FE_OFN173_UUT_Mpath_the_mult_x_operand1_23_,
		\UUT/Mpath/the_mult/x_operand1[22] ,
		FE_OFCN204_FE_OFN126_UUT_Mpath_the_mult_x_operand1_21_,
		\UUT/Mpath/the_mult/x_operand1[20] ,
		FE_OFN130_UUT_Mpath_the_mult_x_operand1_19_,
		\UUT/Mpath/the_mult/x_operand1[18] ,
		FE_OFN134_UUT_Mpath_the_mult_x_operand1_17_,
		\UUT/Mpath/the_mult/x_operand1[16] ,
		FE_OFN138_UUT_Mpath_the_mult_x_operand1_15_,
		\UUT/Mpath/the_mult/x_operand1[14] ,
		FE_OFN142_UUT_Mpath_the_mult_x_operand1_13_,
		\UUT/Mpath/the_mult/x_operand1[12] ,
		FE_OFN146_UUT_Mpath_the_mult_x_operand1_11_,
		\UUT/Mpath/the_mult/x_operand1[10] ,
		FE_OFN149_UUT_Mpath_the_mult_x_operand1_9_,
		\UUT/Mpath/the_mult/x_operand1[8] ,
		FE_OFN152_UUT_Mpath_the_mult_x_operand1_7_,
		\UUT/Mpath/the_mult/x_operand1[6] ,
		FE_OFN156_UUT_Mpath_the_mult_x_operand1_5_,
		\UUT/Mpath/the_mult/x_operand1[4] ,
		FE_OFN165_UUT_Mpath_the_mult_x_operand1_3_,
		\UUT/Mpath/the_mult/x_operand1[2] ,
		FE_OFN171_UUT_Mpath_the_mult_x_operand1_1_,
		\UUT/Mpath/the_mult/x_operand1[0]  }), 
	.b({ \UUT/Mpath/the_mult/x_operand2 [31],
		\UUT/Mpath/the_mult/x_operand2 [30],
		\UUT/Mpath/the_mult/x_operand2 [29],
		\UUT/Mpath/the_mult/x_operand2 [28],
		\UUT/Mpath/the_mult/x_operand2 [27],
		\UUT/Mpath/the_mult/x_operand2 [26],
		FE_OFN120_UUT_Mpath_the_mult_x_operand2_25_,
		\UUT/Mpath/the_mult/x_operand2 [24],
		\UUT/Mpath/the_mult/x_operand2 [23],
		\UUT/Mpath/the_mult/x_operand2 [22],
		\UUT/Mpath/the_mult/x_operand2 [21],
		\UUT/Mpath/the_mult/x_operand2 [20],
		FE_OFN129_UUT_Mpath_the_mult_x_operand2_19_,
		\UUT/Mpath/the_mult/x_operand2 [18],
		FE_OFN133_UUT_Mpath_the_mult_x_operand2_17_,
		FE_OFN136_UUT_Mpath_the_mult_x_operand2_16_,
		FE_OFN137_UUT_Mpath_the_mult_x_operand2_15_,
		FE_OFN140_UUT_Mpath_the_mult_x_operand2_14_,
		\UUT/Mpath/the_mult/x_operand2 [13],
		\UUT/Mpath/the_mult/x_operand2 [12],
		\UUT/Mpath/the_mult/x_operand2 [11],
		\UUT/Mpath/the_mult/x_operand2 [10],
		\UUT/Mpath/the_mult/x_operand2 [9],
		\UUT/Mpath/the_mult/x_operand2 [8],
		\UUT/Mpath/the_mult/x_operand2 [7],
		\UUT/Mpath/the_mult/x_operand2 [6],
		\UUT/Mpath/the_mult/x_operand2 [5],
		\UUT/Mpath/the_mult/x_operand2 [4],
		\UUT/Mpath/the_mult/x_operand2 [3],
		FE_OFN167_UUT_Mpath_the_mult_x_operand2_2_,
		FE_OFN170_UUT_Mpath_the_mult_x_operand2_1_,
		FE_OFN105_UUT_Mpath_the_mult_x_operand2_0_ }), 
	.product({ \UUT/Mpath/the_mult/x_mult_out[63] ,
		\UUT/Mpath/the_mult/x_mult_out[62] ,
		\UUT/Mpath/the_mult/x_mult_out[61] ,
		\UUT/Mpath/the_mult/x_mult_out[60] ,
		\UUT/Mpath/the_mult/x_mult_out[59] ,
		\UUT/Mpath/the_mult/x_mult_out[58] ,
		\UUT/Mpath/the_mult/x_mult_out[57] ,
		\UUT/Mpath/the_mult/x_mult_out[56] ,
		\UUT/Mpath/the_mult/x_mult_out[55] ,
		\UUT/Mpath/the_mult/x_mult_out[54] ,
		\UUT/Mpath/the_mult/x_mult_out[53] ,
		\UUT/Mpath/the_mult/x_mult_out[52] ,
		\UUT/Mpath/the_mult/x_mult_out[51] ,
		\UUT/Mpath/the_mult/x_mult_out[50] ,
		\UUT/Mpath/the_mult/x_mult_out[49] ,
		\UUT/Mpath/the_mult/x_mult_out[48] ,
		\UUT/Mpath/the_mult/x_mult_out[47] ,
		\UUT/Mpath/the_mult/x_mult_out[46] ,
		\UUT/Mpath/the_mult/x_mult_out[45] ,
		\UUT/Mpath/the_mult/x_mult_out[44] ,
		\UUT/Mpath/the_mult/x_mult_out[43] ,
		\UUT/Mpath/the_mult/x_mult_out[42] ,
		\UUT/Mpath/the_mult/x_mult_out[41] ,
		\UUT/Mpath/the_mult/x_mult_out[40] ,
		\UUT/Mpath/the_mult/x_mult_out[39] ,
		\UUT/Mpath/the_mult/x_mult_out[38] ,
		\UUT/Mpath/the_mult/x_mult_out[37] ,
		\UUT/Mpath/the_mult/x_mult_out[36] ,
		\UUT/Mpath/the_mult/x_mult_out[35] ,
		\UUT/Mpath/the_mult/x_mult_out[34] ,
		\UUT/Mpath/the_mult/x_mult_out[33] ,
		\UUT/Mpath/the_mult/x_mult_out[32] ,
		\UUT/Mpath/the_mult/x_mult_out[31] ,
		\UUT/Mpath/the_mult/x_mult_out[30] ,
		\UUT/Mpath/the_mult/x_mult_out[29] ,
		\UUT/Mpath/the_mult/x_mult_out[28] ,
		\UUT/Mpath/the_mult/x_mult_out[27] ,
		\UUT/Mpath/the_mult/x_mult_out[26] ,
		\UUT/Mpath/the_mult/x_mult_out[25] ,
		\UUT/Mpath/the_mult/x_mult_out[24] ,
		\UUT/Mpath/the_mult/x_mult_out[23] ,
		\UUT/Mpath/the_mult/x_mult_out[22] ,
		\UUT/Mpath/the_mult/x_mult_out[21] ,
		\UUT/Mpath/the_mult/x_mult_out[20] ,
		\UUT/Mpath/the_mult/x_mult_out[19] ,
		\UUT/Mpath/the_mult/x_mult_out[18] ,
		\UUT/Mpath/the_mult/x_mult_out[17] ,
		\UUT/Mpath/the_mult/x_mult_out[16] ,
		\UUT/Mpath/the_mult/x_mult_out[15] ,
		\UUT/Mpath/the_mult/x_mult_out[14] ,
		\UUT/Mpath/the_mult/x_mult_out[13] ,
		\UUT/Mpath/the_mult/x_mult_out[12] ,
		\UUT/Mpath/the_mult/x_mult_out[11] ,
		\UUT/Mpath/the_mult/x_mult_out[10] ,
		\UUT/Mpath/the_mult/x_mult_out[9] ,
		\UUT/Mpath/the_mult/x_mult_out[8] ,
		\UUT/Mpath/the_mult/x_mult_out[7] ,
		\UUT/Mpath/the_mult/x_mult_out[6] ,
		\UUT/Mpath/the_mult/x_mult_out[5] ,
		\UUT/Mpath/the_mult/x_mult_out[4] ,
		\UUT/Mpath/the_mult/x_mult_out[3] ,
		\UUT/Mpath/the_mult/x_mult_out[2] ,
		\UUT/Mpath/the_mult/x_mult_out[1] ,
		\UUT/Mpath/the_mult/x_mult_out[0]  }), 
	.FE_PT1_n796(n796), 
	.FE_PT1_n705(n705), 
	.FE_PT1_n654(n654), 
	.FE_PT1_n617(n617), 
	.FE_PT1_n582(n582), 
	.n531(n531), 
	.FE_PT1_n477(n477), 
	.n338(n338), 
	.FE_PT1_n808(n808), 
	.FE_PT1_n949(n949));
   up_island_DW_rightsh_1 \UUT/Mpath/the_shift/S_SRL/srl_128  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.SH({ FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		\UUT/Mpath/out_regB[1] ,
		FE_OFN184_UUT_Mpath_out_regB_0_ }), 
	.B(\UUT/Mpath/the_shift/sh_srl ), 
	.DATA_TC(1'b0), 
	.FE_OFN169_UUT_Mpath_out_regB_2_(FE_OFN169_UUT_Mpath_out_regB_2_), 
	.FE_OFN175_UUT_Mpath_out_regB_1_(FE_OFN175_UUT_Mpath_out_regB_1_), 
	.FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_(FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_));
   up_island_DW_sra_1 \UUT/Mpath/the_shift/S_SRA/sra_106  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.SH({ FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN163_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.B(\UUT/Mpath/the_shift/sh_sra ), 
	.SH_TC(1'b0), 
	.FE_OFN160_UUT_Mpath_out_regB_4_(FE_OFN160_UUT_Mpath_out_regB_4_), 
	.FE_OFN164_UUT_Mpath_out_regB_3_(FE_OFN164_UUT_Mpath_out_regB_3_), 
	.FE_OFN180_UUT_Mpath_out_regB_0_(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.FE_OFN181_UUT_Mpath_out_regB_0_(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.FE_OFN184_UUT_Mpath_out_regB_0_(FE_OFN184_UUT_Mpath_out_regB_0_), 
	.FE_OFN185_UUT_Mpath_out_regB_0_(FE_OFN185_UUT_Mpath_out_regB_0_), 
	.FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_(FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_));
   up_island_DW_rbsh_1 \UUT/Mpath/the_shift/S_ROR/ror_81  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.SH({ FE_OFN160_UUT_Mpath_out_regB_4_,
		FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_,
		FE_OFN169_UUT_Mpath_out_regB_2_,
		FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_,
		FE_OFN185_UUT_Mpath_out_regB_0_ }), 
	.B(\UUT/Mpath/the_shift/sh_ror ), 
	.SH_TC(1'b0), 
	.FE_OFN176_UUT_Mpath_out_regB_1_(FE_OFN176_UUT_Mpath_out_regB_1_), 
	.FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_(FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_), 
	.FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_));
   up_island_DW01_bsh_1 \UUT/Mpath/the_shift/S_ROL/rol_55  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.SH({ FE_OFN160_UUT_Mpath_out_regB_4_,
		FE_OFCN202_FE_OFN164_UUT_Mpath_out_regB_3_,
		FE_OFN169_UUT_Mpath_out_regB_2_,
		FE_OFCN201_FE_OFN176_UUT_Mpath_out_regB_1_,
		FE_OFN185_UUT_Mpath_out_regB_0_ }), 
	.B(\UUT/Mpath/the_shift/sh_rol ), 
	.FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_(FE_OFCN203_FE_OFN160_UUT_Mpath_out_regB_4_));
   up_island_DW_leftsh_1 \UUT/Mpath/the_shift/S_SLL/sll_150  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.SH({ FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.B(\UUT/Mpath/the_shift/sh_sll ), 
	.FE_OFN163_UUT_Mpath_out_regB_3_(FE_OFN163_UUT_Mpath_out_regB_3_), 
	.FE_OFN180_UUT_Mpath_out_regB_0_(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.FE_OFN184_UUT_Mpath_out_regB_0_(FE_OFN184_UUT_Mpath_out_regB_0_));
   up_island_DW_cmp_0 \UUT/Mpath/the_alu/lt_114  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.B({ \UUT/Mpath/out_regB[31] ,
		\UUT/Mpath/out_regB[30] ,
		\UUT/Mpath/out_regB[29] ,
		\UUT/Mpath/out_regB[28] ,
		\UUT/Mpath/out_regB[27] ,
		\UUT/Mpath/out_regB[26] ,
		\UUT/Mpath/out_regB[25] ,
		\UUT/Mpath/out_regB[24] ,
		\UUT/Mpath/out_regB[23] ,
		\UUT/Mpath/out_regB[22] ,
		\UUT/Mpath/out_regB[21] ,
		\UUT/Mpath/out_regB[20] ,
		\UUT/Mpath/out_regB[19] ,
		\UUT/Mpath/out_regB[18] ,
		\UUT/Mpath/out_regB[17] ,
		\UUT/Mpath/out_regB[16] ,
		\UUT/Mpath/out_regB[15] ,
		\UUT/Mpath/out_regB[14] ,
		\UUT/Mpath/out_regB[13] ,
		\UUT/Mpath/out_regB[12] ,
		\UUT/Mpath/out_regB[11] ,
		\UUT/Mpath/out_regB[10] ,
		\UUT/Mpath/out_regB[9] ,
		\UUT/Mpath/out_regB[8] ,
		\UUT/Mpath/out_regB[7] ,
		\UUT/Mpath/out_regB[6] ,
		\UUT/Mpath/out_regB[5] ,
		FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.TC(1'b1), 
	.GE_LT(1'b1), 
	.GE_GT_EQ(1'b0), 
	.GE_LT_GT_LE(\UUT/Mpath/the_alu/N91 ));
   up_island_DW_cmp_1 \UUT/Mpath/the_alu/lt_120  (.A({ \UUT/Mpath/out_regA[31] ,
		\UUT/Mpath/out_regA[30] ,
		\UUT/Mpath/out_regA[29] ,
		\UUT/Mpath/out_regA[28] ,
		\UUT/Mpath/out_regA[27] ,
		\UUT/Mpath/out_regA[26] ,
		\UUT/Mpath/out_regA[25] ,
		\UUT/Mpath/out_regA[24] ,
		\UUT/Mpath/out_regA[23] ,
		\UUT/Mpath/out_regA[22] ,
		\UUT/Mpath/out_regA[21] ,
		\UUT/Mpath/out_regA[20] ,
		\UUT/Mpath/out_regA[19] ,
		\UUT/Mpath/out_regA[18] ,
		\UUT/Mpath/out_regA[17] ,
		\UUT/Mpath/out_regA[16] ,
		\UUT/Mpath/out_regA[15] ,
		\UUT/Mpath/out_regA[14] ,
		\UUT/Mpath/out_regA[13] ,
		\UUT/Mpath/out_regA[12] ,
		\UUT/Mpath/out_regA[11] ,
		\UUT/Mpath/out_regA[10] ,
		\UUT/Mpath/out_regA[9] ,
		\UUT/Mpath/out_regA[8] ,
		\UUT/Mpath/out_regA[7] ,
		\UUT/Mpath/out_regA[6] ,
		\UUT/Mpath/out_regA[5] ,
		\UUT/Mpath/out_regA[4] ,
		\UUT/Mpath/out_regA[3] ,
		FE_OFCN198_UUT_Mpath_out_regA_2_,
		\UUT/Mpath/out_regA[1] ,
		FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_ }), 
	.B({ \UUT/Mpath/out_regB[31] ,
		\UUT/Mpath/out_regB[30] ,
		\UUT/Mpath/out_regB[29] ,
		\UUT/Mpath/out_regB[28] ,
		\UUT/Mpath/out_regB[27] ,
		\UUT/Mpath/out_regB[26] ,
		\UUT/Mpath/out_regB[25] ,
		\UUT/Mpath/out_regB[24] ,
		\UUT/Mpath/out_regB[23] ,
		\UUT/Mpath/out_regB[22] ,
		\UUT/Mpath/out_regB[21] ,
		\UUT/Mpath/out_regB[20] ,
		\UUT/Mpath/out_regB[19] ,
		\UUT/Mpath/out_regB[18] ,
		\UUT/Mpath/out_regB[17] ,
		\UUT/Mpath/out_regB[16] ,
		\UUT/Mpath/out_regB[15] ,
		\UUT/Mpath/out_regB[14] ,
		\UUT/Mpath/out_regB[13] ,
		\UUT/Mpath/out_regB[12] ,
		\UUT/Mpath/out_regB[11] ,
		\UUT/Mpath/out_regB[10] ,
		\UUT/Mpath/out_regB[9] ,
		\UUT/Mpath/out_regB[8] ,
		\UUT/Mpath/out_regB[7] ,
		\UUT/Mpath/out_regB[6] ,
		\UUT/Mpath/out_regB[5] ,
		FE_OFN159_UUT_Mpath_out_regB_4_,
		FE_OFN162_UUT_Mpath_out_regB_3_,
		FE_OFN168_UUT_Mpath_out_regB_2_,
		FE_OFCN200_FE_OFN175_UUT_Mpath_out_regB_1_,
		FE_OFN182_UUT_Mpath_out_regB_0_ }), 
	.TC(1'b0), 
	.GE_LT(1'b1), 
	.GE_GT_EQ(1'b0), 
	.GE_LT_GT_LE(\UUT/Mpath/the_alu/N93 ));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N49 ), 
	.Q(\UUT/Mpath/out_regA[17] ), 
	.D(n3169), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N37 ), 
	.Q(\UUT/Mpath/out_regA[23] ), 
	.D(n3776), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N44 ), 
	.Q(\UUT/Mpath/out_regB[20] ), 
	.D(n3044), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[20]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N43 ), 
	.Q(\UUT/Mpath/out_regA[20] ), 
	.D(n3049), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N46 ), 
	.Q(\UUT/Mpath/out_regB[19] ), 
	.D(n3084), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[19]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N45 ), 
	.Q(\UUT/Mpath/out_regA[19] ), 
	.D(n3089), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[7]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N69 ), 
	.Q(\UUT/Mpath/out_regA[7] ), 
	.D(n3501), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[8]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N67 ), 
	.Q(\UUT/Mpath/out_regA[8] ), 
	.D(n3492), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N55 ), 
	.Q(\UUT/Mpath/out_regA[14] ), 
	.D(n3289), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[29]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N25 ), 
	.Q(\UUT/Mpath/out_regA[29] ), 
	.D(n3943), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N57 ), 
	.Q(\UUT/Mpath/out_regA[13] ), 
	.D(n3329), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N34 ), 
	.Q(\UUT/Mpath/out_regB[25] ), 
	.D(n2918), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[25]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N33 ), 
	.Q(\UUT/Mpath/out_regA[25] ), 
	.D(n3811), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N36 ), 
	.Q(\UUT/Mpath/out_regB[24] ), 
	.D(n2924), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[24]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N35 ), 
	.Q(\UUT/Mpath/out_regA[24] ), 
	.D(n2929), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N30 ), 
	.Q(\UUT/Mpath/out_regB[27] ), 
	.D(n2906), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[27]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N29 ), 
	.Q(\UUT/Mpath/out_regA[27] ), 
	.D(n3877), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[6]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N71 ), 
	.Q(\UUT/Mpath/out_regA[6] ), 
	.D(n3541), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N59 ), 
	.Q(\UUT/Mpath/out_regA[12] ), 
	.D(n3369), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[30]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N23 ), 
	.Q(\UUT/Mpath/out_regA[30] ), 
	.D(n3981), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N48 ), 
	.Q(\UUT/Mpath/out_regB[18] ), 
	.D(n3124), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[18]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N47 ), 
	.Q(\UUT/Mpath/out_regA[18] ), 
	.D(n3129), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regA/data_out_reg[2]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N79 ), 
	.Q(\UUT/Mpath/out_regA[2] ), 
	.D(n3701), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N74 ), 
	.Q(\UUT/Mpath/out_regB[5] ), 
	.D(n3576), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[5]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N73 ), 
	.Q(\UUT/Mpath/out_regA[5] ), 
	.D(n3581), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N32 ), 
	.Q(\UUT/Mpath/out_regB[26] ), 
	.D(n2912), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[26]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N31 ), 
	.Q(\UUT/Mpath/out_regA[26] ), 
	.D(n3844), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[17]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N50 ), 
	.Q(\UUT/Mpath/out_regB[17] ), 
	.D(n3164), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[23]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N38 ), 
	.Q(\UUT/Mpath/out_regB[23] ), 
	.D(n4014), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N28 ), 
	.Q(\UUT/Mpath/out_regB[28] ), 
	.D(n2900), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[28]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N27 ), 
	.Q(\UUT/Mpath/out_regA[28] ), 
	.D(n3910), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[3]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N77 ), 
	.Q(\UUT/Mpath/out_regA[3] ), 
	.D(n3661), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[10]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N63 ), 
	.Q(\UUT/Mpath/out_regA[10] ), 
	.D(n3446), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[9]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N65 ), 
	.Q(\UUT/Mpath/out_regA[9] ), 
	.D(n3454), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N22 ), 
	.Q(\UUT/Mpath/out_regB[31] ), 
	.D(n4327), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N21 ), 
	.Q(\UUT/Mpath/out_regA[31] ), 
	.D(n4057), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[4]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N75 ), 
	.Q(\UUT/Mpath/out_regA[4] ), 
	.D(n3621), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N52 ), 
	.Q(\UUT/Mpath/out_regB[16] ), 
	.D(n3204), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[16]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N51 ), 
	.Q(\UUT/Mpath/out_regA[16] ), 
	.D(n3209), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N40 ), 
	.Q(\UUT/Mpath/out_regB[22] ), 
	.D(n2964), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[22]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N39 ), 
	.Q(\UUT/Mpath/out_regA[22] ), 
	.D(n2969), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N61 ), 
	.Q(\UUT/Mpath/out_regA[11] ), 
	.D(n3409), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N41 ), 
	.Q(\UUT/Mpath/out_regA[21] ), 
	.D(n3009), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N54 ), 
	.Q(\UUT/Mpath/out_regB[15] ), 
	.D(n3244), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regA/data_out_reg[15]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N53 ), 
	.Q(\UUT/Mpath/out_regA[15] ), 
	.D(n3249), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[21]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N42 ), 
	.Q(\UUT/Mpath/out_regB[21] ), 
	.D(n3004), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/the_mult/Pipe_mult_reg/data_out_reg[50]  (.RN(\UUT/Mcontrol/int_reset ), 
	.Q(\UUT/Mpath/the_mult/Mult_out[50] ), 
	.D(n4307), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[14]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N56 ), 
	.Q(\UUT/Mpath/out_regB[14] ), 
	.D(n3284), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[13]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N58 ), 
	.Q(\UUT/Mpath/out_regB[13] ), 
	.D(n3324), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[12]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N60 ), 
	.Q(\UUT/Mpath/out_regB[12] ), 
	.D(n3364), 
	.CK(CLK));
   DFFR_X2 \UUT/Mpath/regB/data_out_reg[11]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N62 ), 
	.Q(\UUT/Mpath/out_regB[11] ), 
	.D(n3404), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regA/data_out_reg[0]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N83 ), 
	.Q(\UUT/Mpath/out_regA[0] ), 
	.D(n4256), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/regA/data_out_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(\UUT/Mpath/the_alu/N81 ), 
	.Q(\UUT/Mpath/out_regA[1] ), 
	.D(n3740), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[5]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2685), 
	.Q(\UUT/Mcontrol/f_currpc [5]), 
	.D(n3574), 
	.CK(CLK));
   DFFS_X2 \UUT/Mcontrol/Program_counter/out_pc_reg[18]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2651), 
	.Q(\UUT/Mcontrol/f_currpc [18]), 
	.D(n3123), 
	.CK(CLK));
   DFFR_X1 \UUT/Mpath/the_mult/MulHi_reg/data_out_reg[31]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n5685), 
	.Q(\UUT/Mpath/the_mult/acc_out[63] ), 
	.D(n4329), 
	.CK(CLK));
   NAND2_X1 syn1555 (.ZN(n6440), 
	.A2(\UUT/Mpath/the_mult/N231 ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[0] ));
   INV_X4 syn1525 (.ZN(net54953), 
	.A(n6445));
   NAND3_X1 syn1524 (.ZN(n6445), 
	.A3(\localbus/N95 ), 
	.A2(n6444), 
	.A1(n6436));
   NAND2_X1 syn1522 (.ZN(n6444), 
	.A2(\localbus/N322 ), 
	.A1(\localbus/N335 ));
   INV_X2 syn868 (.ZN(n139), 
	.A(n6433));
   INV_X1 syn831 (.ZN(n6438), 
	.A(\UUT/Mpath/the_mult/m_mul_command[3] ));
   INV_X2 syn768 (.ZN(n137), 
	.A(n6443));
   NAND2_X1 syn767 (.ZN(n6443), 
	.A2(n6432), 
	.A1(n975));
   NOR2_X1 syn749 (.ZN(n6435), 
	.A2(n6432), 
	.A1(n6426));
   NOR2_X1 syn745 (.ZN(n6434), 
	.A2(net54953), 
	.A1(n6429));
   AND2_X1 syn743 (.ZN(n6430), 
	.A2(n6440), 
	.A1(n6439));
   NOR2_X1 syn741 (.ZN(n6439), 
	.A2(\UUT/Mpath/the_mult/m_mul_command[1] ), 
	.A1(\UUT/Mpath/the_mult/N244 ));
   AND2_X1 syn739 (.ZN(n6431), 
	.A2(n6438), 
	.A1(n6437));
   NOR2_X1 syn737 (.ZN(n6437), 
	.A2(\UUT/Mpath/the_mult/m_mul_command[5] ), 
	.A1(\UUT/Mpath/the_mult/m_mul_command[4] ));
   INV_X1 syn727 (.ZN(n6428), 
	.A(net87679));
   NAND3_X1 syn725 (.ZN(n6433), 
	.A3(n971), 
	.A2(n6435), 
	.A1(n6434));
   INV_X1 syn722 (.ZN(n6432), 
	.A(\UUT/Mpath/the_mult/N285 ));
   NAND2_X1 syn721 (.ZN(n6426), 
	.A2(n6431), 
	.A1(n6430));
   INV_X1 syn720 (.ZN(n6429), 
	.A(n5413));
   NAND3_X1 net89067 (.ZN(n1183), 
	.A3(n971), 
	.A2(n6426), 
	.A1(\UUT/Mpath/the_mult/N285 ));
   DFFR_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[1]  (.RN(\UUT/Mcontrol/int_reset ), 
	.QN(n2698), 
	.Q(\UUT/Mcontrol/f_currpc [1]), 
	.D(n3735), 
	.CK(CLK));
   DFFS_X1 \UUT/Mcontrol/Program_counter/out_pc_reg[15]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n2660), 
	.Q(\UUT/Mcontrol/f_currpc [15]), 
	.D(n3243), 
	.CK(CLK));
   DFFS_X2 \UUT/Mcontrol/ir_xm/out_mem_command_reg[MR]  (.SN(\UUT/Mcontrol/int_reset ), 
	.QN(n5710), 
	.Q(\UUT/m_mem_command[MR] ), 
	.D(n4060), 
	.CK(CLK));
   NOR2_X1 U5278 (.ZN(n6436), 
	.A2(BUS_NREADY), 
	.A1(\localbus/c2_op[MASTER] ));
   INV_X1 U5279 (.ZN(n6868), 
	.A(\UUT/branch_rega [4]));
   OR2_X1 U5281 (.ZN(n6787), 
	.A2(\UUT/branch_rega [4]), 
	.A1(n6794));
   NOR3_X2 U5282 (.ZN(n2074), 
	.A3(n2070), 
	.A2(n6209), 
	.A1(n933));
   NAND2_X2 U5283 (.ZN(n71), 
	.A2(n175), 
	.A1(n147));
   OR2_X1 U5284 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N116 ), 
	.A2(\UUT/Mcontrol/st_logic/N106 ), 
	.A1(\UUT/Mcontrol/d_jump_type[1] ));
   OR2_X1 U5285 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N264 ), 
	.A2(\UUT/Mcontrol/st_logic/N61 ), 
	.A1(\UUT/Mcontrol/d_jump_type[1] ));
   OR2_X1 U5286 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N252 ), 
	.A2(\UUT/Mcontrol/st_logic/N86 ), 
	.A1(\UUT/Mcontrol/d_jump_type[1] ));
   INV_X1 U5289 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N224 ), 
	.A(\UUT/Mcontrol/d_jump_type[1] ));
   NOR2_X1 U5298 (.ZN(\UUT/rs1_addr [1]), 
	.A2(n6322), 
	.A1(n5896));
   INV_X1 U5299 (.ZN(n6854), 
	.A(\UUT/branch_rega [5]));
   INV_X1 U5300 (.ZN(n6832), 
	.A(\UUT/branch_rega [0]));
   AND2_X1 U5302 (.ZN(\UUT/Mpath/the_alu/N107 ), 
	.A2(\UUT/Mpath/out_regB[18] ), 
	.A1(\UUT/Mpath/out_regA[18] ));
   OR2_X1 U5303 (.ZN(\UUT/Mpath/the_alu/N139 ), 
	.A2(\UUT/Mpath/out_regB[18] ), 
	.A1(\UUT/Mpath/out_regA[18] ));
   AND2_X2 U5304 (.ZN(n6347), 
	.A2(\UUT/N3 ), 
	.A1(\localbus/N50 ));
   INV_X1 U5305 (.ZN(\localbus/N50 ), 
	.A(\localbus/c1_op[MASTER] ));
   AND2_X1 U5306 (.ZN(\UUT/Mpath/the_alu/N110 ), 
	.A2(\UUT/Mpath/out_regB[15] ), 
	.A1(\UUT/Mpath/out_regA[15] ));
   OR2_X1 U5307 (.ZN(\UUT/Mpath/the_alu/N142 ), 
	.A2(\UUT/Mpath/out_regB[15] ), 
	.A1(\UUT/Mpath/out_regA[15] ));
   AND2_X1 U5308 (.ZN(\UUT/Mpath/the_alu/N106 ), 
	.A2(\UUT/Mpath/out_regB[19] ), 
	.A1(\UUT/Mpath/out_regA[19] ));
   OR2_X1 U5309 (.ZN(\UUT/Mpath/the_alu/N138 ), 
	.A2(\UUT/Mpath/out_regB[19] ), 
	.A1(\UUT/Mpath/out_regA[19] ));
   AND2_X1 U5310 (.ZN(\UUT/Mpath/the_alu/N105 ), 
	.A2(\UUT/Mpath/out_regB[20] ), 
	.A1(\UUT/Mpath/out_regA[20] ));
   OR2_X1 U5311 (.ZN(\UUT/Mpath/the_alu/N137 ), 
	.A2(\UUT/Mpath/out_regB[20] ), 
	.A1(\UUT/Mpath/out_regA[20] ));
   AND2_X1 U5312 (.ZN(\UUT/Mpath/the_alu/N104 ), 
	.A2(\UUT/Mpath/out_regB[21] ), 
	.A1(\UUT/Mpath/out_regA[21] ));
   OR2_X1 U5313 (.ZN(\UUT/Mpath/the_alu/N136 ), 
	.A2(\UUT/Mpath/out_regB[21] ), 
	.A1(\UUT/Mpath/out_regA[21] ));
   AND2_X1 U5314 (.ZN(\UUT/Mpath/the_alu/N116 ), 
	.A2(\UUT/Mpath/out_regB[9] ), 
	.A1(\UUT/Mpath/out_regA[9] ));
   OR2_X1 U5315 (.ZN(\UUT/Mpath/the_alu/N148 ), 
	.A2(\UUT/Mpath/out_regB[9] ), 
	.A1(\UUT/Mpath/out_regA[9] ));
   AND2_X1 U5316 (.ZN(\UUT/Mpath/the_alu/N115 ), 
	.A2(\UUT/Mpath/out_regB[10] ), 
	.A1(\UUT/Mpath/out_regA[10] ));
   OR2_X1 U5317 (.ZN(\UUT/Mpath/the_alu/N147 ), 
	.A2(\UUT/Mpath/out_regB[10] ), 
	.A1(\UUT/Mpath/out_regA[10] ));
   AND2_X1 U5318 (.ZN(\UUT/Mpath/the_alu/N103 ), 
	.A2(\UUT/Mpath/out_regB[22] ), 
	.A1(\UUT/Mpath/out_regA[22] ));
   OR2_X1 U5319 (.ZN(\UUT/Mpath/the_alu/N135 ), 
	.A2(\UUT/Mpath/out_regB[22] ), 
	.A1(\UUT/Mpath/out_regA[22] ));
   OAI21_X1 U5321 (.ZN(n5529), 
	.B2(n2592), 
	.B1(\UUT/regfile/N262 ), 
	.A(\UUT/Mcontrol/st_logic/N55 ));
   AND3_X2 U5322 (.ZN(n135), 
	.A3(n5413), 
	.A2(net54895), 
	.A1(n1183));
   AND2_X1 U5323 (.ZN(\UUT/Mpath/the_alu/N102 ), 
	.A2(\UUT/Mpath/out_regB[23] ), 
	.A1(\UUT/Mpath/out_regA[23] ));
   OR2_X1 U5324 (.ZN(\UUT/Mpath/the_alu/N134 ), 
	.A2(\UUT/Mpath/out_regB[23] ), 
	.A1(\UUT/Mpath/out_regA[23] ));
   AND2_X2 U5325 (.ZN(n1215), 
	.A2(n2574), 
	.A1(\UUT/Mpath/the_alu/N474 ));
   AND2_X2 U5326 (.ZN(n1213), 
	.A2(\UUT/Mpath/the_alu/N492 ), 
	.A1(n6348));
   AND2_X1 U5327 (.ZN(\UUT/Mpath/the_alu/N117 ), 
	.A2(\UUT/Mpath/out_regB[8] ), 
	.A1(\UUT/Mpath/out_regA[8] ));
   OR2_X1 U5328 (.ZN(\UUT/Mpath/the_alu/N149 ), 
	.A2(\UUT/Mpath/out_regB[8] ), 
	.A1(\UUT/Mpath/out_regA[8] ));
   AND2_X1 U5329 (.ZN(\UUT/Mpath/the_alu/N109 ), 
	.A2(\UUT/Mpath/out_regB[16] ), 
	.A1(\UUT/Mpath/out_regA[16] ));
   OR2_X1 U5330 (.ZN(\UUT/Mpath/the_alu/N141 ), 
	.A2(\UUT/Mpath/out_regB[16] ), 
	.A1(\UUT/Mpath/out_regA[16] ));
   AND2_X1 U5331 (.ZN(\UUT/Mpath/the_alu/N108 ), 
	.A2(\UUT/Mpath/out_regB[17] ), 
	.A1(\UUT/Mpath/out_regA[17] ));
   OR2_X1 U5332 (.ZN(\UUT/Mpath/the_alu/N140 ), 
	.A2(\UUT/Mpath/out_regB[17] ), 
	.A1(\UUT/Mpath/out_regA[17] ));
   AND2_X1 U5333 (.ZN(\UUT/Mpath/the_alu/N97 ), 
	.A2(\UUT/Mpath/out_regB[28] ), 
	.A1(\UUT/Mpath/out_regA[28] ));
   OR2_X1 U5334 (.ZN(\UUT/Mpath/the_alu/N129 ), 
	.A2(\UUT/Mpath/out_regB[28] ), 
	.A1(\UUT/Mpath/out_regA[28] ));
   AND2_X1 U5335 (.ZN(\UUT/Mpath/the_alu/N98 ), 
	.A2(\UUT/Mpath/out_regB[27] ), 
	.A1(\UUT/Mpath/out_regA[27] ));
   OR2_X1 U5336 (.ZN(\UUT/Mpath/the_alu/N130 ), 
	.A2(\UUT/Mpath/out_regB[27] ), 
	.A1(\UUT/Mpath/out_regA[27] ));
   AND2_X1 U5337 (.ZN(\UUT/Mpath/the_alu/N100 ), 
	.A2(\UUT/Mpath/out_regB[25] ), 
	.A1(\UUT/Mpath/out_regA[25] ));
   OR2_X1 U5338 (.ZN(\UUT/Mpath/the_alu/N132 ), 
	.A2(\UUT/Mpath/out_regB[25] ), 
	.A1(\UUT/Mpath/out_regA[25] ));
   AND2_X1 U5339 (.ZN(\UUT/Mpath/the_alu/N95 ), 
	.A2(\UUT/Mpath/out_regB[30] ), 
	.A1(\UUT/Mpath/out_regA[30] ));
   OR2_X1 U5340 (.ZN(\UUT/Mpath/the_alu/N127 ), 
	.A2(\UUT/Mpath/out_regB[30] ), 
	.A1(\UUT/Mpath/out_regA[30] ));
   OR2_X2 U5341 (.ZN(n132), 
	.A2(\UUT/regfile/N269 ), 
	.A1(\UUT/byp_controlB[2] ));
   AND3_X2 U5342 (.ZN(n142), 
	.A3(n5413), 
	.A2(net54895), 
	.A1(n976));
   AND2_X2 U5343 (.ZN(n1291), 
	.A2(n6025), 
	.A1(n6016));
   AND2_X2 U5344 (.ZN(n1937), 
	.A2(n6321), 
	.A1(n6312));
   NOR3_X1 U5346 (.ZN(n1214), 
	.A3(n2577), 
	.A2(n6349), 
	.A1(\UUT/Mpath/the_alu/N486 ));
   AND2_X1 U5347 (.ZN(\UUT/Mpath/the_alu/N118 ), 
	.A2(\UUT/Mpath/out_regB[7] ), 
	.A1(\UUT/Mpath/out_regA[7] ));
   OR2_X1 U5348 (.ZN(\UUT/Mpath/the_alu/N150 ), 
	.A2(\UUT/Mpath/out_regB[7] ), 
	.A1(\UUT/Mpath/out_regA[7] ));
   INV_X2 U5349 (.ZN(n1938), 
	.A(n5553));
   INV_X2 U5350 (.ZN(n1294), 
	.A(n5738));
   AND2_X1 U5351 (.ZN(\UUT/Mpath/the_alu/N111 ), 
	.A2(\UUT/Mpath/out_regB[14] ), 
	.A1(\UUT/Mpath/out_regA[14] ));
   OR2_X1 U5352 (.ZN(\UUT/Mpath/the_alu/N143 ), 
	.A2(\UUT/Mpath/out_regB[14] ), 
	.A1(\UUT/Mpath/out_regA[14] ));
   OR2_X1 U5353 (.ZN(\UUT/Mpath/the_alu/N144 ), 
	.A2(\UUT/Mpath/out_regB[13] ), 
	.A1(\UUT/Mpath/out_regA[13] ));
   AND2_X1 U5354 (.ZN(\UUT/Mpath/the_alu/N112 ), 
	.A2(\UUT/Mpath/out_regB[13] ), 
	.A1(\UUT/Mpath/out_regA[13] ));
   AND2_X1 U5355 (.ZN(\UUT/Mpath/the_alu/N114 ), 
	.A2(\UUT/Mpath/out_regB[11] ), 
	.A1(\UUT/Mpath/out_regA[11] ));
   OR2_X1 U5356 (.ZN(\UUT/Mpath/the_alu/N146 ), 
	.A2(\UUT/Mpath/out_regB[11] ), 
	.A1(\UUT/Mpath/out_regA[11] ));
   AND2_X2 U5357 (.ZN(n5540), 
	.A2(n6308), 
	.A1(n6305));
   AND2_X2 U5358 (.ZN(n5535), 
	.A2(n6302), 
	.A1(n6301));
   AND2_X2 U5359 (.ZN(n5725), 
	.A2(n6012), 
	.A1(n6009));
   AND2_X2 U5360 (.ZN(n5720), 
	.A2(n6006), 
	.A1(n6005));
   AND2_X2 U5361 (.ZN(n6199), 
	.A2(n6324), 
	.A1(\UUT/Mpath/the_shift/N108 ));
   AND3_X2 U5365 (.ZN(n5730), 
	.A3(n6016), 
	.A2(n6007), 
	.A1(\UUT/rs2_addr [4]));
   AND3_X2 U5366 (.ZN(n5557), 
	.A3(n6308), 
	.A2(n6310), 
	.A1(n6318));
   NAND3_X1 U5367 (.ZN(n6369), 
	.A3(n6308), 
	.A2(\UUT/rs1_addr [4]), 
	.A1(FE_OFCN199_UUT_rs1_addr_3_));
   INV_X1 U5368 (.ZN(n6370), 
	.A(n6369));
   INV_X1 U5369 (.ZN(n6371), 
	.A(n6369));
   AND3_X2 U5370 (.ZN(n5742), 
	.A3(n6012), 
	.A2(n6014), 
	.A1(n6022));
   AND3_X2 U5371 (.ZN(n1930), 
	.A3(n6310), 
	.A2(n2591), 
	.A1(n6308));
   AND2_X1 U5372 (.ZN(n6308), 
	.A2(n6303), 
	.A1(n6309));
   AND3_X2 U5373 (.ZN(n5735), 
	.A3(n6012), 
	.A2(\UUT/rs2_addr [4]), 
	.A1(\UUT/rs2_addr [3]));
   AND2_X1 U5374 (.ZN(\UUT/Mpath/the_alu/N113 ), 
	.A2(\UUT/Mpath/out_regB[12] ), 
	.A1(\UUT/Mpath/out_regA[12] ));
   OR2_X1 U5375 (.ZN(\UUT/Mpath/the_alu/N145 ), 
	.A2(\UUT/Mpath/out_regB[12] ), 
	.A1(\UUT/Mpath/out_regA[12] ));
   AND3_X2 U5376 (.ZN(n1282), 
	.A3(n6021), 
	.A2(n6008), 
	.A1(n6010));
   INV_X2 U5377 (.ZN(n1277), 
	.A(n5722));
   NAND2_X2 U5378 (.ZN(n5434), 
	.A2(\UUT/byp_controlB[0] ), 
	.A1(\UUT/byp_controlB[2] ));
   NAND3_X2 U5379 (.ZN(n133), 
	.A3(\UUT/Mpath/the_mult/N311 ), 
	.A2(n975), 
	.A1(\UUT/Mpath/the_mult/N285 ));
   INV_X2 U5380 (.ZN(n1926), 
	.A(n5537));
   NAND2_X2 U5381 (.ZN(n5558), 
	.A2(n6316), 
	.A1(n6319));
   AND3_X2 U5382 (.ZN(n291), 
	.A3(\UUT/Mpath/the_mult/N216 ), 
	.A2(n1194), 
	.A1(\UUT/Mpath/the_mult/N198 ));
   AND2_X1 U5383 (.ZN(\UUT/Mpath/the_alu/N96 ), 
	.A2(\UUT/Mpath/out_regB[29] ), 
	.A1(\UUT/Mpath/out_regA[29] ));
   OR2_X1 U5384 (.ZN(\UUT/Mpath/the_alu/N128 ), 
	.A2(\UUT/Mpath/out_regB[29] ), 
	.A1(\UUT/Mpath/out_regA[29] ));
   NAND2_X2 U5385 (.ZN(n5743), 
	.A2(n6020), 
	.A1(n6023));
   OR2_X1 U5386 (.ZN(\UUT/Mpath/the_alu/N152 ), 
	.A2(\UUT/Mpath/out_regB[5] ), 
	.A1(\UUT/Mpath/out_regA[5] ));
   AND2_X1 U5387 (.ZN(\UUT/Mpath/the_alu/N120 ), 
	.A2(\UUT/Mpath/out_regB[5] ), 
	.A1(\UUT/Mpath/out_regA[5] ));
   AND2_X1 U5388 (.ZN(\UUT/Mpath/the_alu/N99 ), 
	.A2(\UUT/Mpath/out_regB[26] ), 
	.A1(\UUT/Mpath/out_regA[26] ));
   OR2_X1 U5389 (.ZN(\UUT/Mpath/the_alu/N131 ), 
	.A2(\UUT/Mpath/out_regB[26] ), 
	.A1(\UUT/Mpath/out_regA[26] ));
   AND3_X2 U5390 (.ZN(n1931), 
	.A3(n6321), 
	.A2(n2591), 
	.A1(n6309));
   AND3_X2 U5391 (.ZN(n1284), 
	.A3(n6014), 
	.A2(\UUT/rs2_addr [3]), 
	.A1(n6012));
   NAND2_X2 U5392 (.ZN(n129), 
	.A2(\UUT/Mcontrol/st_logic/N42 ), 
	.A1(\UUT/byp_controlB[2] ));
   NAND2_X2 U5393 (.ZN(n5430), 
	.A2(\UUT/Mcontrol/st_logic/N42 ), 
	.A1(\UUT/byp_controlB[2] ));
   AND4_X2 U5394 (.ZN(n145), 
	.A4(n972), 
	.A3(n5413), 
	.A2(n971), 
	.A1(net54895));
   OR2_X2 U5395 (.ZN(n5432), 
	.A2(\UUT/regfile/N269 ), 
	.A1(\UUT/byp_controlB[2] ));
   INV_X2 U5397 (.ZN(n611), 
	.A(n620));
   INV_X2 U5398 (.ZN(n576), 
	.A(n585));
   INV_X2 U5399 (.ZN(n551), 
	.A(n560));
   INV_X2 U5400 (.ZN(n648), 
	.A(n657));
   INV_X2 U5401 (.ZN(n671), 
	.A(n680));
   INV_X2 U5402 (.ZN(n525), 
	.A(n534));
   INV_X2 U5403 (.ZN(n500), 
	.A(n509));
   INV_X2 U5404 (.ZN(n699), 
	.A(n708));
   INV_X2 U5405 (.ZN(n722), 
	.A(n731));
   INV_X2 U5406 (.ZN(n471), 
	.A(n480));
   INV_X2 U5407 (.ZN(n447), 
	.A(n459));
   INV_X2 U5408 (.ZN(n745), 
	.A(n754));
   INV_X2 U5409 (.ZN(n768), 
	.A(n777));
   INV_X2 U5410 (.ZN(n423), 
	.A(n432));
   INV_X2 U5411 (.ZN(n401), 
	.A(n410));
   INV_X2 U5412 (.ZN(n802), 
	.A(n800));
   INV_X2 U5413 (.ZN(n814), 
	.A(n812));
   INV_X2 U5414 (.ZN(n379), 
	.A(n388));
   INV_X2 U5415 (.ZN(n353), 
	.A(n362));
   INV_X2 U5416 (.ZN(n958), 
	.A(n641));
   INV_X2 U5417 (.ZN(n959), 
	.A(n605));
   INV_X2 U5418 (.ZN(n332), 
	.A(n341));
   INV_X2 U5419 (.ZN(n303), 
	.A(n315));
   INV_X2 U5420 (.ZN(n960), 
	.A(n1076));
   NAND2_X2 U5421 (.ZN(n5745), 
	.A2(n6018), 
	.A1(n6023));
   NAND2_X2 U5422 (.ZN(n5560), 
	.A2(n6314), 
	.A1(n6319));
   INV_X2 U5423 (.ZN(n1927), 
	.A(n5542));
   INV_X2 U5424 (.ZN(n1279), 
	.A(n5727));
   NAND3_X2 U5425 (.ZN(n5717), 
	.A3(n6005), 
	.A2(n6008), 
	.A1(n6007));
   NAND3_X2 U5426 (.ZN(n5532), 
	.A3(n6301), 
	.A2(n6304), 
	.A1(n6303));
   NAND3_X2 U5427 (.ZN(n5732), 
	.A3(n6006), 
	.A2(\UUT/rs2_addr [4]), 
	.A1(n6020));
   AND2_X1 U5428 (.ZN(\UUT/Mpath/the_alu/N101 ), 
	.A2(\UUT/Mpath/out_regB[24] ), 
	.A1(\UUT/Mpath/out_regA[24] ));
   OR2_X1 U5429 (.ZN(\UUT/Mpath/the_alu/N133 ), 
	.A2(\UUT/Mpath/out_regB[24] ), 
	.A1(\UUT/Mpath/out_regA[24] ));
   NAND3_X2 U5430 (.ZN(n5746), 
	.A3(n6025), 
	.A2(\UUT/rs2_addr [1]), 
	.A1(n6018));
   NAND3_X2 U5431 (.ZN(n5547), 
	.A3(n6302), 
	.A2(\UUT/rs1_addr [4]), 
	.A1(n6316));
   NOR2_X1 U5432 (.ZN(n6302), 
	.A2(\UUT/rs1_addr [0]), 
	.A1(n6304));
   NAND3_X2 U5433 (.ZN(n5561), 
	.A3(n6321), 
	.A2(FE_OFN98_UUT_rs1_addr_1_), 
	.A1(n6314));
   NAND3_X2 U5434 (.ZN(n5546), 
	.A3(FE_OFN98_UUT_rs1_addr_1_), 
	.A2(n6316), 
	.A1(n6313));
   NAND3_X2 U5435 (.ZN(n5731), 
	.A3(\UUT/rs2_addr [1]), 
	.A2(n6020), 
	.A1(n6017));
   NAND3_X2 U5437 (.ZN(n1934), 
	.A3(n6312), 
	.A2(n6310), 
	.A1(n6303));
   OR2_X1 U5438 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N114 ), 
	.A2(FE_OFN103_UUT_Mcontrol_Nextpc_decoding_N255), 
	.A1(\UUT/Mcontrol/st_logic/N103 ));
   OR2_X1 U5439 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N262 ), 
	.A2(FE_OFN103_UUT_Mcontrol_Nextpc_decoding_N255), 
	.A1(\UUT/Mcontrol/d_jump_type[3] ));
   AND2_X1 U5455 (.ZN(\UUT/Mpath/the_alu/N119 ), 
	.A2(\UUT/Mpath/out_regB[6] ), 
	.A1(\UUT/Mpath/out_regA[6] ));
   OR2_X1 U5456 (.ZN(\UUT/Mpath/the_alu/N151 ), 
	.A2(\UUT/Mpath/out_regB[6] ), 
	.A1(\UUT/Mpath/out_regA[6] ));
   NAND3_X2 U5457 (.ZN(n1287), 
	.A3(n6016), 
	.A2(n6014), 
	.A1(n6007));
   INV_X2 U5458 (.ZN(n1290), 
	.A(n5739));
   INV_X2 U5460 (.ZN(n1275), 
	.A(n5721));
   INV_X2 U5461 (.ZN(n1936), 
	.A(n5554));
   NAND2_X2 U5462 (.ZN(n131), 
	.A2(\UUT/byp_controlB[0] ), 
	.A1(\UUT/byp_controlB[2] ));
   INV_X2 U5463 (.ZN(n1925), 
	.A(n5536));
   NAND3_X2 U5464 (.ZN(n6373), 
	.A3(n6317), 
	.A2(n6304), 
	.A1(n6306));
   INV_X1 U5465 (.ZN(n6306), 
	.A(\UUT/rs1_addr [2]));
   NAND3_X2 U5466 (.ZN(n1288), 
	.A3(n6025), 
	.A2(\UUT/rs2_addr [3]), 
	.A1(n6013));
   NAND2_X1 U5467 (.ZN(n6374), 
	.A2(n6309), 
	.A1(n6317));
   INV_X1 U5468 (.ZN(n6375), 
	.A(n6374));
   INV_X1 U5469 (.ZN(n6376), 
	.A(n6374));
   AND2_X2 U5470 (.ZN(n5741), 
	.A2(n6013), 
	.A1(n6021));
   AND2_X2 U5471 (.ZN(n5544), 
	.A2(n6313), 
	.A1(n6312));
   AND2_X2 U5472 (.ZN(n144), 
	.A2(n973), 
	.A1(n975));
   NAND3_X2 U5473 (.ZN(n5737), 
	.A3(n6021), 
	.A2(n6010), 
	.A1(\UUT/rs2_addr [1]));
   AND2_X2 U5474 (.ZN(n5729), 
	.A2(n6017), 
	.A1(n6016));
   NAND3_X2 U5475 (.ZN(n5744), 
	.A3(n6025), 
	.A2(n6020), 
	.A1(\UUT/rs2_addr [1]));
   NAND3_X2 U5476 (.ZN(n5552), 
	.A3(n6317), 
	.A2(n6306), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   AND3_X2 U5477 (.ZN(n5549), 
	.A3(n6309), 
	.A2(FE_OFCN199_UUT_rs1_addr_3_), 
	.A1(n6313));
   NAND3_X2 U5478 (.ZN(n5559), 
	.A3(n6321), 
	.A2(n6316), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   AND3_X2 U5479 (.ZN(n5724), 
	.A3(n6009), 
	.A2(\UUT/rs2_addr [0]), 
	.A1(n6013));
   AND3_X2 U5480 (.ZN(n5719), 
	.A3(n6005), 
	.A2(\UUT/rs2_addr [0]), 
	.A1(\UUT/rs2_addr [1]));
   AND3_X2 U5481 (.ZN(n5734), 
	.A3(n6013), 
	.A2(\UUT/rs2_addr [3]), 
	.A1(n6017));
   AND3_X2 U5482 (.ZN(n5534), 
	.A3(n6301), 
	.A2(\UUT/rs1_addr [0]), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   NAND3_X2 U5483 (.ZN(n5716), 
	.A3(n6005), 
	.A2(n6008), 
	.A1(\UUT/rs2_addr [0]));
   AND3_X2 U5484 (.ZN(n5539), 
	.A3(n6305), 
	.A2(\UUT/rs1_addr [0]), 
	.A1(n6309));
   NAND3_X2 U5485 (.ZN(n140), 
	.A3(\UUT/Mpath/the_mult/N311 ), 
	.A2(n975), 
	.A1(\UUT/Mpath/the_mult/N255 ));
   NAND3_X2 U5486 (.ZN(n5531), 
	.A3(n6301), 
	.A2(n6304), 
	.A1(\UUT/rs1_addr [0]));
   NAND3_X2 U5487 (.ZN(n5736), 
	.A3(n6023), 
	.A2(n6022), 
	.A1(n6010));
   NAND3_X2 U5488 (.ZN(n5551), 
	.A3(n6319), 
	.A2(n6318), 
	.A1(n6306));
   NAND3_X2 U5489 (.ZN(n5541), 
	.A3(n6314), 
	.A2(n6313), 
	.A1(FE_OFN98_UUT_rs1_addr_1_));
   NAND3_X2 U5490 (.ZN(n5726), 
	.A3(n6018), 
	.A2(n6017), 
	.A1(\UUT/rs2_addr [1]));
   INV_X2 U5491 (.ZN(n181), 
	.A(n831));
   OAI221_X1 U5492 (.ZN(n831), 
	.C2(n5473), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5873), 
	.A(n282));
   INV_X2 U5493 (.ZN(n130), 
	.A(n849));
   OAI221_X1 U5494 (.ZN(n849), 
	.C2(n5464), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5851), 
	.A(n282));
   INV_X2 U5495 (.ZN(n194), 
	.A(n825));
   OAI221_X1 U5496 (.ZN(n825), 
	.C2(n5476), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5882), 
	.A(n282));
   INV_X2 U5497 (.ZN(n153), 
	.A(n843));
   OAI221_X1 U5498 (.ZN(n843), 
	.C2(n5467), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5857), 
	.A(n282));
   INV_X2 U5499 (.ZN(n952), 
	.A(n1171));
   OAI221_X1 U5500 (.ZN(n1171), 
	.C2(n5455), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5825), 
	.A(n282));
   INV_X2 U5501 (.ZN(n209), 
	.A(n280));
   OAI221_X1 U5502 (.ZN(n280), 
	.C2(n5479), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5890), 
	.A(n282));
   INV_X2 U5503 (.ZN(n165), 
	.A(n837));
   OAI221_X1 U5504 (.ZN(n837), 
	.C2(n5470), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5863), 
	.A(n282));
   INV_X2 U5505 (.ZN(n860), 
	.A(n869));
   OAI221_X1 U5506 (.ZN(n869), 
	.C2(n5458), 
	.C1(n5710), 
	.B2(n281), 
	.B1(n5832), 
	.A(n282));
   INV_X2 U5507 (.ZN(n82), 
	.A(n83));
   NOR2_X1 U5508 (.ZN(n319), 
	.A2(FE_OFN96_n5530), 
	.A1(FE_OFN11_net54953));
   NAND2_X2 U5509 (.ZN(n83), 
	.A2(net54859), 
	.A1(n116));
   NOR2_X1 U5510 (.ZN(n318), 
	.A2(FE_OFN97_n5529), 
	.A1(FE_OFN12_net54953));
   NOR2_X1 U5511 (.ZN(n314), 
	.A2(FE_OFN96_n5530), 
	.A1(FE_OFN8_n73));
   NOR2_X4 U5512 (.ZN(n5612), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n6284));
   NOR2_X1 U5513 (.ZN(n312), 
	.A2(FE_OFN97_n5529), 
	.A1(FE_OFN8_n73));
   NOR3_X1 U5514 (.ZN(n325), 
	.A3(n1195), 
	.A2(\UUT/Mpath/N114 ), 
	.A1(FE_OFN91_n285));
   NOR2_X4 U5517 (.ZN(n1208), 
	.A2(\UUT/Mpath/the_alu/N474 ), 
	.A1(n2573));
   NOR2_X4 U5518 (.ZN(n284), 
	.A2(\UUT/Mpath/the_mult/N216 ), 
	.A1(n1193));
   OR2_X1 U5519 (.ZN(\UUT/Mpath/the_mult/N216 ), 
	.A2(\UUT/Mpath/the_mult/N197 ), 
	.A1(\UUT/Mpath/the_mult/x_mul_command[0] ));
   NOR2_X4 U5520 (.ZN(n1210), 
	.A2(n2572), 
	.A1(FE_OFN87_n1211));
   NOR2_X4 U5521 (.ZN(n6198), 
	.A2(\UUT/Mpath/the_shift/N118 ), 
	.A1(n6325));
   NOR2_X4 U5522 (.ZN(n6200), 
	.A2(\UUT/Mpath/the_shift/N108 ), 
	.A1(n6323));
   NOR2_X4 U5523 (.ZN(n1212), 
	.A2(n6349), 
	.A1(n2576));
   NAND2_X2 U5524 (.ZN(n5528), 
	.A2(\UUT/Mcontrol/st_logic/N47 ), 
	.A1(\UUT/byp_controlA[2] ));
   NOR2_X4 U5525 (.ZN(n5779), 
	.A2(\localbus/c2_op[MASTER] ), 
	.A1(n6003));
   AND2_X1 U5527 (.ZN(\localbus/N93 ), 
	.A2(\localbus/N322 ), 
	.A1(\localbus/N335 ));
   NAND2_X1 U5528 (.ZN(n5530), 
	.A2(\UUT/byp_controlA[0] ), 
	.A1(\UUT/byp_controlA[2] ));
   INV_X2 U5531 (.ZN(n6380), 
	.A(n249));
   INV_X2 U5532 (.ZN(n249), 
	.A(n248));
   NOR2_X1 U5533 (.ZN(n285), 
	.A2(\UUT/Mpath/N117 ), 
	.A1(\UUT/exe_outsel [0]));
   INV_X2 U5535 (.ZN(n6381), 
	.A(n253));
   INV_X2 U5536 (.ZN(n6382), 
	.A(n247));
   INV_X2 U5537 (.ZN(n6383), 
	.A(n245));
   INV_X2 U5538 (.ZN(n6384), 
	.A(n251));
   INV_X2 U5539 (.ZN(n253), 
	.A(n252));
   INV_X2 U5540 (.ZN(n247), 
	.A(n246));
   INV_X2 U5541 (.ZN(n245), 
	.A(n244));
   INV_X2 U5542 (.ZN(n251), 
	.A(n250));
   INV_X2 U5543 (.ZN(n6385), 
	.A(n243));
   INV_X2 U5544 (.ZN(n6386), 
	.A(n257));
   INV_X2 U5545 (.ZN(n6387), 
	.A(n255));
   INV_X2 U5546 (.ZN(n6388), 
	.A(n241));
   INV_X2 U5547 (.ZN(n243), 
	.A(n242));
   INV_X2 U5548 (.ZN(n257), 
	.A(n256));
   INV_X2 U5549 (.ZN(n255), 
	.A(n254));
   INV_X2 U5550 (.ZN(n241), 
	.A(n240));
   INV_X2 U5551 (.ZN(n6389), 
	.A(n263));
   INV_X2 U5552 (.ZN(n6390), 
	.A(n239));
   INV_X2 U5553 (.ZN(n6391), 
	.A(n237));
   INV_X2 U5554 (.ZN(n6392), 
	.A(n259));
   INV_X2 U5555 (.ZN(n263), 
	.A(n262));
   INV_X2 U5556 (.ZN(n239), 
	.A(n238));
   INV_X2 U5557 (.ZN(n237), 
	.A(n236));
   INV_X2 U5558 (.ZN(n259), 
	.A(n258));
   INV_X2 U5559 (.ZN(n6393), 
	.A(n235));
   INV_X2 U5560 (.ZN(n6394), 
	.A(n261));
   INV_X2 U5561 (.ZN(n6395), 
	.A(n265));
   INV_X2 U5562 (.ZN(n6396), 
	.A(n233));
   INV_X2 U5563 (.ZN(n235), 
	.A(n234));
   INV_X2 U5564 (.ZN(n261), 
	.A(n260));
   INV_X2 U5565 (.ZN(n265), 
	.A(n264));
   INV_X2 U5566 (.ZN(n233), 
	.A(n232));
   INV_X2 U5567 (.ZN(n6397), 
	.A(n271));
   INV_X2 U5568 (.ZN(n6398), 
	.A(n231));
   INV_X2 U5569 (.ZN(n6399), 
	.A(n227));
   INV_X2 U5570 (.ZN(n6400), 
	.A(n267));
   INV_X2 U5571 (.ZN(n271), 
	.A(n270));
   INV_X2 U5572 (.ZN(n231), 
	.A(n230));
   INV_X2 U5573 (.ZN(n227), 
	.A(n226));
   INV_X2 U5574 (.ZN(n267), 
	.A(n266));
   INV_X2 U5575 (.ZN(n6401), 
	.A(n223));
   INV_X2 U5576 (.ZN(n6402), 
	.A(n269));
   INV_X2 U5577 (.ZN(n6403), 
	.A(n273));
   INV_X2 U5578 (.ZN(n6404), 
	.A(n229));
   INV_X2 U5579 (.ZN(n223), 
	.A(n222));
   INV_X2 U5580 (.ZN(n269), 
	.A(n268));
   INV_X2 U5581 (.ZN(n273), 
	.A(n272));
   INV_X2 U5582 (.ZN(n229), 
	.A(n228));
   INV_X2 U5583 (.ZN(n6405), 
	.A(n277));
   INV_X2 U5584 (.ZN(n6406), 
	.A(n225));
   INV_X2 U5585 (.ZN(n6407), 
	.A(n219));
   INV_X2 U5586 (.ZN(n6408), 
	.A(n275));
   INV_X2 U5587 (.ZN(n277), 
	.A(n276));
   INV_X2 U5588 (.ZN(n225), 
	.A(n224));
   INV_X2 U5589 (.ZN(n219), 
	.A(n218));
   INV_X2 U5590 (.ZN(n275), 
	.A(n274));
   INV_X2 U5592 (.ZN(n6410), 
	.A(n221));
   INV_X2 U5593 (.ZN(n6411), 
	.A(n279));
   INV_X2 U5594 (.ZN(n147), 
	.A(FE_OFN8_n73));
   NOR2_X4 U5595 (.ZN(n5564), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(\UUT/Mpath/N115 ));
   INV_X2 U5596 (.ZN(n221), 
	.A(n220));
   INV_X2 U5597 (.ZN(n279), 
	.A(n278));
   INV_X1 U5598 (.ZN(n6650), 
	.A(\UUT/jar_in [7]));
   INV_X1 U5599 (.ZN(n6648), 
	.A(\UUT/jar_in [3]));
   INV_X1 U5600 (.ZN(n6655), 
	.A(\UUT/jar_in [6]));
   NAND2_X1 U5601 (.ZN(n6412), 
	.A2(n6467), 
	.A1(n6466));
   NAND2_X1 U5602 (.ZN(n2895), 
	.A2(n6413), 
	.A1(n136));
   INV_X1 U5603 (.ZN(n6413), 
	.A(n6412));
   AOI21_X1 U5604 (.ZN(n136), 
	.B2(\UUT/Mpath/the_mult/Mad_out [61]), 
	.B1(n139), 
	.A(n6428));
   OR2_X1 U5605 (.ZN(n6466), 
	.A2(n134), 
	.A1(n133));
   OR2_X1 U5606 (.ZN(n6414), 
	.A2(n154), 
	.A1(n133));
   OR2_X1 U5607 (.ZN(n6415), 
	.A2(n135), 
	.A1(n5689));
   NAND3_X1 U5608 (.ZN(n2901), 
	.A3(n155), 
	.A2(n6415), 
	.A1(n6414));
   AND2_X1 U5609 (.ZN(n155), 
	.A2(n6458), 
	.A1(n6457));
   OR2_X1 U5610 (.ZN(n6416), 
	.A2(n466), 
	.A1(n294));
   OR2_X1 U5611 (.ZN(n6417), 
	.A2(n2660), 
	.A1(n295));
   NAND3_X1 U5612 (.ZN(n3243), 
	.A3(n468), 
	.A2(n6417), 
	.A1(n6416));
   AND3_X1 U5613 (.ZN(n468), 
	.A3(n6618), 
	.A2(n6617), 
	.A1(n6616));
   AOI22_X1 U5614 (.ZN(n2327), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/Bta [2]), 
	.B1(n6449), 
	.A2(\UUT/break_code[2] ), 
	.A1(n908));
   OR2_X1 U5615 (.ZN(n6633), 
	.A2(n6488), 
	.A1(n6634));
   OR2_X1 U5616 (.ZN(n6418), 
	.A2(n294), 
	.A1(n787));
   OR2_X1 U5617 (.ZN(n6419), 
	.A2(n2698), 
	.A1(n295));
   NAND3_X1 U5618 (.ZN(n3735), 
	.A3(n790), 
	.A2(n6419), 
	.A1(n6418));
   AND3_X1 U5619 (.ZN(n790), 
	.A3(n6538), 
	.A2(n6537), 
	.A1(n6536));
   AND3_X1 U5620 (.ZN(n571), 
	.A3(n2374), 
	.A2(n6704), 
	.A1(n6703));
   OR2_X1 U5621 (.ZN(n6420), 
	.A2(n6687), 
	.A1(n6531));
   OR2_X1 U5622 (.ZN(n6421), 
	.A2(n6688), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N125 ));
   NAND3_X1 U5623 (.ZN(n6686), 
	.A3(n2351), 
	.A2(n6421), 
	.A1(n6420));
   INV_X1 U5624 (.ZN(n6687), 
	.A(\UUT/jar_in [12]));
   INV_X1 U5625 (.ZN(n6688), 
	.A(\UUT/branch_rega [12]));
   NAND2_X1 U5626 (.ZN(n6422), 
	.A2(n6907), 
	.A1(n6906));
   NAND3_X1 U5627 (.ZN(n6909), 
	.A3(n6905), 
	.A2(n6423), 
	.A1(n6908));
   INV_X1 U5628 (.ZN(n6423), 
	.A(n6422));
   NAND2_X1 U5629 (.ZN(n6424), 
	.A2(\localbus/c1_addr_outbus[29] ), 
	.A1(\localbus/c1_addr_outbus[30] ));
   INV_X1 U5630 (.ZN(n6425), 
	.A(n6595));
   AND2_X1 U5631 (.ZN(n6903), 
	.A2(n6425), 
	.A1(n6424));
   AND2_X1 U5632 (.ZN(n6595), 
	.A2(n6644), 
	.A1(n6347));
   NOR2_X1 U5633 (.ZN(n5456), 
	.A2(n6481), 
	.A1(n6480));
   AND2_X1 U5634 (.ZN(n6481), 
	.A2(n5564), 
	.A1(n5563));
   NAND4_X1 U5636 (.ZN(n6128), 
	.A4(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A3(n6045), 
	.A2(n6285), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N89 ));
   AND4_X1 U5637 (.ZN(n6915), 
	.A4(n4358), 
	.A3(n4357), 
	.A2(n4359), 
	.A1(n6447));
   NOR4_X1 U5638 (.ZN(n6447), 
	.A4(\localbus/c1_addr_outbus[29] ), 
	.A3(n6595), 
	.A2(\localbus/c1_addr_outbus[27] ), 
	.A1(\localbus/c1_addr_outbus[28] ));
   NOR2_X1 U5640 (.ZN(n6449), 
	.A2(n6615), 
	.A1(n6693));
   NAND2_X1 U5643 (.ZN(n6451), 
	.A2(n6469), 
	.A1(n6468));
   OR2_X1 U5647 (.ZN(n6454), 
	.A2(n294), 
	.A1(n395));
   OR2_X1 U5648 (.ZN(n6455), 
	.A2(n2651), 
	.A1(n295));
   NAND3_X1 U5649 (.ZN(n3123), 
	.A3(n398), 
	.A2(n6455), 
	.A1(n6454));
   AND2_X1 U5651 (.ZN(n297), 
	.A2(n295), 
	.A1(n2324));
   AND2_X1 U5653 (.ZN(n6711), 
	.A2(n295), 
	.A1(n2324));
   OR2_X1 U5655 (.ZN(n6469), 
	.A2(n6456), 
	.A1(n6693));
   NAND2_X1 U5656 (.ZN(n6456), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/Bta [9]), 
	.A1(n6614));
   NAND2_X1 U5657 (.ZN(n6457), 
	.A2(n156), 
	.A1(n137));
   NAND2_X1 U5658 (.ZN(n6458), 
	.A2(n139), 
	.A1(\UUT/Mpath/the_mult/Mad_out [60]));
   NAND2_X1 U5659 (.ZN(n6459), 
	.A2(n6583), 
	.A1(n6582));
   NAND2_X1 U5660 (.ZN(n4041), 
	.A2(n6460), 
	.A1(n905));
   INV_X1 U5661 (.ZN(n6460), 
	.A(n6459));
   NAND2_X1 U5662 (.ZN(n6461), 
	.A2(n139), 
	.A1(\UUT/Mpath/the_mult/Mad_out [63]));
   NAND2_X1 U5663 (.ZN(n4329), 
	.A2(net56414), 
	.A1(n6461));
   OAI22_X2 U5664 (.ZN(n6641), 
	.B2(\UUT/Mcontrol/st_logic/N89 ), 
	.B1(n6293), 
	.A2(n6292), 
	.A1(n6633));
   NAND2_X1 U5665 (.ZN(n6462), 
	.A2(n6573), 
	.A1(n6572));
   AND3_X1 U5666 (.ZN(n6463), 
	.A3(n2536), 
	.A2(n6513), 
	.A1(n6512));
   OR2_X1 U5667 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N27 ), 
	.A2(n6488), 
	.A1(n6831));
   AND2_X1 U5668 (.ZN(n299), 
	.A2(n295), 
	.A1(n6714));
   AND2_X1 U5669 (.ZN(n6511), 
	.A2(n295), 
	.A1(n6714));
   AOI22_X1 U5671 (.ZN(n5462), 
	.B2(n5564), 
	.B1(n5571), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5570));
   OR2_X1 U5672 (.ZN(n6573), 
	.A2(n6465), 
	.A1(n6693));
   NAND2_X1 U5673 (.ZN(n6465), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/Bta [10]), 
	.A1(n6614));
   OR3_X1 U5674 (.ZN(n6637), 
	.A3(n4339), 
	.A2(n4340), 
	.A1(\localbus/N57 ));
   OR2_X1 U5675 (.ZN(n6467), 
	.A2(n135), 
	.A1(n5688));
   OAI22_X1 U5676 (.ZN(n6289), 
	.B2(\UUT/Mcontrol/st_logic/N89 ), 
	.B1(n6293), 
	.A2(n6292), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N27 ));
   OAI222_X1 U5677 (.ZN(n6488), 
	.C2(FE_OFN96_n5530), 
	.C1(n5455), 
	.B2(FE_OFN97_n5529), 
	.B1(n5414), 
	.A2(n5528), 
	.A1(n6619));
   AND2_X1 U5678 (.ZN(n6872), 
	.A2(n6519), 
	.A1(n6845));
   NOR3_X1 U5679 (.ZN(n979), 
	.A3(n6462), 
	.A2(n6677), 
	.A1(n6676));
   NAND2_X1 U5680 (.ZN(net87679), 
	.A2(n138), 
	.A1(n137));
   NAND2_X1 U5681 (.ZN(n6468), 
	.A2(\UUT/break_code[9] ), 
	.A1(n908));
   OAI222_X1 U5682 (.ZN(\UUT/branch_regb [31]), 
	.C2(n5434), 
	.C1(n5455), 
	.B2(n5432), 
	.B1(n5454), 
	.A2(n6619), 
	.A1(n5430));
   NAND2_X1 U5683 (.ZN(n6470), 
	.A2(n1259), 
	.A1(n1260));
   NAND2_X1 U5684 (.ZN(n5563), 
	.A2(n6471), 
	.A1(n1261));
   INV_X1 U5685 (.ZN(n6471), 
	.A(n6470));
   AOI21_X1 U5686 (.ZN(n6472), 
	.B2(\UUT/Mcontrol/st_logic/N70 ), 
	.B1(n6641), 
	.A(n6291));
   NAND2_X1 U5688 (.ZN(n6473), 
	.A2(n139), 
	.A1(\UUT/Mpath/the_mult/Mad_out [62]));
   NAND2_X1 U5689 (.ZN(n3977), 
	.A2(n6474), 
	.A1(n6473));
   AND2_X1 U5690 (.ZN(n6474), 
	.A2(n6694), 
	.A1(n6483));
   NAND2_X1 U5691 (.ZN(n6476), 
	.A2(\UUT/jar_in [20]), 
	.A1(n6711));
   NAND2_X1 U5692 (.ZN(n6477), 
	.A2(\UUT/branch_rega [20]), 
	.A1(n298));
   NAND2_X1 U5693 (.ZN(n6478), 
	.A2(n299), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [20]));
   AND3_X1 U5694 (.ZN(n350), 
	.A3(n6478), 
	.A2(n6477), 
	.A1(n6476));
   OAI22_X1 U5695 (.ZN(n6479), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), 
	.B1(n6472), 
	.A2(n6287), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N22 ));
   AND2_X1 U5696 (.ZN(n6480), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5562));
   NAND2_X1 U5698 (.ZN(n6482), 
	.A2(n6844), 
	.A1(n6843));
   INV_X1 U5699 (.ZN(n6483), 
	.A(n6482));
   AOI22_X1 U5700 (.ZN(n6619), 
	.B2(n5564), 
	.B1(n6690), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n6197));
   OR2_X1 U5701 (.ZN(n6769), 
	.A2(n6776), 
	.A1(\UUT/branch_rega [16]));
   AOI222_X2 U5702 (.ZN(n5486), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[21] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n346), 
	.A2(n5564), 
	.A1(n6107));
   AND2_X1 U5703 (.ZN(n6581), 
	.A2(n6736), 
	.A1(n6484));
   INV_X1 U5704 (.ZN(n6484), 
	.A(n6621));
   NAND2_X1 U5705 (.ZN(n5571), 
	.A2(n6561), 
	.A1(n1255));
   NAND3_X1 U5708 (.ZN(n6487), 
	.A3(n2374), 
	.A2(n6704), 
	.A1(n6703));
   OAI222_X1 U5709 (.ZN(n6489), 
	.C2(FE_OFN96_n5530), 
	.C1(n5455), 
	.B2(FE_OFN97_n5529), 
	.B1(n5414), 
	.A2(n5528), 
	.A1(n6619));
   OAI222_X1 U5710 (.ZN(\UUT/branch_rega [31]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5455), 
	.B2(FE_OFN97_n5529), 
	.B1(n5414), 
	.A2(n5528), 
	.A1(n6619));
   OR2_X1 U5712 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1945 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1938 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   INV_X1 U5713 (.ZN(n643), 
	.A(n6649));
   OAI221_X1 U5714 (.ZN(n6649), 
	.C2(n6733), 
	.C1(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.B2(n6650), 
	.B1(n6531), 
	.A(n2466));
   NAND2_X1 U5715 (.ZN(n6490), 
	.A2(n297), 
	.A1(\UUT/jar_in [17]));
   NAND2_X1 U5716 (.ZN(n6491), 
	.A2(\UUT/branch_rega [17]), 
	.A1(n298));
   NAND2_X1 U5717 (.ZN(n6492), 
	.A2(n299), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [17]));
   AND3_X1 U5718 (.ZN(n420), 
	.A3(n6492), 
	.A2(n6491), 
	.A1(n6490));
   OAI222_X1 U5719 (.ZN(\UUT/branch_rega [17]), 
	.C2(n5501), 
	.C1(n5528), 
	.B2(n2223), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5503));
   NAND2_X1 U5720 (.ZN(n6493), 
	.A2(\UUT/break_code[4] ), 
	.A1(n908));
   NAND2_X1 U5721 (.ZN(n6494), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/Bta [4]), 
	.A1(n6449));
   AND2_X1 U5722 (.ZN(n2536), 
	.A2(n6494), 
	.A1(n6493));
   AND3_X1 U5723 (.ZN(n6640), 
	.A3(n6544), 
	.A2(n6545), 
	.A1(n6530));
   AOI22_X1 U5724 (.ZN(n764), 
	.B2(\UUT/Mcontrol/d_sampled_finstr [2]), 
	.B1(n2329), 
	.A2(n2328), 
	.A1(n6263));
   NAND2_X1 U5725 (.ZN(n6495), 
	.A2(n6631), 
	.A1(n6630));
   NAND2_X1 U5726 (.ZN(n2963), 
	.A2(n6496), 
	.A1(n296));
   INV_X1 U5727 (.ZN(n6496), 
	.A(n6495));
   NAND2_X1 U5728 (.ZN(n6497), 
	.A2(n297), 
	.A1(\UUT/jar_in [22]));
   NAND2_X1 U5729 (.ZN(n6498), 
	.A2(\UUT/branch_rega [22]), 
	.A1(n298));
   NAND2_X1 U5730 (.ZN(n6499), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/Bta [22]), 
	.A1(n6511));
   AND3_X1 U5731 (.ZN(n296), 
	.A3(n6499), 
	.A2(n6498), 
	.A1(n6497));
   OAI22_X1 U5732 (.ZN(n6294), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/N242 ), 
	.B1(n6298), 
	.A2(n6489), 
	.A1(n6297));
   AND2_X1 U5734 (.ZN(\UUT/Mpath/the_alu/N121 ), 
	.A2(\UUT/Mpath/out_regB[4] ), 
	.A1(\UUT/Mpath/out_regA[4] ));
   OR2_X1 U5735 (.ZN(\UUT/Mpath/the_alu/N153 ), 
	.A2(FE_OFN159_UUT_Mpath_out_regB_4_), 
	.A1(\UUT/Mpath/out_regA[4] ));
   NAND2_X1 U5736 (.ZN(n6500), 
	.A2(n297), 
	.A1(\UUT/jar_in [16]));
   NAND2_X1 U5737 (.ZN(n6501), 
	.A2(\UUT/branch_rega [16]), 
	.A1(n298));
   NAND2_X1 U5738 (.ZN(n6502), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/Bta [16]), 
	.A1(n299));
   AND3_X1 U5739 (.ZN(n442), 
	.A3(n6502), 
	.A2(n6501), 
	.A1(n6500));
   OAI222_X1 U5740 (.ZN(\UUT/branch_rega [16]), 
	.C2(n5504), 
	.C1(n5528), 
	.B2(n2243), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5506));
   NOR2_X1 U5741 (.ZN(n6862), 
	.A2(n6504), 
	.A1(n6725));
   NAND2_X1 U5742 (.ZN(n6504), 
	.A2(n6876), 
	.A1(n6505));
   AND2_X1 U5743 (.ZN(n6505), 
	.A2(n6712), 
	.A1(n6868));
   OR2_X1 U5744 (.ZN(n6506), 
	.A2(n6849), 
	.A1(n6531));
   OR2_X1 U5745 (.ZN(n6507), 
	.A2(n6854), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N125 ));
   NAND3_X1 U5746 (.ZN(n6848), 
	.A3(n2512), 
	.A2(n6507), 
	.A1(n6506));
   INV_X1 U5747 (.ZN(n6849), 
	.A(\UUT/jar_in [5]));
   OAI21_X1 U5749 (.ZN(n907), 
	.B2(n2560), 
	.B1(n6479), 
	.A(n2561));
   INV_X1 U5750 (.ZN(n666), 
	.A(n6654));
   NOR2_X1 U5751 (.ZN(n6714), 
	.A2(n6693), 
	.A1(n6615));
   NAND2_X1 U5752 (.ZN(n6508), 
	.A2(n6597), 
	.A1(n6596));
   NAND2_X1 U5753 (.ZN(n3043), 
	.A2(n6509), 
	.A1(n350));
   INV_X1 U5754 (.ZN(n6509), 
	.A(n6508));
   AND2_X1 U5755 (.ZN(n6510), 
	.A2(n295), 
	.A1(n6714));
   OR2_X1 U5756 (.ZN(n6512), 
	.A2(n6856), 
	.A1(n6531));
   OR2_X1 U5757 (.ZN(n6513), 
	.A2(n6868), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N125 ));
   NAND3_X1 U5758 (.ZN(n6855), 
	.A3(n2536), 
	.A2(n6513), 
	.A1(n6512));
   INV_X1 U5759 (.ZN(n6856), 
	.A(\UUT/jar_in [4]));
   NAND2_X1 U5761 (.ZN(n6514), 
	.A2(n6624), 
	.A1(n6623));
   NAND2_X1 U5762 (.ZN(n3163), 
	.A2(n6515), 
	.A1(n420));
   INV_X1 U5763 (.ZN(n6515), 
	.A(n6514));
   OR2_X1 U5764 (.ZN(n6690), 
	.A2(n6576), 
	.A1(n6516));
   NAND2_X1 U5765 (.ZN(n6516), 
	.A2(n6696), 
	.A1(n6530));
   NOR2_X1 U5768 (.ZN(n1261), 
	.A2(n6666), 
	.A1(n6522));
   NAND2_X1 U5769 (.ZN(n6522), 
	.A2(n6524), 
	.A1(n6523));
   NOR2_X1 U5770 (.ZN(n6519), 
	.A2(n6745), 
	.A1(\UUT/branch_rega [26]));
   NAND2_X1 U5771 (.ZN(n6520), 
	.A2(n1247), 
	.A1(n1248));
   NAND2_X1 U5772 (.ZN(n5578), 
	.A2(n6521), 
	.A1(n1249));
   INV_X1 U5773 (.ZN(n6521), 
	.A(n6520));
   NAND2_X1 U5774 (.ZN(n6523), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[30] ));
   NAND2_X1 U5775 (.ZN(n6524), 
	.A2(n1262), 
	.A1(n1208));
   AND2_X1 U5776 (.ZN(n6676), 
	.A2(\UUT/jar_in [10]), 
	.A1(n2324));
   AND2_X1 U5777 (.ZN(n6672), 
	.A2(\UUT/jar_in [9]), 
	.A1(n2324));
   NAND2_X1 U5779 (.ZN(n6526), 
	.A2(\UUT/break_code[5] ), 
	.A1(n908));
   NAND2_X1 U5780 (.ZN(n6527), 
	.A2(n6449), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [5]));
   AND2_X1 U5781 (.ZN(n2512), 
	.A2(n6526), 
	.A1(n6527));
   INV_X1 U5782 (.ZN(n740), 
	.A(n6647));
   NAND2_X1 U5783 (.ZN(n6528), 
	.A2(\UUT/Mcontrol/d_instr [6]), 
	.A1(n935));
   NAND2_X1 U5784 (.ZN(n2076), 
	.A2(n6529), 
	.A1(n6086));
   INV_X1 U5785 (.ZN(n6529), 
	.A(n6528));
   NAND2_X1 U5786 (.ZN(n6057), 
	.A2(n6067), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1945 ));
   INV_X1 U5787 (.ZN(n6079), 
	.A(n6046));
   NOR2_X1 U5788 (.ZN(n6045), 
	.A2(n6057), 
	.A1(n6079));
   NAND2_X1 U5789 (.ZN(n6530), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[31] ));
   OAI22_X1 U5790 (.ZN(n6693), 
	.B2(\UUT/Mcontrol/Nextpc_decoding/N266 ), 
	.B1(n6288), 
	.A2(n6287), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N22 ));
   OAI21_X1 U5791 (.ZN(n6531), 
	.B2(n2560), 
	.B1(n6479), 
	.A(n2561));
   NAND3_X1 U5792 (.ZN(n6053), 
	.A3(n6210), 
	.A2(n6040), 
	.A1(n6328));
   OR2_X1 U5793 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1889 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1875 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1876 ));
   OR2_X1 U5796 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1923 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1875 ), 
	.A1(\UUT/Mcontrol/d_instr [30]));
   INV_X1 U5805 (.ZN(n545), 
	.A(n6686));
   NOR2_X1 U5806 (.ZN(n6819), 
	.A2(n6532), 
	.A1(n6575));
   NAND2_X1 U5807 (.ZN(n6532), 
	.A2(n6851), 
	.A1(n6533));
   AND2_X1 U5808 (.ZN(n6533), 
	.A2(n6775), 
	.A1(n6549));
   NAND2_X1 U5809 (.ZN(n6534), 
	.A2(n1241), 
	.A1(n1242));
   NAND2_X1 U5810 (.ZN(n5585), 
	.A2(n6535), 
	.A1(n1243));
   INV_X1 U5811 (.ZN(n6535), 
	.A(n6534));
   NAND2_X1 U5812 (.ZN(n6536), 
	.A2(n6711), 
	.A1(\UUT/jar_in [1]));
   NAND2_X1 U5813 (.ZN(n6537), 
	.A2(FE_OFN187_UUT_branch_rega_1_), 
	.A1(n298));
   NAND2_X1 U5814 (.ZN(n6538), 
	.A2(n299), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [1]));
   OR2_X1 U5819 (.ZN(\UUT/Mpath/the_alu/N154 ), 
	.A2(\UUT/Mpath/out_regB[3] ), 
	.A1(\UUT/Mpath/out_regA[3] ));
   AND2_X1 U5820 (.ZN(\UUT/Mpath/the_alu/N122 ), 
	.A2(\UUT/Mpath/out_regB[3] ), 
	.A1(\UUT/Mpath/out_regA[3] ));
   OR2_X1 U5821 (.ZN(n6543), 
	.A2(n6910), 
	.A1(\localbus/c1_addr_outbus[30] ));
   NAND2_X1 U5822 (.ZN(\localbus/N56 ), 
	.A2(n6909), 
	.A1(n6543));
   NAND2_X1 U5823 (.ZN(n6544), 
	.A2(n1209), 
	.A1(n1208));
   NAND2_X1 U5824 (.ZN(n6545), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[31] ));
   OR2_X1 U5825 (.ZN(n6875), 
	.A2(\UUT/branch_rega [29]), 
	.A1(\UUT/branch_rega [28]));
   AND3_X1 U5826 (.ZN(n1255), 
	.A3(n6548), 
	.A2(n6547), 
	.A1(n6546));
   INV_X1 U5827 (.ZN(n6546), 
	.A(n6629));
   NAND2_X1 U5828 (.ZN(n6547), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[29] ));
   NAND2_X1 U5829 (.ZN(n6548), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[29] ));
   OR2_X1 U5830 (.ZN(n6608), 
	.A2(n5528), 
	.A1(n5462));
   AND2_X1 U5831 (.ZN(n6720), 
	.A2(n6723), 
	.A1(n6825));
   NOR2_X1 U5834 (.ZN(n6736), 
	.A2(\UUT/branch_rega [29]), 
	.A1(\UUT/branch_rega [28]));
   AND2_X1 U5835 (.ZN(n6549), 
	.A2(n6834), 
	.A1(n6833));
   NOR2_X1 U5836 (.ZN(n6838), 
	.A2(n6550), 
	.A1(n6850));
   NAND2_X1 U5837 (.ZN(n6550), 
	.A2(n6885), 
	.A1(n6697));
   NAND2_X1 U5838 (.ZN(n6551), 
	.A2(n1235), 
	.A1(n1236));
   NAND2_X1 U5839 (.ZN(n5592), 
	.A2(n6552), 
	.A1(n1237));
   INV_X1 U5840 (.ZN(n6552), 
	.A(n6551));
   NAND2_X1 U5841 (.ZN(n6553), 
	.A2(n6556), 
	.A1(n1237));
   NAND2_X1 U5842 (.ZN(n5471), 
	.A2(n6554), 
	.A1(n6553));
   OR2_X1 U5843 (.ZN(n6554), 
	.A2(n5564), 
	.A1(n6555));
   INV_X1 U5844 (.ZN(n6555), 
	.A(n6578));
   AND2_X1 U5845 (.ZN(n6556), 
	.A2(n6578), 
	.A1(n6552));
   OAI222_X1 U5846 (.ZN(\UUT/branch_rega [28]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5467), 
	.B2(FE_OFN97_n5529), 
	.B1(n5417), 
	.A2(n5528), 
	.A1(n5465));
   AOI222_X2 U5847 (.ZN(n1249), 
	.C2(FE_OFN87_n1211), 
	.C1(\UUT/Mpath/the_alu/sum[28] ), 
	.B2(n1210), 
	.B1(\UUT/Mpath/the_alu/diff[28] ), 
	.A2(n1250), 
	.A1(n1208));
   AOI22_X2 U5848 (.ZN(n5465), 
	.B2(n5564), 
	.B1(n5578), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5577));
   NAND2_X1 U5850 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N222 ), 
	.A2(n6559), 
	.A1(n6558));
   AND2_X2 U5851 (.ZN(n6558), 
	.A2(n6813), 
	.A1(n6829));
   NOR2_X1 U5852 (.ZN(n6559), 
	.A2(n6721), 
	.A1(n6671));
   NAND2_X1 U5853 (.ZN(n6560), 
	.A2(n1253), 
	.A1(n1254));
   INV_X1 U5854 (.ZN(n6561), 
	.A(n6560));
   NAND2_X1 U5855 (.ZN(n6562), 
	.A2(n6711), 
	.A1(\UUT/jar_in [18]));
   NAND2_X1 U5856 (.ZN(n6563), 
	.A2(\UUT/branch_rega [18]), 
	.A1(n298));
   NAND2_X1 U5857 (.ZN(n6564), 
	.A2(n6511), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [18]));
   AND3_X1 U5858 (.ZN(n398), 
	.A3(n6564), 
	.A2(n6563), 
	.A1(n6562));
   OAI222_X1 U5859 (.ZN(\UUT/branch_regb [29]), 
	.C2(n5434), 
	.C1(n5464), 
	.B2(n5432), 
	.B1(n5463), 
	.A2(n5430), 
	.A1(n5462));
   NAND2_X1 U5860 (.ZN(n6565), 
	.A2(n6610), 
	.A1(n6609));
   NAND2_X1 U5861 (.ZN(\UUT/branch_rega [29]), 
	.A2(n6566), 
	.A1(n6608));
   INV_X1 U5862 (.ZN(n6566), 
	.A(n6565));
   OR2_X1 U5863 (.ZN(n6567), 
	.A2(n294), 
	.A1(n369));
   OR2_X1 U5864 (.ZN(n6568), 
	.A2(n2648), 
	.A1(n295));
   NAND3_X1 U5865 (.ZN(n3083), 
	.A3(n372), 
	.A2(n6568), 
	.A1(n6567));
   NAND2_X1 U5866 (.ZN(n6569), 
	.A2(n6711), 
	.A1(\UUT/jar_in [19]));
   NAND2_X1 U5867 (.ZN(n6570), 
	.A2(\UUT/branch_rega [19]), 
	.A1(n298));
   NAND2_X1 U5868 (.ZN(n6571), 
	.A2(n6511), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [19]));
   AND3_X1 U5869 (.ZN(n372), 
	.A3(n6571), 
	.A2(n6570), 
	.A1(n6569));
   OR2_X1 U5870 (.ZN(n6610), 
	.A2(FE_OFN96_n5530), 
	.A1(n5464));
   NAND2_X1 U5871 (.ZN(n6572), 
	.A2(\UUT/break_code[10] ), 
	.A1(n908));
   OR2_X1 U5872 (.ZN(n6663), 
	.A2(n5528), 
	.A1(n5456));
   AND2_X1 U5873 (.ZN(\UUT/Mpath/the_alu/N123 ), 
	.A2(FE_OFN168_UUT_Mpath_out_regB_2_), 
	.A1(FE_OFCN198_UUT_Mpath_out_regA_2_));
   OR2_X1 U5874 (.ZN(\UUT/Mpath/the_alu/N155 ), 
	.A2(FE_OFN168_UUT_Mpath_out_regB_2_), 
	.A1(FE_OFCN198_UUT_Mpath_out_regA_2_));
   NAND2_X1 U5876 (.ZN(n6575), 
	.A2(n6836), 
	.A1(n6838));
   AND2_X1 U5877 (.ZN(n6829), 
	.A2(n6870), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N159 ));
   AND2_X1 U5878 (.ZN(n6813), 
	.A2(n6814), 
	.A1(n6819));
   OAI22_X1 U5879 (.ZN(n1211), 
	.B2(\UUT/Mpath/the_alu/N468 ), 
	.B1(\UUT/Mpath/the_alu/N520 ), 
	.A2(n2575), 
	.A1(\UUT/Mpath/the_alu/N520 ));
   OR2_X1 U5880 (.ZN(n6754), 
	.A2(\UUT/branch_rega [6]), 
	.A1(n6764));
   INV_X1 U5881 (.ZN(n6721), 
	.A(n6720));
   INV_X1 U5882 (.ZN(n6724), 
	.A(\UUT/branch_rega [6]));
   OAI222_X1 U5883 (.ZN(\UUT/branch_rega [6]), 
	.C2(FE_OFN18_n5441), 
	.C1(n5528), 
	.B2(n2491), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5443));
   NAND2_X1 U5884 (.ZN(n6576), 
	.A2(n6577), 
	.A1(n6545));
   INV_X1 U5885 (.ZN(n6577), 
	.A(n6632));
   OR2_X1 U5886 (.ZN(n6858), 
	.A2(\UUT/branch_rega [25]), 
	.A1(\UUT/branch_rega [26]));
   AND2_X1 U5887 (.ZN(n6591), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[27] ));
   INV_X1 U5888 (.ZN(n6578), 
	.A(n6700));
   NOR2_X1 U5889 (.ZN(n6789), 
	.A2(n6579), 
	.A1(n6742));
   NAND2_X1 U5890 (.ZN(n6579), 
	.A2(n6724), 
	.A1(n6580));
   AND2_X1 U5891 (.ZN(n6580), 
	.A2(n6719), 
	.A1(n6733));
   NAND2_X1 U5892 (.ZN(n6689), 
	.A2(n6581), 
	.A1(n6663));
   OR2_X1 U5893 (.ZN(n6582), 
	.A2(n294), 
	.A1(FE_OFN102_n117));
   OR2_X1 U5894 (.ZN(n6583), 
	.A2(n2727), 
	.A1(n295));
   NAND2_X1 U5895 (.ZN(n6584), 
	.A2(n297), 
	.A1(\UUT/jar_in [23]));
   NAND2_X1 U5896 (.ZN(n6585), 
	.A2(\UUT/branch_rega [23]), 
	.A1(n298));
   NAND2_X1 U5897 (.ZN(n6586), 
	.A2(n6510), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [23]));
   AND3_X1 U5898 (.ZN(n905), 
	.A3(n6584), 
	.A2(n6585), 
	.A1(n6586));
   OAI222_X1 U5899 (.ZN(n6272), 
	.C2(n6035), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n5881), 
	.B1(n6163), 
	.A2(n6026), 
	.A1(n6128));
   NAND3_X1 U5900 (.ZN(n6587), 
	.A3(\UUT/Mcontrol/Operation_decoding32/N2030 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2036 ), 
	.A1(n6028));
   INV_X1 U5901 (.ZN(n931), 
	.A(n6587));
   INV_X1 U5902 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2037 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N2036 ));
   OR2_X1 U5903 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2036 ), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N2029 ), 
	.A1(\UUT/Mcontrol/d_instr [26]));
   OAI222_X1 U5905 (.ZN(\UUT/branch_rega [22]), 
	.C2(n5483), 
	.C1(n5528), 
	.B2(n2098), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5485));
   OR2_X1 U5906 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2086 ), 
	.A2(\UUT/Mcontrol/d_instr [31]), 
	.A1(\UUT/Mcontrol/d_instr [30]));
   OR2_X1 U5913 (.ZN(\UUT/Mcontrol/Operation_decoding32/N2020 ), 
	.A2(\UUT/Mcontrol/d_instr [31]), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1876 ));
   AND2_X1 U5926 (.ZN(n6210), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1963 ), 
	.A1(\UUT/Mcontrol/Operation_decoding32/N1969 ));
   INV_X1 U5927 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1970 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1969 ));
   INV_X1 U5928 (.ZN(\UUT/Mcontrol/Operation_decoding32/N1964 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1963 ));
   OAI222_X1 U5929 (.ZN(n6181), 
	.C2(n6032), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n6035), 
	.B1(n6163), 
	.A2(n6128), 
	.A1(n6029));
   OAI222_X1 U5930 (.ZN(n6188), 
	.C2(n6033), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n6036), 
	.B1(n6163), 
	.A2(n6128), 
	.A1(n6031));
   OAI222_X1 U5931 (.ZN(n6278), 
	.C2(n6036), 
	.C1(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.B2(n5889), 
	.B1(n6163), 
	.A2(n6128), 
	.A1(n6034));
   AND2_X1 U5932 (.ZN(n6589), 
	.A2(n1244), 
	.A1(n1208));
   AND2_X1 U5933 (.ZN(n6590), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[27] ));
   NOR3_X1 U5934 (.ZN(n1243), 
	.A3(n6591), 
	.A2(n6590), 
	.A1(n6589));
   OR2_X1 U5935 (.ZN(n6592), 
	.A2(n5528), 
	.A1(n5468));
   OR2_X1 U5936 (.ZN(n6593), 
	.A2(FE_OFN97_n5529), 
	.A1(n5418));
   OR2_X1 U5937 (.ZN(n6594), 
	.A2(FE_OFN96_n5530), 
	.A1(n5470));
   NAND3_X1 U5938 (.ZN(\UUT/branch_rega [27]), 
	.A3(n6594), 
	.A2(n6593), 
	.A1(n6592));
   AND2_X1 U5939 (.ZN(n6826), 
	.A2(n6851), 
	.A1(n6814));
   INV_X1 U5940 (.ZN(n6851), 
	.A(\UUT/branch_rega [16]));
   NAND2_X1 U5942 (.ZN(n6788), 
	.A2(n6834), 
	.A1(n6803));
   NOR2_X1 U5943 (.ZN(n6735), 
	.A2(n6751), 
	.A1(\UUT/branch_rega [12]));
   INV_X1 U5944 (.ZN(n6803), 
	.A(n6802));
   NAND2_X1 U5945 (.ZN(n6163), 
	.A2(\UUT/Mcontrol/Operation_decoding32/N1975 ), 
	.A1(n6155));
   OR2_X1 U5947 (.ZN(n6596), 
	.A2(n294), 
	.A1(FE_OFN99_n348));
   OR2_X1 U5948 (.ZN(n6597), 
	.A2(n2645), 
	.A1(n295));
   OR2_X1 U5949 (.ZN(n4337), 
	.A2(\localbus/N62 ), 
	.A1(\localbus/N57 ));
   NAND2_X1 U5950 (.ZN(\localbus/N227 ), 
	.A2(\localbus/N338 ), 
	.A1(n4337));
   INV_X1 U5951 (.ZN(\UUT/Mcontrol/d_instr [29]), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1877 ));
   AOI22_X1 U5952 (.ZN(n2061), 
	.B2(n2077), 
	.B1(n6030), 
	.A2(n6085), 
	.A1(n935));
   INV_X1 U5953 (.ZN(\UUT/Mcontrol/d_instr [30]), 
	.A(n6070));
   OR2_X1 U5954 (.ZN(n6598), 
	.A2(n294), 
	.A1(FE_OFN100_n327));
   OR2_X1 U5955 (.ZN(n6599), 
	.A2(n2642), 
	.A1(n295));
   NAND3_X1 U5956 (.ZN(n3003), 
	.A3(n329), 
	.A2(n6599), 
	.A1(n6598));
   NAND2_X1 U5957 (.ZN(n6600), 
	.A2(n297), 
	.A1(\UUT/jar_in [21]));
   NAND2_X1 U5958 (.ZN(n6601), 
	.A2(\UUT/branch_rega [21]), 
	.A1(n298));
   NAND2_X1 U5959 (.ZN(n6602), 
	.A2(n6510), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [21]));
   AND3_X1 U5960 (.ZN(n329), 
	.A3(n6602), 
	.A2(n6601), 
	.A1(n6600));
   OR2_X1 U5961 (.ZN(n6604), 
	.A2(n6603), 
	.A1(FE_OFN187_UUT_branch_rega_1_));
   INV_X1 U5962 (.ZN(n6603), 
	.A(n6790));
   AND2_X1 U5963 (.ZN(n6660), 
	.A2(n6789), 
	.A1(n6605));
   INV_X1 U5964 (.ZN(n6605), 
	.A(n6604));
   OR2_X1 U5965 (.ZN(n6606), 
	.A2(n294), 
	.A1(n495));
   OR2_X1 U5966 (.ZN(n6607), 
	.A2(n2663), 
	.A1(n295));
   NAND3_X1 U5967 (.ZN(n3283), 
	.A3(n497), 
	.A2(n6607), 
	.A1(n6606));
   OR2_X1 U5968 (.ZN(n6609), 
	.A2(FE_OFN97_n5529), 
	.A1(n5416));
   NAND2_X1 U5969 (.ZN(n6611), 
	.A2(n297), 
	.A1(\UUT/jar_in [14]));
   NAND2_X1 U5970 (.ZN(n6612), 
	.A2(\UUT/branch_rega [14]), 
	.A1(n298));
   NAND2_X1 U5971 (.ZN(n6613), 
	.A2(n6511), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [14]));
   AND3_X1 U5972 (.ZN(n497), 
	.A3(n6613), 
	.A2(n6612), 
	.A1(n6611));
   OAI222_X1 U5973 (.ZN(\UUT/branch_rega [14]), 
	.C2(n5510), 
	.C1(n5528), 
	.B2(n2283), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5512));
   OAI222_X1 U5974 (.ZN(\UUT/branch_regb [27]), 
	.C2(n5434), 
	.C1(n5470), 
	.B2(n5432), 
	.B1(n5469), 
	.A2(n5430), 
	.A1(n5468));
   INV_X1 U5975 (.ZN(n6744), 
	.A(\UUT/branch_rega [27]));
   NOR2_X1 U5977 (.ZN(n6614), 
	.A2(n2560), 
	.A1(n2559));
   INV_X1 U5978 (.ZN(n6615), 
	.A(n6614));
   NAND2_X1 U5979 (.ZN(n6616), 
	.A2(n6711), 
	.A1(\UUT/jar_in [15]));
   NAND2_X1 U5980 (.ZN(n6617), 
	.A2(\UUT/branch_rega [15]), 
	.A1(n298));
   NAND2_X1 U5981 (.ZN(n6618), 
	.A2(n6510), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [15]));
   OAI222_X1 U5982 (.ZN(\UUT/branch_rega [15]), 
	.C2(n5507), 
	.C1(n5528), 
	.B2(n2263), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5509));
   INV_X1 U5983 (.ZN(\UUT/Mcontrol/d_instr [31]), 
	.A(n6069));
   INV_X1 U5984 (.ZN(\UUT/Mcontrol/Operation_decoding32/N89 ), 
	.A(\UUT/Mcontrol/Operation_decoding32/N1882 ));
   NAND2_X1 U5985 (.ZN(n6621), 
	.A2(n6665), 
	.A1(n6664));
   NAND2_X1 U5986 (.ZN(\UUT/branch_rega [30]), 
	.A2(n6484), 
	.A1(n6663));
   OR2_X1 U5988 (.ZN(n6623), 
	.A2(n294), 
	.A1(n417));
   OR2_X1 U5989 (.ZN(n6624), 
	.A2(n2654), 
	.A1(n295));
   OR2_X1 U5990 (.ZN(n6665), 
	.A2(FE_OFN96_n5530), 
	.A1(n5458));
   AOI22_X1 U5993 (.ZN(n5468), 
	.B2(n5564), 
	.B1(n5585), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5584));
   NOR2_X1 U5994 (.ZN(n6626), 
	.A2(FE_OFN187_UUT_branch_rega_1_), 
	.A1(n6785));
   AND2_X1 U5995 (.ZN(n6831), 
	.A2(n6627), 
	.A1(n6626));
   AND2_X1 U5996 (.ZN(n6627), 
	.A2(n6876), 
	.A1(n6628));
   INV_X1 U5997 (.ZN(n6628), 
	.A(n6657));
   AND2_X1 U5998 (.ZN(n6629), 
	.A2(n1256), 
	.A1(n1208));
   OR2_X1 U5999 (.ZN(n6630), 
	.A2(n294), 
	.A1(FE_OFN101_n292));
   OR2_X1 U6000 (.ZN(n6631), 
	.A2(n2639), 
	.A1(n295));
   AND2_X1 U6001 (.ZN(n6632), 
	.A2(n1209), 
	.A1(n1208));
   NOR2_X1 U6002 (.ZN(n6634), 
	.A2(n6657), 
	.A1(n6777));
   AND2_X1 U6003 (.ZN(n6681), 
	.A2(n6636), 
	.A1(n6635));
   NOR2_X1 U6004 (.ZN(n6635), 
	.A2(\UUT/branch_rega [29]), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N160 ));
   NOR2_X1 U6005 (.ZN(n6636), 
	.A2(\UUT/branch_rega [28]), 
	.A1(\UUT/branch_rega [27]));
   INV_X1 U6006 (.ZN(\localbus/c1_op[SLAVE][0] ), 
	.A(n6637));
   NOR3_X1 U6008 (.ZN(n909), 
	.A3(n6673), 
	.A2(n6451), 
	.A1(n6672));
   NOR3_X1 U6010 (.ZN(n6642), 
	.A3(n6451), 
	.A2(n6673), 
	.A1(n6672));
   NAND2_X1 U6012 (.ZN(n6644), 
	.A2(n6696), 
	.A1(n6640));
   AOI21_X1 U6013 (.ZN(n6288), 
	.B2(\UUT/Mcontrol/st_logic/N70 ), 
	.B1(n6289), 
	.A(n6291));
   OAI221_X1 U6014 (.ZN(n6647), 
	.C2(n6876), 
	.C1(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.B2(n6648), 
	.B1(n6531), 
	.A(n2558));
   INV_X1 U6015 (.ZN(n6876), 
	.A(\UUT/branch_rega [3]));
   OAI222_X1 U6016 (.ZN(\UUT/branch_rega [7]), 
	.C2(FE_OFN195_n5438), 
	.C1(n5528), 
	.B2(n2468), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5440));
   AND2_X1 U6018 (.ZN(n6651), 
	.A2(\UUT/Mcontrol/st_logic/N96 ), 
	.A1(n6489));
   NOR2_X1 U6019 (.ZN(n6298), 
	.A2(n6651), 
	.A1(n6299));
   NAND2_X1 U6020 (.ZN(n6652), 
	.A2(\UUT/jar_in [8]), 
	.A1(n2324));
   NAND2_X1 U6021 (.ZN(n6653), 
	.A2(\UUT/branch_rega [8]), 
	.A1(\UUT/Mcontrol/st_logic/N109 ));
   AND3_X1 U6022 (.ZN(n631), 
	.A3(n2443), 
	.A2(n6653), 
	.A1(n6652));
   OAI222_X1 U6024 (.ZN(\UUT/branch_rega [8]), 
	.C2(FE_OFN191_n5435), 
	.C1(n5528), 
	.B2(n2445), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5437));
   OAI221_X1 U6025 (.ZN(n6654), 
	.C2(n6724), 
	.C1(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.B2(n6655), 
	.B1(n6531), 
	.A(n2489));
   NAND2_X1 U6027 (.ZN(n6657), 
	.A2(n6832), 
	.A1(n6779));
   NAND2_X1 U6029 (.ZN(n6777), 
	.A2(n6876), 
	.A1(n6660));
   OR2_X1 U6031 (.ZN(n6661), 
	.A2(n294), 
	.A1(n520));
   OR2_X1 U6032 (.ZN(n6662), 
	.A2(n2666), 
	.A1(n295));
   NAND3_X1 U6033 (.ZN(n3323), 
	.A3(n522), 
	.A2(n6662), 
	.A1(n6661));
   OR2_X1 U6034 (.ZN(n6664), 
	.A2(FE_OFN97_n5529), 
	.A1(n5415));
   AND2_X1 U6035 (.ZN(n6666), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[30] ));
   NAND2_X1 U6036 (.ZN(n6667), 
	.A2(n297), 
	.A1(\UUT/jar_in [13]));
   NAND2_X1 U6037 (.ZN(n6668), 
	.A2(\UUT/branch_rega [13]), 
	.A1(n298));
   NAND2_X1 U6038 (.ZN(n6669), 
	.A2(n6510), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/Bta [13]));
   AND3_X1 U6039 (.ZN(n522), 
	.A3(n6669), 
	.A2(n6668), 
	.A1(n6667));
   OAI222_X1 U6040 (.ZN(\UUT/branch_rega [13]), 
	.C2(n5513), 
	.C1(n5528), 
	.B2(n2303), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5515));
   INV_X1 U6041 (.ZN(n6670), 
	.A(n6705));
   NAND2_X1 U6042 (.ZN(n6671), 
	.A2(n6670), 
	.A1(n6688));
   AND2_X1 U6043 (.ZN(n6673), 
	.A2(\UUT/branch_rega [9]), 
	.A1(\UUT/Mcontrol/st_logic/N109 ));
   OR2_X1 U6044 (.ZN(n6865), 
	.A2(\UUT/branch_rega [12]), 
	.A1(\UUT/branch_rega [13]));
   OAI222_X1 U6047 (.ZN(\UUT/branch_rega [12]), 
	.C2(n5516), 
	.C1(n5528), 
	.B2(n2353), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5518));
   INV_X1 U6048 (.ZN(n6859), 
	.A(n6858));
   AND2_X1 U6049 (.ZN(n6677), 
	.A2(\UUT/branch_rega [10]), 
	.A1(\UUT/Mcontrol/st_logic/N109 ));
   OAI222_X1 U6050 (.ZN(\UUT/branch_rega [10]), 
	.C2(FE_OFN193_n5522), 
	.C1(n5528), 
	.B2(n2399), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5524));
   NOR2_X1 U6052 (.ZN(n906), 
	.A2(n6615), 
	.A1(n6479));
   OR2_X1 U6054 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N160 ), 
	.A2(\UUT/branch_rega [30]), 
	.A1(n6489));
   INV_X1 U6055 (.ZN(n6680), 
	.A(n6809));
   NAND2_X1 U6056 (.ZN(n6725), 
	.A2(n6682), 
	.A1(n6681));
   NOR2_X1 U6057 (.ZN(n6682), 
	.A2(n6680), 
	.A1(\UUT/branch_rega [26]));
   NAND2_X1 U6059 (.ZN(n6684), 
	.A2(\UUT/jar_in [2]), 
	.A1(n2324));
   NAND2_X1 U6060 (.ZN(n6685), 
	.A2(\UUT/branch_rega [2]), 
	.A1(\UUT/Mcontrol/st_logic/N109 ));
   AND3_X1 U6061 (.ZN(n763), 
	.A3(n2327), 
	.A2(n6685), 
	.A1(n6684));
   OAI222_X1 U6062 (.ZN(\UUT/branch_rega [2]), 
	.C2(FE_OFN189_n5459), 
	.C1(n5528), 
	.B2(n2330), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5461));
   NOR2_X1 U6063 (.ZN(n6845), 
	.A2(n6488), 
	.A1(n6689));
   OR2_X1 U6064 (.ZN(n6691), 
	.A2(n294), 
	.A1(n439));
   OR2_X1 U6065 (.ZN(n6692), 
	.A2(n2657), 
	.A1(n295));
   NAND3_X1 U6066 (.ZN(n3203), 
	.A3(n442), 
	.A2(n6692), 
	.A1(n6691));
   NAND2_X1 U6067 (.ZN(n6694), 
	.A2(n863), 
	.A1(n137));
   NAND2_X1 U6068 (.ZN(n6695), 
	.A2(n1206), 
	.A1(n1205));
   INV_X1 U6069 (.ZN(n6696), 
	.A(n6695));
   OR2_X1 U6070 (.ZN(n6794), 
	.A2(\UUT/branch_rega [3]), 
	.A1(n6799));
   OAI222_X1 U6071 (.ZN(\UUT/branch_rega [3]), 
	.C2(FE_OFN30_n5450), 
	.C1(n5528), 
	.B2(n2565), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5452));
   OR2_X1 U6072 (.ZN(\UUT/Mpath/the_alu/N157 ), 
	.A2(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.A1(FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_));
   AND2_X1 U6073 (.ZN(\UUT/Mpath/the_alu/N125 ), 
	.A2(FE_OFN182_UUT_Mpath_out_regB_0_), 
	.A1(FE_OFCN205_FE_OFN104_UUT_Mpath_out_regA_0_));
   NOR2_X1 U6074 (.ZN(n6697), 
	.A2(\UUT/branch_rega [22]), 
	.A1(\UUT/branch_rega [21]));
   AND2_X1 U6075 (.ZN(n6699), 
	.A2(n6744), 
	.A1(n6877));
   AND2_X1 U6077 (.ZN(n6700), 
	.A2(\UUT/Mpath/N119 ), 
	.A1(n5591));
   NAND2_X1 U6080 (.ZN(n6703), 
	.A2(\UUT/jar_in [11]), 
	.A1(n2324));
   NAND2_X1 U6081 (.ZN(n6704), 
	.A2(\UUT/branch_rega [11]), 
	.A1(\UUT/Mcontrol/st_logic/N109 ));
   OR2_X1 U6082 (.ZN(n6705), 
	.A2(\UUT/branch_rega [13]), 
	.A1(\UUT/branch_rega [14]));
   AND2_X1 U6084 (.ZN(n6707), 
	.A2(n1238), 
	.A1(n1208));
   AND2_X1 U6085 (.ZN(n6708), 
	.A2(n1210), 
	.A1(\UUT/Mpath/the_alu/diff[26] ));
   AND2_X1 U6086 (.ZN(n6709), 
	.A2(FE_OFN87_n1211), 
	.A1(\UUT/Mpath/the_alu/sum[26] ));
   NOR3_X1 U6087 (.ZN(n1237), 
	.A3(n6709), 
	.A2(n6708), 
	.A1(n6707));
   OAI222_X1 U6088 (.ZN(\UUT/branch_rega [11]), 
	.C2(n5519), 
	.C1(n5528), 
	.B2(n2376), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5521));
   INV_X1 U6089 (.ZN(n694), 
	.A(n6848));
   OAI222_X1 U6090 (.ZN(\UUT/branch_regb [26]), 
	.C2(n5434), 
	.C1(n5473), 
	.B2(n5432), 
	.B1(n5472), 
	.A2(n5430), 
	.A1(n5471));
   NAND2_X1 U6092 (.ZN(n546), 
	.A2(n978), 
	.A1(net54875));
   INV_X4 U6093 (.ZN(n295), 
	.A(FE_OFCN206_FE_OFN186_n546));
   INV_X1 U6094 (.ZN(n6712), 
	.A(n6718));
   AND2_X1 U6096 (.ZN(net56414), 
	.A2(n6883), 
	.A1(n6882));
   INV_X1 U6097 (.ZN(n6717), 
	.A(n6726));
   NAND2_X1 U6098 (.ZN(n6718), 
	.A2(n6717), 
	.A1(n6854));
   AND2_X1 U6099 (.ZN(n6732), 
	.A2(n6733), 
	.A1(n6740));
   OR2_X1 U6100 (.ZN(n6792), 
	.A2(\UUT/branch_rega [21]), 
	.A1(n6796));
   INV_X1 U6101 (.ZN(n6834), 
	.A(\UUT/branch_rega [18]));
   OAI222_X1 U6102 (.ZN(\UUT/branch_rega [18]), 
	.C2(n5498), 
	.C1(n5528), 
	.B2(n2203), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5500));
   AOI222_X1 U6103 (.ZN(n5498), 
	.C2(n5612), 
	.C1(\UUT/Mpath/out_jar[18] ), 
	.B2(\UUT/Mpath/N119 ), 
	.B1(n415), 
	.A2(n5564), 
	.A1(n6134));
   INV_X1 U6104 (.ZN(n6719), 
	.A(n6727));
   NOR2_X1 U6106 (.ZN(n6723), 
	.A2(n6752), 
	.A1(n6730));
   NAND2_X1 U6108 (.ZN(n6726), 
	.A2(n6724), 
	.A1(n6732));
   NAND2_X1 U6109 (.ZN(n6727), 
	.A2(n6805), 
	.A1(n6728));
   AND2_X1 U6110 (.ZN(n6728), 
	.A2(n6729), 
	.A1(n6757));
   INV_X1 U6111 (.ZN(n6729), 
	.A(n6734));
   NAND2_X1 U6112 (.ZN(n6730), 
	.A2(n6731), 
	.A1(n6757));
   INV_X1 U6113 (.ZN(n6731), 
	.A(n6737));
   INV_X1 U6114 (.ZN(n6733), 
	.A(\UUT/branch_rega [7]));
   NAND2_X1 U6115 (.ZN(n6734), 
	.A2(n6825), 
	.A1(n6735));
   OR2_X1 U6116 (.ZN(n6737), 
	.A2(\UUT/branch_rega [9]), 
	.A1(\UUT/branch_rega [8]));
   AND2_X1 U6119 (.ZN(n6740), 
	.A2(n6741), 
	.A1(n6746));
   INV_X1 U6120 (.ZN(n6741), 
	.A(\UUT/branch_rega [8]));
   NAND2_X1 U6121 (.ZN(n6742), 
	.A2(n6885), 
	.A1(n6822));
   NAND2_X1 U6123 (.ZN(n6745), 
	.A2(n6852), 
	.A1(n6744));
   INV_X1 U6124 (.ZN(n6885), 
	.A(\UUT/branch_rega [23]));
   OAI222_X1 U6125 (.ZN(\UUT/branch_rega [23]), 
	.C2(n5480), 
	.C1(n5528), 
	.B2(n2078), 
	.B1(FE_OFN97_n5529), 
	.A2(FE_OFN96_n5530), 
	.A1(n5482));
   AND2_X1 U6126 (.ZN(n6746), 
	.A2(n6747), 
	.A1(n6756));
   INV_X1 U6127 (.ZN(n6747), 
	.A(\UUT/branch_rega [9]));
   INV_X1 U6128 (.ZN(n6748), 
	.A(n6759));
   NAND2_X1 U6129 (.ZN(n6749), 
	.A2(n6748), 
	.A1(n6880));
   INV_X1 U6130 (.ZN(n6750), 
	.A(n6749));
   NAND2_X1 U6131 (.ZN(n6751), 
	.A2(n6750), 
	.A1(n6830));
   OR2_X1 U6132 (.ZN(n6752), 
	.A2(n6754), 
	.A1(\UUT/branch_rega [7]));
   AND2_X1 U6134 (.ZN(n6756), 
	.A2(n6757), 
	.A1(n6761));
   INV_X1 U6135 (.ZN(n6757), 
	.A(\UUT/branch_rega [10]));
   NAND2_X1 U6137 (.ZN(n6759), 
	.A2(n6846), 
	.A1(n6763));
   INV_X1 U6138 (.ZN(n6760), 
	.A(n6824));
   NOR2_X1 U6139 (.ZN(n6761), 
	.A2(n6760), 
	.A1(n6767));
   NOR2_X1 U6141 (.ZN(n6763), 
	.A2(\UUT/branch_rega [15]), 
	.A1(n6769));
   INV_X1 U6142 (.ZN(n6833), 
	.A(\UUT/branch_rega [19]));
   OR2_X1 U6146 (.ZN(n6764), 
	.A2(n6765), 
	.A1(\UUT/branch_rega [5]));
   INV_X1 U6147 (.ZN(n6765), 
	.A(n6774));
   OR2_X1 U6148 (.ZN(n6767), 
	.A2(\UUT/branch_rega [14]), 
	.A1(n6771));
   NAND2_X1 U6151 (.ZN(n6771), 
	.A2(n6826), 
	.A1(n6772));
   NOR2_X1 U6152 (.ZN(n6772), 
	.A2(\UUT/branch_rega [17]), 
	.A1(n6786));
   NOR2_X1 U6154 (.ZN(n6774), 
	.A2(n6832), 
	.A1(n6787));
   INV_X1 U6155 (.ZN(n6775), 
	.A(\UUT/branch_rega [17]));
   NAND2_X1 U6156 (.ZN(n6776), 
	.A2(n6775), 
	.A1(n6781));
   INV_X1 U6158 (.ZN(n6779), 
	.A(\UUT/branch_rega [2]));
   INV_X1 U6159 (.ZN(n6877), 
	.A(\UUT/branch_rega [24]));
   OAI222_X1 U6160 (.ZN(\UUT/branch_rega [24]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5479), 
	.B2(FE_OFN97_n5529), 
	.B1(n5421), 
	.A2(n5528), 
	.A1(n5477));
   NOR2_X1 U6162 (.ZN(n6781), 
	.A2(\UUT/branch_rega [19]), 
	.A1(n6788));
   NAND2_X1 U6166 (.ZN(n6785), 
	.A2(n6790), 
	.A1(n6789));
   OR2_X1 U6167 (.ZN(n6786), 
	.A2(n6792), 
	.A1(\UUT/branch_rega [22]));
   AND2_X1 U6168 (.ZN(n6790), 
	.A2(n6854), 
	.A1(n6868));
   OR2_X1 U6172 (.ZN(n6796), 
	.A2(n6797), 
	.A1(\UUT/branch_rega [20]));
   INV_X1 U6173 (.ZN(n6797), 
	.A(n6801));
   OR2_X1 U6174 (.ZN(n6799), 
	.A2(\UUT/branch_rega [2]), 
	.A1(FE_OFN187_UUT_branch_rega_1_));
   AND2_X1 U6176 (.ZN(n6801), 
	.A2(n6833), 
	.A1(n6834));
   OR2_X1 U6178 (.ZN(n6802), 
	.A2(\UUT/branch_rega [20]), 
	.A1(\UUT/branch_rega [21]));
   OR2_X1 U6179 (.ZN(n6804), 
	.A2(\UUT/branch_rega [8]), 
	.A1(\UUT/branch_rega [9]));
   INV_X1 U6180 (.ZN(n6805), 
	.A(n6804));
   AND2_X1 U6182 (.ZN(n6809), 
	.A2(n6816), 
	.A1(n6885));
   INV_X1 U6184 (.ZN(n6816), 
	.A(n6815));
   INV_X1 U6188 (.ZN(n6814), 
	.A(\UUT/branch_rega [15]));
   OR2_X1 U6189 (.ZN(n6815), 
	.A2(\UUT/branch_rega [24]), 
	.A1(\UUT/branch_rega [25]));
   AND2_X1 U6194 (.ZN(n6822), 
	.A2(n6872), 
	.A1(n6877));
   AND2_X1 U6196 (.ZN(n6824), 
	.A2(n6866), 
	.A1(n6825));
   INV_X1 U6197 (.ZN(n6825), 
	.A(\UUT/branch_rega [11]));
   INV_X1 U6200 (.ZN(n6830), 
	.A(\UUT/branch_rega [22]));
   INV_X1 U6202 (.ZN(n6836), 
	.A(\UUT/branch_rega [20]));
   OR2_X1 U6206 (.ZN(n6843), 
	.A2(n861), 
	.A1(n133));
   OR2_X1 U6207 (.ZN(n6844), 
	.A2(n135), 
	.A1(n5686));
   OAI222_X1 U6208 (.ZN(\UUT/branch_rega [26]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5473), 
	.B2(FE_OFN97_n5529), 
	.B1(n5419), 
	.A2(n5528), 
	.A1(n5471));
   OAI222_X1 U6209 (.ZN(\UUT/branch_rega [25]), 
	.C2(FE_OFN96_n5530), 
	.C1(n5476), 
	.B2(FE_OFN97_n5529), 
	.B1(n5420), 
	.A2(n5528), 
	.A1(n5474));
   INV_X1 U6210 (.ZN(n6846), 
	.A(\UUT/branch_rega [14]));
   INV_X1 U6211 (.ZN(n2324), 
	.A(n907));
   OR2_X1 U6212 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N125 ), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N116 ), 
	.A1(\UUT/Mcontrol/st_logic/N65 ));
   NAND2_X1 U6213 (.ZN(n6850), 
	.A2(n6859), 
	.A1(n6699));
   INV_X1 U6214 (.ZN(n6852), 
	.A(\UUT/branch_rega [25]));
   INV_X1 U6215 (.ZN(n6861), 
	.A(n6488));
   INV_X1 U6216 (.ZN(n6860), 
	.A(n6489));
   NAND2_X1 U6217 (.ZN(n6887), 
	.A2(n6863), 
	.A1(n6862));
   AND2_X1 U6218 (.ZN(n6863), 
	.A2(n6890), 
	.A1(n6864));
   INV_X1 U6219 (.ZN(n6864), 
	.A(n6889));
   INV_X1 U6220 (.ZN(n6866), 
	.A(n6865));
   NOR2_X1 U6222 (.ZN(n6870), 
	.A2(n6875), 
	.A1(\UUT/branch_rega [30]));
   INV_X1 U6226 (.ZN(n6880), 
	.A(\UUT/branch_rega [13]));
   NAND2_X1 U6227 (.ZN(n6881), 
	.A2(n6894), 
	.A1(n6893));
   INV_X1 U6228 (.ZN(n6882), 
	.A(n6881));
   NAND2_X1 U6229 (.ZN(n6883), 
	.A2(n948), 
	.A1(n137));
   NAND2_X1 U6231 (.ZN(n6296), 
	.A2(n6888), 
	.A1(n6887));
   OR2_X1 U6232 (.ZN(n6888), 
	.A2(n6861), 
	.A1(\UUT/Mcontrol/Nextpc_decoding/N247 ));
   OR2_X1 U6233 (.ZN(n6889), 
	.A2(\UUT/Mcontrol/Nextpc_decoding/N247 ), 
	.A1(\UUT/branch_rega [0]));
   NOR2_X1 U6234 (.ZN(n6890), 
	.A2(FE_OFN187_UUT_branch_rega_1_), 
	.A1(\UUT/branch_rega [2]));
   AOI21_X2 U6235 (.ZN(n6299), 
	.B2(\UUT/Mcontrol/st_logic/N102 ), 
	.B1(\UUT/Mcontrol/Nextpc_decoding/N32 ), 
	.A(\UUT/Mcontrol/st_logic/N96 ));
   INV_X1 U6237 (.ZN(\UUT/Mcontrol/Nextpc_decoding/N159 ), 
	.A(\UUT/branch_rega [31]));
   OR2_X1 U6238 (.ZN(n6893), 
	.A2(n1142), 
	.A1(n133));
   OR2_X1 U6239 (.ZN(n6894), 
	.A2(n135), 
	.A1(n5685));
   INV_X1 U6243 (.ZN(net54843), 
	.A(net54953));
   INV_X1 U6244 (.ZN(net54845), 
	.A(net54953));
   INV_X1 U6245 (.ZN(net54847), 
	.A(FE_OFN10_net54953));
   INV_X1 U6246 (.ZN(net54849), 
	.A(FE_OFN10_net54953));
   INV_X1 U6247 (.ZN(net54851), 
	.A(FE_OFN10_net54953));
   INV_X1 U6248 (.ZN(net54853), 
	.A(FE_OFN10_net54953));
   INV_X1 U6249 (.ZN(net54855), 
	.A(FE_OFN10_net54953));
   INV_X1 U6250 (.ZN(net54857), 
	.A(FE_OFN10_net54953));
   INV_X1 U6251 (.ZN(net54859), 
	.A(FE_OFN12_net54953));
   INV_X1 U6252 (.ZN(net54861), 
	.A(FE_OFN12_net54953));
   INV_X1 U6253 (.ZN(net54863), 
	.A(FE_OFN12_net54953));
   INV_X1 U6254 (.ZN(net54865), 
	.A(net54953));
   INV_X1 U6255 (.ZN(net54867), 
	.A(net54953));
   INV_X1 U6256 (.ZN(net54869), 
	.A(FE_OFN12_net54953));
   INV_X1 U6257 (.ZN(net54871), 
	.A(net54953));
   INV_X1 U6258 (.ZN(net54873), 
	.A(FE_OFN10_net54953));
   INV_X1 U6259 (.ZN(net54875), 
	.A(FE_OFN11_net54953));
   INV_X1 U6260 (.ZN(net54877), 
	.A(FE_OFN12_net54953));
   INV_X1 U6261 (.ZN(net54879), 
	.A(net54953));
   INV_X1 U6262 (.ZN(net54881), 
	.A(FE_OFN12_net54953));
   INV_X1 U6263 (.ZN(net54883), 
	.A(FE_OFN10_net54953));
   INV_X1 U6264 (.ZN(net54885), 
	.A(net54953));
   INV_X1 U6265 (.ZN(net54887), 
	.A(FE_OFN12_net54953));
   INV_X1 U6266 (.ZN(net54889), 
	.A(FE_OFN12_net54953));
   INV_X1 U6267 (.ZN(net54891), 
	.A(FE_OFN12_net54953));
   INV_X1 U6268 (.ZN(net54893), 
	.A(net54953));
   INV_X1 U6269 (.ZN(net54895), 
	.A(FE_OFN12_net54953));
   NAND4_X1 U6294 (.ZN(\localbus/N61 ), 
	.A4(\localbus/c1_addr_outbus[28] ), 
	.A3(\localbus/c1_addr_outbus[29] ), 
	.A2(\localbus/c1_addr_outbus[30] ), 
	.A1(n6595));
   OAI21_X1 U6295 (.ZN(n6902), 
	.B2(\localbus/c1_addr_outbus[28] ), 
	.B1(\localbus/c1_addr_outbus[29] ), 
	.A(\localbus/c1_addr_outbus[30] ));
   NAND2_X1 U6297 (.ZN(\localbus/N60 ), 
	.A2(n6425), 
	.A1(n6902));
   INV_X1 U6298 (.ZN(n6910), 
	.A(n6903));
   OR2_X1 U6299 (.ZN(n6904), 
	.A2(\localbus/c1_addr_outbus[13] ), 
	.A1(\localbus/c1_addr_outbus[14] ));
   AOI221_X1 U6300 (.ZN(n6908), 
	.C2(n6904), 
	.C1(\localbus/c1_addr_outbus[16] ), 
	.B2(\localbus/c1_addr_outbus[15] ), 
	.B1(\localbus/c1_addr_outbus[16] ), 
	.A(n6910));
   NOR4_X1 U6301 (.ZN(n6907), 
	.A4(\localbus/c1_addr_outbus[17] ), 
	.A3(\localbus/c1_addr_outbus[18] ), 
	.A2(\localbus/c1_addr_outbus[19] ), 
	.A1(\localbus/c1_addr_outbus[20] ));
   NOR4_X1 U6302 (.ZN(n6906), 
	.A4(\localbus/c1_addr_outbus[21] ), 
	.A3(\localbus/c1_addr_outbus[22] ), 
	.A2(\localbus/c1_addr_outbus[23] ), 
	.A1(\localbus/c1_addr_outbus[24] ));
   NOR4_X1 U6303 (.ZN(n6905), 
	.A4(\localbus/c1_addr_outbus[25] ), 
	.A3(\localbus/c1_addr_outbus[26] ), 
	.A2(\localbus/c1_addr_outbus[27] ), 
	.A1(\localbus/c1_addr_outbus[28] ));
   NOR2_X1 U6304 (.ZN(n6914), 
	.A2(\localbus/c1_addr_outbus[30] ), 
	.A1(n6595));
   NOR4_X1 U6305 (.ZN(n6912), 
	.A4(\localbus/c1_addr_outbus[16] ), 
	.A3(\localbus/c1_addr_outbus[17] ), 
	.A2(\localbus/c1_addr_outbus[18] ), 
	.A1(\localbus/c1_addr_outbus[19] ));
   NOR4_X1 U6306 (.ZN(n6911), 
	.A4(\localbus/c1_addr_outbus[20] ), 
	.A3(\localbus/c1_addr_outbus[21] ), 
	.A2(\localbus/c1_addr_outbus[22] ), 
	.A1(\localbus/c1_addr_outbus[23] ));
   AND2_X1 U6307 (.ZN(n6913), 
	.A2(n6911), 
	.A1(n6912));
   OAI22_X1 U6308 (.ZN(\localbus/N55 ), 
	.B2(n6914), 
	.B1(n6913), 
	.A2(n6914), 
	.A1(n6915));
   XNOR2_X1 U6309 (.ZN(n6918), 
	.B(\UUT/rs2_addr [0]), 
	.A(\UUT/Mcontrol/x_rd[0] ));
   XNOR2_X1 U6310 (.ZN(n6917), 
	.B(\UUT/rs2_addr [2]), 
	.A(\UUT/Mcontrol/x_rd[2] ));
   XNOR2_X1 U6311 (.ZN(n6916), 
	.B(\UUT/rs2_addr [1]), 
	.A(\UUT/Mcontrol/x_rd[1] ));
   NAND3_X1 U6312 (.ZN(n6921), 
	.A3(n6916), 
	.A2(n6917), 
	.A1(n6918));
   XOR2_X1 U6313 (.Z(n6920), 
	.B(\UUT/rs2_addr [3]), 
	.A(\UUT/Mcontrol/x_rd[3] ));
   XOR2_X1 U6314 (.Z(n6919), 
	.B(\UUT/rs2_addr [4]), 
	.A(\UUT/Mcontrol/x_rd[4] ));
   NOR3_X1 U6315 (.ZN(\UUT/Mcontrol/bp_logicB/N2 ), 
	.A3(n6919), 
	.A2(n6920), 
	.A1(n6921));
   XNOR2_X1 U6316 (.ZN(n6924), 
	.B(\UUT/rs2_addr [0]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[0] ));
   XNOR2_X1 U6317 (.ZN(n6923), 
	.B(\UUT/rs2_addr [2]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[2] ));
   XNOR2_X1 U6318 (.ZN(n6922), 
	.B(\UUT/rs2_addr [1]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[1] ));
   NAND3_X1 U6319 (.ZN(n6927), 
	.A3(n6922), 
	.A2(n6923), 
	.A1(n6924));
   XOR2_X1 U6320 (.Z(n6926), 
	.B(\UUT/rs2_addr [3]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[3] ));
   XOR2_X1 U6321 (.Z(n6925), 
	.B(\UUT/rs2_addr [4]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[4] ));
   NOR3_X1 U6322 (.ZN(\UUT/Mcontrol/bp_logicB/N3 ), 
	.A3(n6925), 
	.A2(n6926), 
	.A1(n6927));
   XNOR2_X1 U6323 (.ZN(n6930), 
	.B(\UUT/rs1_addr [0]), 
	.A(\UUT/Mcontrol/x_rd[0] ));
   XNOR2_X1 U6324 (.ZN(n6929), 
	.B(\UUT/rs1_addr [2]), 
	.A(\UUT/Mcontrol/x_rd[2] ));
   XNOR2_X1 U6325 (.ZN(n6928), 
	.B(FE_OFN98_UUT_rs1_addr_1_), 
	.A(\UUT/Mcontrol/x_rd[1] ));
   NAND3_X1 U6326 (.ZN(n6933), 
	.A3(n6928), 
	.A2(n6929), 
	.A1(n6930));
   XOR2_X1 U6327 (.Z(n6932), 
	.B(FE_OFCN199_UUT_rs1_addr_3_), 
	.A(\UUT/Mcontrol/x_rd[3] ));
   XOR2_X1 U6328 (.Z(n6931), 
	.B(\UUT/rs1_addr [4]), 
	.A(\UUT/Mcontrol/x_rd[4] ));
   NOR3_X1 U6329 (.ZN(\UUT/Mcontrol/bp_logicA/N2 ), 
	.A3(n6931), 
	.A2(n6932), 
	.A1(n6933));
   XNOR2_X1 U6330 (.ZN(n6936), 
	.B(\UUT/rs1_addr [0]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[0] ));
   XNOR2_X1 U6331 (.ZN(n6935), 
	.B(\UUT/rs1_addr [2]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[2] ));
   XNOR2_X1 U6332 (.ZN(n6934), 
	.B(FE_OFN98_UUT_rs1_addr_1_), 
	.A(\UUT/Mcontrol/m_sampled_xrd[1] ));
   NAND3_X1 U6333 (.ZN(n6939), 
	.A3(n6934), 
	.A2(n6935), 
	.A1(n6936));
   XOR2_X1 U6334 (.Z(n6938), 
	.B(FE_OFCN199_UUT_rs1_addr_3_), 
	.A(\UUT/Mcontrol/m_sampled_xrd[3] ));
   XOR2_X1 U6335 (.Z(n6937), 
	.B(\UUT/rs1_addr [4]), 
	.A(\UUT/Mcontrol/m_sampled_xrd[4] ));
   NOR3_X1 U6336 (.ZN(\UUT/Mcontrol/bp_logicA/N3 ), 
	.A3(n6937), 
	.A2(n6938), 
	.A1(n6939));
endmodule

